// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

module IssueUnitCollapsing_2(
  input         clock,
                reset,
                io_dis_uops_0_valid,
  input  [6:0]  io_dis_uops_0_bits_uopc,
  input         io_dis_uops_0_bits_is_rvc,
  input  [9:0]  io_dis_uops_0_bits_fu_code,
  input         io_dis_uops_0_bits_is_br,
                io_dis_uops_0_bits_is_jalr,
                io_dis_uops_0_bits_is_jal,
                io_dis_uops_0_bits_is_sfb,
  input  [19:0] io_dis_uops_0_bits_br_mask,
  input  [4:0]  io_dis_uops_0_bits_br_tag,
  input  [5:0]  io_dis_uops_0_bits_ftq_idx,
  input         io_dis_uops_0_bits_edge_inst,
  input  [5:0]  io_dis_uops_0_bits_pc_lob,
  input         io_dis_uops_0_bits_taken,
  input  [19:0] io_dis_uops_0_bits_imm_packed,
  input  [6:0]  io_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_dis_uops_0_bits_ldq_idx,
                io_dis_uops_0_bits_stq_idx,
  input  [6:0]  io_dis_uops_0_bits_pdst,
                io_dis_uops_0_bits_prs1,
                io_dis_uops_0_bits_prs2,
                io_dis_uops_0_bits_prs3,
  input         io_dis_uops_0_bits_prs1_busy,
                io_dis_uops_0_bits_prs2_busy,
                io_dis_uops_0_bits_exception,
                io_dis_uops_0_bits_bypassable,
  input  [4:0]  io_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_dis_uops_0_bits_mem_size,
  input         io_dis_uops_0_bits_mem_signed,
                io_dis_uops_0_bits_is_fence,
                io_dis_uops_0_bits_is_fencei,
                io_dis_uops_0_bits_is_amo,
                io_dis_uops_0_bits_uses_ldq,
                io_dis_uops_0_bits_uses_stq,
                io_dis_uops_0_bits_ldst_val,
  input  [1:0]  io_dis_uops_0_bits_dst_rtype,
                io_dis_uops_0_bits_lrs1_rtype,
                io_dis_uops_0_bits_lrs2_rtype,
  input         io_dis_uops_0_bits_fp_val,
                io_dis_uops_1_valid,
  input  [6:0]  io_dis_uops_1_bits_uopc,
  input         io_dis_uops_1_bits_is_rvc,
  input  [9:0]  io_dis_uops_1_bits_fu_code,
  input         io_dis_uops_1_bits_is_br,
                io_dis_uops_1_bits_is_jalr,
                io_dis_uops_1_bits_is_jal,
                io_dis_uops_1_bits_is_sfb,
  input  [19:0] io_dis_uops_1_bits_br_mask,
  input  [4:0]  io_dis_uops_1_bits_br_tag,
  input  [5:0]  io_dis_uops_1_bits_ftq_idx,
  input         io_dis_uops_1_bits_edge_inst,
  input  [5:0]  io_dis_uops_1_bits_pc_lob,
  input         io_dis_uops_1_bits_taken,
  input  [19:0] io_dis_uops_1_bits_imm_packed,
  input  [6:0]  io_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_dis_uops_1_bits_ldq_idx,
                io_dis_uops_1_bits_stq_idx,
  input  [6:0]  io_dis_uops_1_bits_pdst,
                io_dis_uops_1_bits_prs1,
                io_dis_uops_1_bits_prs2,
                io_dis_uops_1_bits_prs3,
  input         io_dis_uops_1_bits_prs1_busy,
                io_dis_uops_1_bits_prs2_busy,
                io_dis_uops_1_bits_exception,
                io_dis_uops_1_bits_bypassable,
  input  [4:0]  io_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_dis_uops_1_bits_mem_size,
  input         io_dis_uops_1_bits_mem_signed,
                io_dis_uops_1_bits_is_fence,
                io_dis_uops_1_bits_is_fencei,
                io_dis_uops_1_bits_is_amo,
                io_dis_uops_1_bits_uses_ldq,
                io_dis_uops_1_bits_uses_stq,
                io_dis_uops_1_bits_ldst_val,
  input  [1:0]  io_dis_uops_1_bits_dst_rtype,
                io_dis_uops_1_bits_lrs1_rtype,
                io_dis_uops_1_bits_lrs2_rtype,
  input         io_dis_uops_1_bits_fp_val,
                io_dis_uops_2_valid,
  input  [6:0]  io_dis_uops_2_bits_uopc,
  input         io_dis_uops_2_bits_is_rvc,
  input  [9:0]  io_dis_uops_2_bits_fu_code,
  input         io_dis_uops_2_bits_is_br,
                io_dis_uops_2_bits_is_jalr,
                io_dis_uops_2_bits_is_jal,
                io_dis_uops_2_bits_is_sfb,
  input  [19:0] io_dis_uops_2_bits_br_mask,
  input  [4:0]  io_dis_uops_2_bits_br_tag,
  input  [5:0]  io_dis_uops_2_bits_ftq_idx,
  input         io_dis_uops_2_bits_edge_inst,
  input  [5:0]  io_dis_uops_2_bits_pc_lob,
  input         io_dis_uops_2_bits_taken,
  input  [19:0] io_dis_uops_2_bits_imm_packed,
  input  [6:0]  io_dis_uops_2_bits_rob_idx,
  input  [4:0]  io_dis_uops_2_bits_ldq_idx,
                io_dis_uops_2_bits_stq_idx,
  input  [6:0]  io_dis_uops_2_bits_pdst,
                io_dis_uops_2_bits_prs1,
                io_dis_uops_2_bits_prs2,
                io_dis_uops_2_bits_prs3,
  input         io_dis_uops_2_bits_prs1_busy,
                io_dis_uops_2_bits_prs2_busy,
                io_dis_uops_2_bits_exception,
                io_dis_uops_2_bits_bypassable,
  input  [4:0]  io_dis_uops_2_bits_mem_cmd,
  input  [1:0]  io_dis_uops_2_bits_mem_size,
  input         io_dis_uops_2_bits_mem_signed,
                io_dis_uops_2_bits_is_fence,
                io_dis_uops_2_bits_is_fencei,
                io_dis_uops_2_bits_is_amo,
                io_dis_uops_2_bits_uses_ldq,
                io_dis_uops_2_bits_uses_stq,
                io_dis_uops_2_bits_ldst_val,
  input  [1:0]  io_dis_uops_2_bits_dst_rtype,
                io_dis_uops_2_bits_lrs1_rtype,
                io_dis_uops_2_bits_lrs2_rtype,
  input         io_dis_uops_2_bits_fp_val,
                io_dis_uops_3_valid,
  input  [6:0]  io_dis_uops_3_bits_uopc,
  input         io_dis_uops_3_bits_is_rvc,
  input  [9:0]  io_dis_uops_3_bits_fu_code,
  input         io_dis_uops_3_bits_is_br,
                io_dis_uops_3_bits_is_jalr,
                io_dis_uops_3_bits_is_jal,
                io_dis_uops_3_bits_is_sfb,
  input  [19:0] io_dis_uops_3_bits_br_mask,
  input  [4:0]  io_dis_uops_3_bits_br_tag,
  input  [5:0]  io_dis_uops_3_bits_ftq_idx,
  input         io_dis_uops_3_bits_edge_inst,
  input  [5:0]  io_dis_uops_3_bits_pc_lob,
  input         io_dis_uops_3_bits_taken,
  input  [19:0] io_dis_uops_3_bits_imm_packed,
  input  [6:0]  io_dis_uops_3_bits_rob_idx,
  input  [4:0]  io_dis_uops_3_bits_ldq_idx,
                io_dis_uops_3_bits_stq_idx,
  input  [6:0]  io_dis_uops_3_bits_pdst,
                io_dis_uops_3_bits_prs1,
                io_dis_uops_3_bits_prs2,
                io_dis_uops_3_bits_prs3,
  input         io_dis_uops_3_bits_prs1_busy,
                io_dis_uops_3_bits_prs2_busy,
                io_dis_uops_3_bits_exception,
                io_dis_uops_3_bits_bypassable,
  input  [4:0]  io_dis_uops_3_bits_mem_cmd,
  input  [1:0]  io_dis_uops_3_bits_mem_size,
  input         io_dis_uops_3_bits_mem_signed,
                io_dis_uops_3_bits_is_fence,
                io_dis_uops_3_bits_is_fencei,
                io_dis_uops_3_bits_is_amo,
                io_dis_uops_3_bits_uses_ldq,
                io_dis_uops_3_bits_uses_stq,
                io_dis_uops_3_bits_ldst_val,
  input  [1:0]  io_dis_uops_3_bits_dst_rtype,
                io_dis_uops_3_bits_lrs1_rtype,
                io_dis_uops_3_bits_lrs2_rtype,
  input         io_dis_uops_3_bits_fp_val,
                io_wakeup_ports_0_valid,
  input  [6:0]  io_wakeup_ports_0_bits_pdst,
  input         io_wakeup_ports_1_valid,
  input  [6:0]  io_wakeup_ports_1_bits_pdst,
  input         io_wakeup_ports_2_valid,
  input  [6:0]  io_wakeup_ports_2_bits_pdst,
  input         io_wakeup_ports_3_valid,
  input  [6:0]  io_wakeup_ports_3_bits_pdst,
  input         io_wakeup_ports_4_valid,
  input  [6:0]  io_wakeup_ports_4_bits_pdst,
  input         io_wakeup_ports_5_valid,
  input  [6:0]  io_wakeup_ports_5_bits_pdst,
  input         io_wakeup_ports_6_valid,
  input  [6:0]  io_wakeup_ports_6_bits_pdst,
  input         io_wakeup_ports_7_valid,
  input  [6:0]  io_wakeup_ports_7_bits_pdst,
  input         io_wakeup_ports_8_valid,
  input  [6:0]  io_wakeup_ports_8_bits_pdst,
  input         io_wakeup_ports_9_valid,
  input  [6:0]  io_wakeup_ports_9_bits_pdst,
  input         io_spec_ld_wakeup_0_valid,
  input  [6:0]  io_spec_ld_wakeup_0_bits,
  input         io_spec_ld_wakeup_1_valid,
  input  [6:0]  io_spec_ld_wakeup_1_bits,
  input  [9:0]  io_fu_types_0,
                io_fu_types_2,
                io_fu_types_3,
  input  [19:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input         io_flush_pipeline,
                io_ld_miss,
  output        io_dis_uops_0_ready,
                io_dis_uops_1_ready,
                io_dis_uops_2_ready,
                io_dis_uops_3_ready,
                io_iss_valids_0,
                io_iss_valids_1,
                io_iss_valids_2,
                io_iss_valids_3,
  output [6:0]  io_iss_uops_0_uopc,
  output        io_iss_uops_0_is_rvc,
  output [9:0]  io_iss_uops_0_fu_code,
  output        io_iss_uops_0_iw_p1_poisoned,
                io_iss_uops_0_iw_p2_poisoned,
                io_iss_uops_0_is_br,
                io_iss_uops_0_is_jalr,
                io_iss_uops_0_is_jal,
                io_iss_uops_0_is_sfb,
  output [19:0] io_iss_uops_0_br_mask,
  output [4:0]  io_iss_uops_0_br_tag,
  output [5:0]  io_iss_uops_0_ftq_idx,
  output        io_iss_uops_0_edge_inst,
  output [5:0]  io_iss_uops_0_pc_lob,
  output        io_iss_uops_0_taken,
  output [19:0] io_iss_uops_0_imm_packed,
  output [6:0]  io_iss_uops_0_rob_idx,
  output [4:0]  io_iss_uops_0_ldq_idx,
                io_iss_uops_0_stq_idx,
  output [6:0]  io_iss_uops_0_pdst,
                io_iss_uops_0_prs1,
                io_iss_uops_0_prs2,
  output        io_iss_uops_0_bypassable,
  output [4:0]  io_iss_uops_0_mem_cmd,
  output        io_iss_uops_0_is_amo,
                io_iss_uops_0_uses_stq,
                io_iss_uops_0_ldst_val,
  output [1:0]  io_iss_uops_0_dst_rtype,
                io_iss_uops_0_lrs1_rtype,
                io_iss_uops_0_lrs2_rtype,
  output        io_iss_uops_0_fp_val,
  output [6:0]  io_iss_uops_1_uopc,
  output        io_iss_uops_1_is_rvc,
  output [9:0]  io_iss_uops_1_fu_code,
  output        io_iss_uops_1_iw_p1_poisoned,
                io_iss_uops_1_iw_p2_poisoned,
                io_iss_uops_1_is_br,
                io_iss_uops_1_is_jalr,
                io_iss_uops_1_is_jal,
                io_iss_uops_1_is_sfb,
  output [19:0] io_iss_uops_1_br_mask,
  output [4:0]  io_iss_uops_1_br_tag,
  output [5:0]  io_iss_uops_1_ftq_idx,
  output        io_iss_uops_1_edge_inst,
  output [5:0]  io_iss_uops_1_pc_lob,
  output        io_iss_uops_1_taken,
  output [19:0] io_iss_uops_1_imm_packed,
  output [6:0]  io_iss_uops_1_rob_idx,
  output [4:0]  io_iss_uops_1_ldq_idx,
                io_iss_uops_1_stq_idx,
  output [6:0]  io_iss_uops_1_pdst,
                io_iss_uops_1_prs1,
                io_iss_uops_1_prs2,
  output        io_iss_uops_1_bypassable,
  output [4:0]  io_iss_uops_1_mem_cmd,
  output        io_iss_uops_1_is_amo,
                io_iss_uops_1_uses_stq,
                io_iss_uops_1_ldst_val,
  output [1:0]  io_iss_uops_1_dst_rtype,
                io_iss_uops_1_lrs1_rtype,
                io_iss_uops_1_lrs2_rtype,
  output [6:0]  io_iss_uops_2_uopc,
  output        io_iss_uops_2_is_rvc,
  output [9:0]  io_iss_uops_2_fu_code,
  output        io_iss_uops_2_iw_p1_poisoned,
                io_iss_uops_2_iw_p2_poisoned,
                io_iss_uops_2_is_br,
                io_iss_uops_2_is_jalr,
                io_iss_uops_2_is_jal,
                io_iss_uops_2_is_sfb,
  output [19:0] io_iss_uops_2_br_mask,
  output [4:0]  io_iss_uops_2_br_tag,
  output [5:0]  io_iss_uops_2_ftq_idx,
  output        io_iss_uops_2_edge_inst,
  output [5:0]  io_iss_uops_2_pc_lob,
  output        io_iss_uops_2_taken,
  output [19:0] io_iss_uops_2_imm_packed,
  output [6:0]  io_iss_uops_2_rob_idx,
  output [4:0]  io_iss_uops_2_ldq_idx,
                io_iss_uops_2_stq_idx,
  output [6:0]  io_iss_uops_2_pdst,
                io_iss_uops_2_prs1,
                io_iss_uops_2_prs2,
  output        io_iss_uops_2_bypassable,
  output [4:0]  io_iss_uops_2_mem_cmd,
  output        io_iss_uops_2_is_amo,
                io_iss_uops_2_uses_stq,
                io_iss_uops_2_ldst_val,
  output [1:0]  io_iss_uops_2_dst_rtype,
                io_iss_uops_2_lrs1_rtype,
                io_iss_uops_2_lrs2_rtype,
  output [6:0]  io_iss_uops_3_uopc,
  output        io_iss_uops_3_is_rvc,
  output [9:0]  io_iss_uops_3_fu_code,
  output        io_iss_uops_3_iw_p1_poisoned,
                io_iss_uops_3_iw_p2_poisoned,
                io_iss_uops_3_is_br,
                io_iss_uops_3_is_jalr,
                io_iss_uops_3_is_jal,
                io_iss_uops_3_is_sfb,
  output [19:0] io_iss_uops_3_br_mask,
  output [4:0]  io_iss_uops_3_br_tag,
  output [5:0]  io_iss_uops_3_ftq_idx,
  output        io_iss_uops_3_edge_inst,
  output [5:0]  io_iss_uops_3_pc_lob,
  output        io_iss_uops_3_taken,
  output [19:0] io_iss_uops_3_imm_packed,
  output [6:0]  io_iss_uops_3_rob_idx,
  output [4:0]  io_iss_uops_3_ldq_idx,
                io_iss_uops_3_stq_idx,
  output [6:0]  io_iss_uops_3_pdst,
                io_iss_uops_3_prs1,
                io_iss_uops_3_prs2,
  output        io_iss_uops_3_bypassable,
  output [4:0]  io_iss_uops_3_mem_cmd,
  output        io_iss_uops_3_is_amo,
                io_iss_uops_3_uses_stq,
                io_iss_uops_3_ldst_val,
  output [1:0]  io_iss_uops_3_dst_rtype,
                io_iss_uops_3_lrs1_rtype,
                io_iss_uops_3_lrs2_rtype
);

  wire [3:0]  _GEN_97;
  wire [3:0]  _GEN_95;
  wire [3:0]  _GEN_93;
  wire [3:0]  _GEN_91;
  wire [3:0]  _GEN_89;
  wire [3:0]  _GEN_87;
  wire [3:0]  _GEN_85;
  wire [3:0]  _GEN_83;
  wire [3:0]  _GEN_81;
  wire [3:0]  _GEN_79;
  wire [3:0]  _GEN_77;
  wire [3:0]  _GEN_75;
  wire [3:0]  _GEN_73;
  wire [3:0]  _GEN_71;
  wire [3:0]  _GEN_69;
  wire [3:0]  _GEN_67;
  wire [3:0]  _GEN_65;
  wire [3:0]  _GEN_63;
  wire [3:0]  _GEN_61;
  wire [3:0]  _GEN_59;
  wire [3:0]  _GEN_57;
  wire [3:0]  _GEN_55;
  wire [3:0]  _GEN_53;
  wire [3:0]  _GEN_51;
  wire [3:0]  _GEN_49;
  wire [3:0]  _GEN_47;
  wire [3:0]  _GEN_45;
  wire [3:0]  _GEN_43;
  wire [3:0]  _GEN_41;
  wire [3:0]  _GEN_39;
  wire [3:0]  _GEN_37;
  wire [3:0]  _GEN_35;
  wire [3:0]  _GEN_33;
  wire [3:0]  _GEN_31;
  wire [3:0]  _GEN_29;
  wire [3:0]  _GEN_27;
  wire [3:0]  _GEN_25;
  wire [1:0]  _GEN_23_1to0;
  wire        _slots_39_io_valid;
  wire        _slots_39_io_will_be_valid;
  wire        _slots_39_io_request;
  wire [6:0]  _slots_39_io_out_uop_uopc;
  wire        _slots_39_io_out_uop_is_rvc;
  wire [9:0]  _slots_39_io_out_uop_fu_code;
  wire [1:0]  _slots_39_io_out_uop_iw_state;
  wire        _slots_39_io_out_uop_iw_p1_poisoned;
  wire        _slots_39_io_out_uop_iw_p2_poisoned;
  wire        _slots_39_io_out_uop_is_br;
  wire        _slots_39_io_out_uop_is_jalr;
  wire        _slots_39_io_out_uop_is_jal;
  wire        _slots_39_io_out_uop_is_sfb;
  wire [19:0] _slots_39_io_out_uop_br_mask;
  wire [4:0]  _slots_39_io_out_uop_br_tag;
  wire [5:0]  _slots_39_io_out_uop_ftq_idx;
  wire        _slots_39_io_out_uop_edge_inst;
  wire [5:0]  _slots_39_io_out_uop_pc_lob;
  wire        _slots_39_io_out_uop_taken;
  wire [19:0] _slots_39_io_out_uop_imm_packed;
  wire [6:0]  _slots_39_io_out_uop_rob_idx;
  wire [4:0]  _slots_39_io_out_uop_ldq_idx;
  wire [4:0]  _slots_39_io_out_uop_stq_idx;
  wire [6:0]  _slots_39_io_out_uop_pdst;
  wire [6:0]  _slots_39_io_out_uop_prs1;
  wire [6:0]  _slots_39_io_out_uop_prs2;
  wire [6:0]  _slots_39_io_out_uop_prs3;
  wire        _slots_39_io_out_uop_prs1_busy;
  wire        _slots_39_io_out_uop_prs2_busy;
  wire        _slots_39_io_out_uop_prs3_busy;
  wire        _slots_39_io_out_uop_ppred_busy;
  wire        _slots_39_io_out_uop_bypassable;
  wire [4:0]  _slots_39_io_out_uop_mem_cmd;
  wire [1:0]  _slots_39_io_out_uop_mem_size;
  wire        _slots_39_io_out_uop_mem_signed;
  wire        _slots_39_io_out_uop_is_fence;
  wire        _slots_39_io_out_uop_is_amo;
  wire        _slots_39_io_out_uop_uses_ldq;
  wire        _slots_39_io_out_uop_uses_stq;
  wire        _slots_39_io_out_uop_ldst_val;
  wire [1:0]  _slots_39_io_out_uop_dst_rtype;
  wire [1:0]  _slots_39_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_39_io_out_uop_lrs2_rtype;
  wire        _slots_39_io_out_uop_fp_val;
  wire [6:0]  _slots_39_io_uop_uopc;
  wire        _slots_39_io_uop_is_rvc;
  wire [9:0]  _slots_39_io_uop_fu_code;
  wire        _slots_39_io_uop_iw_p1_poisoned;
  wire        _slots_39_io_uop_iw_p2_poisoned;
  wire        _slots_39_io_uop_is_br;
  wire        _slots_39_io_uop_is_jalr;
  wire        _slots_39_io_uop_is_jal;
  wire        _slots_39_io_uop_is_sfb;
  wire [19:0] _slots_39_io_uop_br_mask;
  wire [4:0]  _slots_39_io_uop_br_tag;
  wire [5:0]  _slots_39_io_uop_ftq_idx;
  wire        _slots_39_io_uop_edge_inst;
  wire [5:0]  _slots_39_io_uop_pc_lob;
  wire        _slots_39_io_uop_taken;
  wire [19:0] _slots_39_io_uop_imm_packed;
  wire [6:0]  _slots_39_io_uop_rob_idx;
  wire [4:0]  _slots_39_io_uop_ldq_idx;
  wire [4:0]  _slots_39_io_uop_stq_idx;
  wire [6:0]  _slots_39_io_uop_pdst;
  wire [6:0]  _slots_39_io_uop_prs1;
  wire [6:0]  _slots_39_io_uop_prs2;
  wire        _slots_39_io_uop_bypassable;
  wire [4:0]  _slots_39_io_uop_mem_cmd;
  wire        _slots_39_io_uop_is_amo;
  wire        _slots_39_io_uop_uses_stq;
  wire        _slots_39_io_uop_ldst_val;
  wire [1:0]  _slots_39_io_uop_dst_rtype;
  wire [1:0]  _slots_39_io_uop_lrs1_rtype;
  wire [1:0]  _slots_39_io_uop_lrs2_rtype;
  wire        _slots_39_io_uop_fp_val;
  wire        _slots_38_io_valid;
  wire        _slots_38_io_will_be_valid;
  wire        _slots_38_io_request;
  wire [6:0]  _slots_38_io_out_uop_uopc;
  wire        _slots_38_io_out_uop_is_rvc;
  wire [9:0]  _slots_38_io_out_uop_fu_code;
  wire [1:0]  _slots_38_io_out_uop_iw_state;
  wire        _slots_38_io_out_uop_iw_p1_poisoned;
  wire        _slots_38_io_out_uop_iw_p2_poisoned;
  wire        _slots_38_io_out_uop_is_br;
  wire        _slots_38_io_out_uop_is_jalr;
  wire        _slots_38_io_out_uop_is_jal;
  wire        _slots_38_io_out_uop_is_sfb;
  wire [19:0] _slots_38_io_out_uop_br_mask;
  wire [4:0]  _slots_38_io_out_uop_br_tag;
  wire [5:0]  _slots_38_io_out_uop_ftq_idx;
  wire        _slots_38_io_out_uop_edge_inst;
  wire [5:0]  _slots_38_io_out_uop_pc_lob;
  wire        _slots_38_io_out_uop_taken;
  wire [19:0] _slots_38_io_out_uop_imm_packed;
  wire [6:0]  _slots_38_io_out_uop_rob_idx;
  wire [4:0]  _slots_38_io_out_uop_ldq_idx;
  wire [4:0]  _slots_38_io_out_uop_stq_idx;
  wire [6:0]  _slots_38_io_out_uop_pdst;
  wire [6:0]  _slots_38_io_out_uop_prs1;
  wire [6:0]  _slots_38_io_out_uop_prs2;
  wire [6:0]  _slots_38_io_out_uop_prs3;
  wire        _slots_38_io_out_uop_prs1_busy;
  wire        _slots_38_io_out_uop_prs2_busy;
  wire        _slots_38_io_out_uop_prs3_busy;
  wire        _slots_38_io_out_uop_ppred_busy;
  wire        _slots_38_io_out_uop_bypassable;
  wire [4:0]  _slots_38_io_out_uop_mem_cmd;
  wire [1:0]  _slots_38_io_out_uop_mem_size;
  wire        _slots_38_io_out_uop_mem_signed;
  wire        _slots_38_io_out_uop_is_fence;
  wire        _slots_38_io_out_uop_is_amo;
  wire        _slots_38_io_out_uop_uses_ldq;
  wire        _slots_38_io_out_uop_uses_stq;
  wire        _slots_38_io_out_uop_ldst_val;
  wire [1:0]  _slots_38_io_out_uop_dst_rtype;
  wire [1:0]  _slots_38_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_38_io_out_uop_lrs2_rtype;
  wire        _slots_38_io_out_uop_fp_val;
  wire [6:0]  _slots_38_io_uop_uopc;
  wire        _slots_38_io_uop_is_rvc;
  wire [9:0]  _slots_38_io_uop_fu_code;
  wire        _slots_38_io_uop_iw_p1_poisoned;
  wire        _slots_38_io_uop_iw_p2_poisoned;
  wire        _slots_38_io_uop_is_br;
  wire        _slots_38_io_uop_is_jalr;
  wire        _slots_38_io_uop_is_jal;
  wire        _slots_38_io_uop_is_sfb;
  wire [19:0] _slots_38_io_uop_br_mask;
  wire [4:0]  _slots_38_io_uop_br_tag;
  wire [5:0]  _slots_38_io_uop_ftq_idx;
  wire        _slots_38_io_uop_edge_inst;
  wire [5:0]  _slots_38_io_uop_pc_lob;
  wire        _slots_38_io_uop_taken;
  wire [19:0] _slots_38_io_uop_imm_packed;
  wire [6:0]  _slots_38_io_uop_rob_idx;
  wire [4:0]  _slots_38_io_uop_ldq_idx;
  wire [4:0]  _slots_38_io_uop_stq_idx;
  wire [6:0]  _slots_38_io_uop_pdst;
  wire [6:0]  _slots_38_io_uop_prs1;
  wire [6:0]  _slots_38_io_uop_prs2;
  wire        _slots_38_io_uop_bypassable;
  wire [4:0]  _slots_38_io_uop_mem_cmd;
  wire        _slots_38_io_uop_is_amo;
  wire        _slots_38_io_uop_uses_stq;
  wire        _slots_38_io_uop_ldst_val;
  wire [1:0]  _slots_38_io_uop_dst_rtype;
  wire [1:0]  _slots_38_io_uop_lrs1_rtype;
  wire [1:0]  _slots_38_io_uop_lrs2_rtype;
  wire        _slots_38_io_uop_fp_val;
  wire        _slots_37_io_valid;
  wire        _slots_37_io_will_be_valid;
  wire        _slots_37_io_request;
  wire [6:0]  _slots_37_io_out_uop_uopc;
  wire        _slots_37_io_out_uop_is_rvc;
  wire [9:0]  _slots_37_io_out_uop_fu_code;
  wire [1:0]  _slots_37_io_out_uop_iw_state;
  wire        _slots_37_io_out_uop_iw_p1_poisoned;
  wire        _slots_37_io_out_uop_iw_p2_poisoned;
  wire        _slots_37_io_out_uop_is_br;
  wire        _slots_37_io_out_uop_is_jalr;
  wire        _slots_37_io_out_uop_is_jal;
  wire        _slots_37_io_out_uop_is_sfb;
  wire [19:0] _slots_37_io_out_uop_br_mask;
  wire [4:0]  _slots_37_io_out_uop_br_tag;
  wire [5:0]  _slots_37_io_out_uop_ftq_idx;
  wire        _slots_37_io_out_uop_edge_inst;
  wire [5:0]  _slots_37_io_out_uop_pc_lob;
  wire        _slots_37_io_out_uop_taken;
  wire [19:0] _slots_37_io_out_uop_imm_packed;
  wire [6:0]  _slots_37_io_out_uop_rob_idx;
  wire [4:0]  _slots_37_io_out_uop_ldq_idx;
  wire [4:0]  _slots_37_io_out_uop_stq_idx;
  wire [6:0]  _slots_37_io_out_uop_pdst;
  wire [6:0]  _slots_37_io_out_uop_prs1;
  wire [6:0]  _slots_37_io_out_uop_prs2;
  wire [6:0]  _slots_37_io_out_uop_prs3;
  wire        _slots_37_io_out_uop_prs1_busy;
  wire        _slots_37_io_out_uop_prs2_busy;
  wire        _slots_37_io_out_uop_prs3_busy;
  wire        _slots_37_io_out_uop_ppred_busy;
  wire        _slots_37_io_out_uop_bypassable;
  wire [4:0]  _slots_37_io_out_uop_mem_cmd;
  wire [1:0]  _slots_37_io_out_uop_mem_size;
  wire        _slots_37_io_out_uop_mem_signed;
  wire        _slots_37_io_out_uop_is_fence;
  wire        _slots_37_io_out_uop_is_amo;
  wire        _slots_37_io_out_uop_uses_ldq;
  wire        _slots_37_io_out_uop_uses_stq;
  wire        _slots_37_io_out_uop_ldst_val;
  wire [1:0]  _slots_37_io_out_uop_dst_rtype;
  wire [1:0]  _slots_37_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_37_io_out_uop_lrs2_rtype;
  wire        _slots_37_io_out_uop_fp_val;
  wire [6:0]  _slots_37_io_uop_uopc;
  wire        _slots_37_io_uop_is_rvc;
  wire [9:0]  _slots_37_io_uop_fu_code;
  wire        _slots_37_io_uop_iw_p1_poisoned;
  wire        _slots_37_io_uop_iw_p2_poisoned;
  wire        _slots_37_io_uop_is_br;
  wire        _slots_37_io_uop_is_jalr;
  wire        _slots_37_io_uop_is_jal;
  wire        _slots_37_io_uop_is_sfb;
  wire [19:0] _slots_37_io_uop_br_mask;
  wire [4:0]  _slots_37_io_uop_br_tag;
  wire [5:0]  _slots_37_io_uop_ftq_idx;
  wire        _slots_37_io_uop_edge_inst;
  wire [5:0]  _slots_37_io_uop_pc_lob;
  wire        _slots_37_io_uop_taken;
  wire [19:0] _slots_37_io_uop_imm_packed;
  wire [6:0]  _slots_37_io_uop_rob_idx;
  wire [4:0]  _slots_37_io_uop_ldq_idx;
  wire [4:0]  _slots_37_io_uop_stq_idx;
  wire [6:0]  _slots_37_io_uop_pdst;
  wire [6:0]  _slots_37_io_uop_prs1;
  wire [6:0]  _slots_37_io_uop_prs2;
  wire        _slots_37_io_uop_bypassable;
  wire [4:0]  _slots_37_io_uop_mem_cmd;
  wire        _slots_37_io_uop_is_amo;
  wire        _slots_37_io_uop_uses_stq;
  wire        _slots_37_io_uop_ldst_val;
  wire [1:0]  _slots_37_io_uop_dst_rtype;
  wire [1:0]  _slots_37_io_uop_lrs1_rtype;
  wire [1:0]  _slots_37_io_uop_lrs2_rtype;
  wire        _slots_37_io_uop_fp_val;
  wire        _slots_36_io_valid;
  wire        _slots_36_io_will_be_valid;
  wire        _slots_36_io_request;
  wire [6:0]  _slots_36_io_out_uop_uopc;
  wire        _slots_36_io_out_uop_is_rvc;
  wire [9:0]  _slots_36_io_out_uop_fu_code;
  wire [1:0]  _slots_36_io_out_uop_iw_state;
  wire        _slots_36_io_out_uop_iw_p1_poisoned;
  wire        _slots_36_io_out_uop_iw_p2_poisoned;
  wire        _slots_36_io_out_uop_is_br;
  wire        _slots_36_io_out_uop_is_jalr;
  wire        _slots_36_io_out_uop_is_jal;
  wire        _slots_36_io_out_uop_is_sfb;
  wire [19:0] _slots_36_io_out_uop_br_mask;
  wire [4:0]  _slots_36_io_out_uop_br_tag;
  wire [5:0]  _slots_36_io_out_uop_ftq_idx;
  wire        _slots_36_io_out_uop_edge_inst;
  wire [5:0]  _slots_36_io_out_uop_pc_lob;
  wire        _slots_36_io_out_uop_taken;
  wire [19:0] _slots_36_io_out_uop_imm_packed;
  wire [6:0]  _slots_36_io_out_uop_rob_idx;
  wire [4:0]  _slots_36_io_out_uop_ldq_idx;
  wire [4:0]  _slots_36_io_out_uop_stq_idx;
  wire [6:0]  _slots_36_io_out_uop_pdst;
  wire [6:0]  _slots_36_io_out_uop_prs1;
  wire [6:0]  _slots_36_io_out_uop_prs2;
  wire [6:0]  _slots_36_io_out_uop_prs3;
  wire        _slots_36_io_out_uop_prs1_busy;
  wire        _slots_36_io_out_uop_prs2_busy;
  wire        _slots_36_io_out_uop_prs3_busy;
  wire        _slots_36_io_out_uop_ppred_busy;
  wire        _slots_36_io_out_uop_bypassable;
  wire [4:0]  _slots_36_io_out_uop_mem_cmd;
  wire [1:0]  _slots_36_io_out_uop_mem_size;
  wire        _slots_36_io_out_uop_mem_signed;
  wire        _slots_36_io_out_uop_is_fence;
  wire        _slots_36_io_out_uop_is_amo;
  wire        _slots_36_io_out_uop_uses_ldq;
  wire        _slots_36_io_out_uop_uses_stq;
  wire        _slots_36_io_out_uop_ldst_val;
  wire [1:0]  _slots_36_io_out_uop_dst_rtype;
  wire [1:0]  _slots_36_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_36_io_out_uop_lrs2_rtype;
  wire        _slots_36_io_out_uop_fp_val;
  wire [6:0]  _slots_36_io_uop_uopc;
  wire        _slots_36_io_uop_is_rvc;
  wire [9:0]  _slots_36_io_uop_fu_code;
  wire        _slots_36_io_uop_iw_p1_poisoned;
  wire        _slots_36_io_uop_iw_p2_poisoned;
  wire        _slots_36_io_uop_is_br;
  wire        _slots_36_io_uop_is_jalr;
  wire        _slots_36_io_uop_is_jal;
  wire        _slots_36_io_uop_is_sfb;
  wire [19:0] _slots_36_io_uop_br_mask;
  wire [4:0]  _slots_36_io_uop_br_tag;
  wire [5:0]  _slots_36_io_uop_ftq_idx;
  wire        _slots_36_io_uop_edge_inst;
  wire [5:0]  _slots_36_io_uop_pc_lob;
  wire        _slots_36_io_uop_taken;
  wire [19:0] _slots_36_io_uop_imm_packed;
  wire [6:0]  _slots_36_io_uop_rob_idx;
  wire [4:0]  _slots_36_io_uop_ldq_idx;
  wire [4:0]  _slots_36_io_uop_stq_idx;
  wire [6:0]  _slots_36_io_uop_pdst;
  wire [6:0]  _slots_36_io_uop_prs1;
  wire [6:0]  _slots_36_io_uop_prs2;
  wire        _slots_36_io_uop_bypassable;
  wire [4:0]  _slots_36_io_uop_mem_cmd;
  wire        _slots_36_io_uop_is_amo;
  wire        _slots_36_io_uop_uses_stq;
  wire        _slots_36_io_uop_ldst_val;
  wire [1:0]  _slots_36_io_uop_dst_rtype;
  wire [1:0]  _slots_36_io_uop_lrs1_rtype;
  wire [1:0]  _slots_36_io_uop_lrs2_rtype;
  wire        _slots_36_io_uop_fp_val;
  wire        _slots_35_io_valid;
  wire        _slots_35_io_will_be_valid;
  wire        _slots_35_io_request;
  wire [6:0]  _slots_35_io_out_uop_uopc;
  wire        _slots_35_io_out_uop_is_rvc;
  wire [9:0]  _slots_35_io_out_uop_fu_code;
  wire [1:0]  _slots_35_io_out_uop_iw_state;
  wire        _slots_35_io_out_uop_iw_p1_poisoned;
  wire        _slots_35_io_out_uop_iw_p2_poisoned;
  wire        _slots_35_io_out_uop_is_br;
  wire        _slots_35_io_out_uop_is_jalr;
  wire        _slots_35_io_out_uop_is_jal;
  wire        _slots_35_io_out_uop_is_sfb;
  wire [19:0] _slots_35_io_out_uop_br_mask;
  wire [4:0]  _slots_35_io_out_uop_br_tag;
  wire [5:0]  _slots_35_io_out_uop_ftq_idx;
  wire        _slots_35_io_out_uop_edge_inst;
  wire [5:0]  _slots_35_io_out_uop_pc_lob;
  wire        _slots_35_io_out_uop_taken;
  wire [19:0] _slots_35_io_out_uop_imm_packed;
  wire [6:0]  _slots_35_io_out_uop_rob_idx;
  wire [4:0]  _slots_35_io_out_uop_ldq_idx;
  wire [4:0]  _slots_35_io_out_uop_stq_idx;
  wire [6:0]  _slots_35_io_out_uop_pdst;
  wire [6:0]  _slots_35_io_out_uop_prs1;
  wire [6:0]  _slots_35_io_out_uop_prs2;
  wire [6:0]  _slots_35_io_out_uop_prs3;
  wire        _slots_35_io_out_uop_prs1_busy;
  wire        _slots_35_io_out_uop_prs2_busy;
  wire        _slots_35_io_out_uop_prs3_busy;
  wire        _slots_35_io_out_uop_ppred_busy;
  wire        _slots_35_io_out_uop_bypassable;
  wire [4:0]  _slots_35_io_out_uop_mem_cmd;
  wire [1:0]  _slots_35_io_out_uop_mem_size;
  wire        _slots_35_io_out_uop_mem_signed;
  wire        _slots_35_io_out_uop_is_fence;
  wire        _slots_35_io_out_uop_is_amo;
  wire        _slots_35_io_out_uop_uses_ldq;
  wire        _slots_35_io_out_uop_uses_stq;
  wire        _slots_35_io_out_uop_ldst_val;
  wire [1:0]  _slots_35_io_out_uop_dst_rtype;
  wire [1:0]  _slots_35_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_35_io_out_uop_lrs2_rtype;
  wire        _slots_35_io_out_uop_fp_val;
  wire [6:0]  _slots_35_io_uop_uopc;
  wire        _slots_35_io_uop_is_rvc;
  wire [9:0]  _slots_35_io_uop_fu_code;
  wire        _slots_35_io_uop_iw_p1_poisoned;
  wire        _slots_35_io_uop_iw_p2_poisoned;
  wire        _slots_35_io_uop_is_br;
  wire        _slots_35_io_uop_is_jalr;
  wire        _slots_35_io_uop_is_jal;
  wire        _slots_35_io_uop_is_sfb;
  wire [19:0] _slots_35_io_uop_br_mask;
  wire [4:0]  _slots_35_io_uop_br_tag;
  wire [5:0]  _slots_35_io_uop_ftq_idx;
  wire        _slots_35_io_uop_edge_inst;
  wire [5:0]  _slots_35_io_uop_pc_lob;
  wire        _slots_35_io_uop_taken;
  wire [19:0] _slots_35_io_uop_imm_packed;
  wire [6:0]  _slots_35_io_uop_rob_idx;
  wire [4:0]  _slots_35_io_uop_ldq_idx;
  wire [4:0]  _slots_35_io_uop_stq_idx;
  wire [6:0]  _slots_35_io_uop_pdst;
  wire [6:0]  _slots_35_io_uop_prs1;
  wire [6:0]  _slots_35_io_uop_prs2;
  wire        _slots_35_io_uop_bypassable;
  wire [4:0]  _slots_35_io_uop_mem_cmd;
  wire        _slots_35_io_uop_is_amo;
  wire        _slots_35_io_uop_uses_stq;
  wire        _slots_35_io_uop_ldst_val;
  wire [1:0]  _slots_35_io_uop_dst_rtype;
  wire [1:0]  _slots_35_io_uop_lrs1_rtype;
  wire [1:0]  _slots_35_io_uop_lrs2_rtype;
  wire        _slots_35_io_uop_fp_val;
  wire        _slots_34_io_valid;
  wire        _slots_34_io_will_be_valid;
  wire        _slots_34_io_request;
  wire [6:0]  _slots_34_io_out_uop_uopc;
  wire        _slots_34_io_out_uop_is_rvc;
  wire [9:0]  _slots_34_io_out_uop_fu_code;
  wire [1:0]  _slots_34_io_out_uop_iw_state;
  wire        _slots_34_io_out_uop_iw_p1_poisoned;
  wire        _slots_34_io_out_uop_iw_p2_poisoned;
  wire        _slots_34_io_out_uop_is_br;
  wire        _slots_34_io_out_uop_is_jalr;
  wire        _slots_34_io_out_uop_is_jal;
  wire        _slots_34_io_out_uop_is_sfb;
  wire [19:0] _slots_34_io_out_uop_br_mask;
  wire [4:0]  _slots_34_io_out_uop_br_tag;
  wire [5:0]  _slots_34_io_out_uop_ftq_idx;
  wire        _slots_34_io_out_uop_edge_inst;
  wire [5:0]  _slots_34_io_out_uop_pc_lob;
  wire        _slots_34_io_out_uop_taken;
  wire [19:0] _slots_34_io_out_uop_imm_packed;
  wire [6:0]  _slots_34_io_out_uop_rob_idx;
  wire [4:0]  _slots_34_io_out_uop_ldq_idx;
  wire [4:0]  _slots_34_io_out_uop_stq_idx;
  wire [6:0]  _slots_34_io_out_uop_pdst;
  wire [6:0]  _slots_34_io_out_uop_prs1;
  wire [6:0]  _slots_34_io_out_uop_prs2;
  wire [6:0]  _slots_34_io_out_uop_prs3;
  wire        _slots_34_io_out_uop_prs1_busy;
  wire        _slots_34_io_out_uop_prs2_busy;
  wire        _slots_34_io_out_uop_prs3_busy;
  wire        _slots_34_io_out_uop_ppred_busy;
  wire        _slots_34_io_out_uop_bypassable;
  wire [4:0]  _slots_34_io_out_uop_mem_cmd;
  wire [1:0]  _slots_34_io_out_uop_mem_size;
  wire        _slots_34_io_out_uop_mem_signed;
  wire        _slots_34_io_out_uop_is_fence;
  wire        _slots_34_io_out_uop_is_amo;
  wire        _slots_34_io_out_uop_uses_ldq;
  wire        _slots_34_io_out_uop_uses_stq;
  wire        _slots_34_io_out_uop_ldst_val;
  wire [1:0]  _slots_34_io_out_uop_dst_rtype;
  wire [1:0]  _slots_34_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_34_io_out_uop_lrs2_rtype;
  wire        _slots_34_io_out_uop_fp_val;
  wire [6:0]  _slots_34_io_uop_uopc;
  wire        _slots_34_io_uop_is_rvc;
  wire [9:0]  _slots_34_io_uop_fu_code;
  wire        _slots_34_io_uop_iw_p1_poisoned;
  wire        _slots_34_io_uop_iw_p2_poisoned;
  wire        _slots_34_io_uop_is_br;
  wire        _slots_34_io_uop_is_jalr;
  wire        _slots_34_io_uop_is_jal;
  wire        _slots_34_io_uop_is_sfb;
  wire [19:0] _slots_34_io_uop_br_mask;
  wire [4:0]  _slots_34_io_uop_br_tag;
  wire [5:0]  _slots_34_io_uop_ftq_idx;
  wire        _slots_34_io_uop_edge_inst;
  wire [5:0]  _slots_34_io_uop_pc_lob;
  wire        _slots_34_io_uop_taken;
  wire [19:0] _slots_34_io_uop_imm_packed;
  wire [6:0]  _slots_34_io_uop_rob_idx;
  wire [4:0]  _slots_34_io_uop_ldq_idx;
  wire [4:0]  _slots_34_io_uop_stq_idx;
  wire [6:0]  _slots_34_io_uop_pdst;
  wire [6:0]  _slots_34_io_uop_prs1;
  wire [6:0]  _slots_34_io_uop_prs2;
  wire        _slots_34_io_uop_bypassable;
  wire [4:0]  _slots_34_io_uop_mem_cmd;
  wire        _slots_34_io_uop_is_amo;
  wire        _slots_34_io_uop_uses_stq;
  wire        _slots_34_io_uop_ldst_val;
  wire [1:0]  _slots_34_io_uop_dst_rtype;
  wire [1:0]  _slots_34_io_uop_lrs1_rtype;
  wire [1:0]  _slots_34_io_uop_lrs2_rtype;
  wire        _slots_34_io_uop_fp_val;
  wire        _slots_33_io_valid;
  wire        _slots_33_io_will_be_valid;
  wire        _slots_33_io_request;
  wire [6:0]  _slots_33_io_out_uop_uopc;
  wire        _slots_33_io_out_uop_is_rvc;
  wire [9:0]  _slots_33_io_out_uop_fu_code;
  wire [1:0]  _slots_33_io_out_uop_iw_state;
  wire        _slots_33_io_out_uop_iw_p1_poisoned;
  wire        _slots_33_io_out_uop_iw_p2_poisoned;
  wire        _slots_33_io_out_uop_is_br;
  wire        _slots_33_io_out_uop_is_jalr;
  wire        _slots_33_io_out_uop_is_jal;
  wire        _slots_33_io_out_uop_is_sfb;
  wire [19:0] _slots_33_io_out_uop_br_mask;
  wire [4:0]  _slots_33_io_out_uop_br_tag;
  wire [5:0]  _slots_33_io_out_uop_ftq_idx;
  wire        _slots_33_io_out_uop_edge_inst;
  wire [5:0]  _slots_33_io_out_uop_pc_lob;
  wire        _slots_33_io_out_uop_taken;
  wire [19:0] _slots_33_io_out_uop_imm_packed;
  wire [6:0]  _slots_33_io_out_uop_rob_idx;
  wire [4:0]  _slots_33_io_out_uop_ldq_idx;
  wire [4:0]  _slots_33_io_out_uop_stq_idx;
  wire [6:0]  _slots_33_io_out_uop_pdst;
  wire [6:0]  _slots_33_io_out_uop_prs1;
  wire [6:0]  _slots_33_io_out_uop_prs2;
  wire [6:0]  _slots_33_io_out_uop_prs3;
  wire        _slots_33_io_out_uop_prs1_busy;
  wire        _slots_33_io_out_uop_prs2_busy;
  wire        _slots_33_io_out_uop_prs3_busy;
  wire        _slots_33_io_out_uop_ppred_busy;
  wire        _slots_33_io_out_uop_bypassable;
  wire [4:0]  _slots_33_io_out_uop_mem_cmd;
  wire [1:0]  _slots_33_io_out_uop_mem_size;
  wire        _slots_33_io_out_uop_mem_signed;
  wire        _slots_33_io_out_uop_is_fence;
  wire        _slots_33_io_out_uop_is_amo;
  wire        _slots_33_io_out_uop_uses_ldq;
  wire        _slots_33_io_out_uop_uses_stq;
  wire        _slots_33_io_out_uop_ldst_val;
  wire [1:0]  _slots_33_io_out_uop_dst_rtype;
  wire [1:0]  _slots_33_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_33_io_out_uop_lrs2_rtype;
  wire        _slots_33_io_out_uop_fp_val;
  wire [6:0]  _slots_33_io_uop_uopc;
  wire        _slots_33_io_uop_is_rvc;
  wire [9:0]  _slots_33_io_uop_fu_code;
  wire        _slots_33_io_uop_iw_p1_poisoned;
  wire        _slots_33_io_uop_iw_p2_poisoned;
  wire        _slots_33_io_uop_is_br;
  wire        _slots_33_io_uop_is_jalr;
  wire        _slots_33_io_uop_is_jal;
  wire        _slots_33_io_uop_is_sfb;
  wire [19:0] _slots_33_io_uop_br_mask;
  wire [4:0]  _slots_33_io_uop_br_tag;
  wire [5:0]  _slots_33_io_uop_ftq_idx;
  wire        _slots_33_io_uop_edge_inst;
  wire [5:0]  _slots_33_io_uop_pc_lob;
  wire        _slots_33_io_uop_taken;
  wire [19:0] _slots_33_io_uop_imm_packed;
  wire [6:0]  _slots_33_io_uop_rob_idx;
  wire [4:0]  _slots_33_io_uop_ldq_idx;
  wire [4:0]  _slots_33_io_uop_stq_idx;
  wire [6:0]  _slots_33_io_uop_pdst;
  wire [6:0]  _slots_33_io_uop_prs1;
  wire [6:0]  _slots_33_io_uop_prs2;
  wire        _slots_33_io_uop_bypassable;
  wire [4:0]  _slots_33_io_uop_mem_cmd;
  wire        _slots_33_io_uop_is_amo;
  wire        _slots_33_io_uop_uses_stq;
  wire        _slots_33_io_uop_ldst_val;
  wire [1:0]  _slots_33_io_uop_dst_rtype;
  wire [1:0]  _slots_33_io_uop_lrs1_rtype;
  wire [1:0]  _slots_33_io_uop_lrs2_rtype;
  wire        _slots_33_io_uop_fp_val;
  wire        _slots_32_io_valid;
  wire        _slots_32_io_will_be_valid;
  wire        _slots_32_io_request;
  wire [6:0]  _slots_32_io_out_uop_uopc;
  wire        _slots_32_io_out_uop_is_rvc;
  wire [9:0]  _slots_32_io_out_uop_fu_code;
  wire [1:0]  _slots_32_io_out_uop_iw_state;
  wire        _slots_32_io_out_uop_iw_p1_poisoned;
  wire        _slots_32_io_out_uop_iw_p2_poisoned;
  wire        _slots_32_io_out_uop_is_br;
  wire        _slots_32_io_out_uop_is_jalr;
  wire        _slots_32_io_out_uop_is_jal;
  wire        _slots_32_io_out_uop_is_sfb;
  wire [19:0] _slots_32_io_out_uop_br_mask;
  wire [4:0]  _slots_32_io_out_uop_br_tag;
  wire [5:0]  _slots_32_io_out_uop_ftq_idx;
  wire        _slots_32_io_out_uop_edge_inst;
  wire [5:0]  _slots_32_io_out_uop_pc_lob;
  wire        _slots_32_io_out_uop_taken;
  wire [19:0] _slots_32_io_out_uop_imm_packed;
  wire [6:0]  _slots_32_io_out_uop_rob_idx;
  wire [4:0]  _slots_32_io_out_uop_ldq_idx;
  wire [4:0]  _slots_32_io_out_uop_stq_idx;
  wire [6:0]  _slots_32_io_out_uop_pdst;
  wire [6:0]  _slots_32_io_out_uop_prs1;
  wire [6:0]  _slots_32_io_out_uop_prs2;
  wire [6:0]  _slots_32_io_out_uop_prs3;
  wire        _slots_32_io_out_uop_prs1_busy;
  wire        _slots_32_io_out_uop_prs2_busy;
  wire        _slots_32_io_out_uop_prs3_busy;
  wire        _slots_32_io_out_uop_ppred_busy;
  wire        _slots_32_io_out_uop_bypassable;
  wire [4:0]  _slots_32_io_out_uop_mem_cmd;
  wire [1:0]  _slots_32_io_out_uop_mem_size;
  wire        _slots_32_io_out_uop_mem_signed;
  wire        _slots_32_io_out_uop_is_fence;
  wire        _slots_32_io_out_uop_is_amo;
  wire        _slots_32_io_out_uop_uses_ldq;
  wire        _slots_32_io_out_uop_uses_stq;
  wire        _slots_32_io_out_uop_ldst_val;
  wire [1:0]  _slots_32_io_out_uop_dst_rtype;
  wire [1:0]  _slots_32_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_32_io_out_uop_lrs2_rtype;
  wire        _slots_32_io_out_uop_fp_val;
  wire [6:0]  _slots_32_io_uop_uopc;
  wire        _slots_32_io_uop_is_rvc;
  wire [9:0]  _slots_32_io_uop_fu_code;
  wire        _slots_32_io_uop_iw_p1_poisoned;
  wire        _slots_32_io_uop_iw_p2_poisoned;
  wire        _slots_32_io_uop_is_br;
  wire        _slots_32_io_uop_is_jalr;
  wire        _slots_32_io_uop_is_jal;
  wire        _slots_32_io_uop_is_sfb;
  wire [19:0] _slots_32_io_uop_br_mask;
  wire [4:0]  _slots_32_io_uop_br_tag;
  wire [5:0]  _slots_32_io_uop_ftq_idx;
  wire        _slots_32_io_uop_edge_inst;
  wire [5:0]  _slots_32_io_uop_pc_lob;
  wire        _slots_32_io_uop_taken;
  wire [19:0] _slots_32_io_uop_imm_packed;
  wire [6:0]  _slots_32_io_uop_rob_idx;
  wire [4:0]  _slots_32_io_uop_ldq_idx;
  wire [4:0]  _slots_32_io_uop_stq_idx;
  wire [6:0]  _slots_32_io_uop_pdst;
  wire [6:0]  _slots_32_io_uop_prs1;
  wire [6:0]  _slots_32_io_uop_prs2;
  wire        _slots_32_io_uop_bypassable;
  wire [4:0]  _slots_32_io_uop_mem_cmd;
  wire        _slots_32_io_uop_is_amo;
  wire        _slots_32_io_uop_uses_stq;
  wire        _slots_32_io_uop_ldst_val;
  wire [1:0]  _slots_32_io_uop_dst_rtype;
  wire [1:0]  _slots_32_io_uop_lrs1_rtype;
  wire [1:0]  _slots_32_io_uop_lrs2_rtype;
  wire        _slots_32_io_uop_fp_val;
  wire        _slots_31_io_valid;
  wire        _slots_31_io_will_be_valid;
  wire        _slots_31_io_request;
  wire [6:0]  _slots_31_io_out_uop_uopc;
  wire        _slots_31_io_out_uop_is_rvc;
  wire [9:0]  _slots_31_io_out_uop_fu_code;
  wire [1:0]  _slots_31_io_out_uop_iw_state;
  wire        _slots_31_io_out_uop_iw_p1_poisoned;
  wire        _slots_31_io_out_uop_iw_p2_poisoned;
  wire        _slots_31_io_out_uop_is_br;
  wire        _slots_31_io_out_uop_is_jalr;
  wire        _slots_31_io_out_uop_is_jal;
  wire        _slots_31_io_out_uop_is_sfb;
  wire [19:0] _slots_31_io_out_uop_br_mask;
  wire [4:0]  _slots_31_io_out_uop_br_tag;
  wire [5:0]  _slots_31_io_out_uop_ftq_idx;
  wire        _slots_31_io_out_uop_edge_inst;
  wire [5:0]  _slots_31_io_out_uop_pc_lob;
  wire        _slots_31_io_out_uop_taken;
  wire [19:0] _slots_31_io_out_uop_imm_packed;
  wire [6:0]  _slots_31_io_out_uop_rob_idx;
  wire [4:0]  _slots_31_io_out_uop_ldq_idx;
  wire [4:0]  _slots_31_io_out_uop_stq_idx;
  wire [6:0]  _slots_31_io_out_uop_pdst;
  wire [6:0]  _slots_31_io_out_uop_prs1;
  wire [6:0]  _slots_31_io_out_uop_prs2;
  wire [6:0]  _slots_31_io_out_uop_prs3;
  wire        _slots_31_io_out_uop_prs1_busy;
  wire        _slots_31_io_out_uop_prs2_busy;
  wire        _slots_31_io_out_uop_prs3_busy;
  wire        _slots_31_io_out_uop_ppred_busy;
  wire        _slots_31_io_out_uop_bypassable;
  wire [4:0]  _slots_31_io_out_uop_mem_cmd;
  wire [1:0]  _slots_31_io_out_uop_mem_size;
  wire        _slots_31_io_out_uop_mem_signed;
  wire        _slots_31_io_out_uop_is_fence;
  wire        _slots_31_io_out_uop_is_amo;
  wire        _slots_31_io_out_uop_uses_ldq;
  wire        _slots_31_io_out_uop_uses_stq;
  wire        _slots_31_io_out_uop_ldst_val;
  wire [1:0]  _slots_31_io_out_uop_dst_rtype;
  wire [1:0]  _slots_31_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_31_io_out_uop_lrs2_rtype;
  wire        _slots_31_io_out_uop_fp_val;
  wire [6:0]  _slots_31_io_uop_uopc;
  wire        _slots_31_io_uop_is_rvc;
  wire [9:0]  _slots_31_io_uop_fu_code;
  wire        _slots_31_io_uop_iw_p1_poisoned;
  wire        _slots_31_io_uop_iw_p2_poisoned;
  wire        _slots_31_io_uop_is_br;
  wire        _slots_31_io_uop_is_jalr;
  wire        _slots_31_io_uop_is_jal;
  wire        _slots_31_io_uop_is_sfb;
  wire [19:0] _slots_31_io_uop_br_mask;
  wire [4:0]  _slots_31_io_uop_br_tag;
  wire [5:0]  _slots_31_io_uop_ftq_idx;
  wire        _slots_31_io_uop_edge_inst;
  wire [5:0]  _slots_31_io_uop_pc_lob;
  wire        _slots_31_io_uop_taken;
  wire [19:0] _slots_31_io_uop_imm_packed;
  wire [6:0]  _slots_31_io_uop_rob_idx;
  wire [4:0]  _slots_31_io_uop_ldq_idx;
  wire [4:0]  _slots_31_io_uop_stq_idx;
  wire [6:0]  _slots_31_io_uop_pdst;
  wire [6:0]  _slots_31_io_uop_prs1;
  wire [6:0]  _slots_31_io_uop_prs2;
  wire        _slots_31_io_uop_bypassable;
  wire [4:0]  _slots_31_io_uop_mem_cmd;
  wire        _slots_31_io_uop_is_amo;
  wire        _slots_31_io_uop_uses_stq;
  wire        _slots_31_io_uop_ldst_val;
  wire [1:0]  _slots_31_io_uop_dst_rtype;
  wire [1:0]  _slots_31_io_uop_lrs1_rtype;
  wire [1:0]  _slots_31_io_uop_lrs2_rtype;
  wire        _slots_31_io_uop_fp_val;
  wire        _slots_30_io_valid;
  wire        _slots_30_io_will_be_valid;
  wire        _slots_30_io_request;
  wire [6:0]  _slots_30_io_out_uop_uopc;
  wire        _slots_30_io_out_uop_is_rvc;
  wire [9:0]  _slots_30_io_out_uop_fu_code;
  wire [1:0]  _slots_30_io_out_uop_iw_state;
  wire        _slots_30_io_out_uop_iw_p1_poisoned;
  wire        _slots_30_io_out_uop_iw_p2_poisoned;
  wire        _slots_30_io_out_uop_is_br;
  wire        _slots_30_io_out_uop_is_jalr;
  wire        _slots_30_io_out_uop_is_jal;
  wire        _slots_30_io_out_uop_is_sfb;
  wire [19:0] _slots_30_io_out_uop_br_mask;
  wire [4:0]  _slots_30_io_out_uop_br_tag;
  wire [5:0]  _slots_30_io_out_uop_ftq_idx;
  wire        _slots_30_io_out_uop_edge_inst;
  wire [5:0]  _slots_30_io_out_uop_pc_lob;
  wire        _slots_30_io_out_uop_taken;
  wire [19:0] _slots_30_io_out_uop_imm_packed;
  wire [6:0]  _slots_30_io_out_uop_rob_idx;
  wire [4:0]  _slots_30_io_out_uop_ldq_idx;
  wire [4:0]  _slots_30_io_out_uop_stq_idx;
  wire [6:0]  _slots_30_io_out_uop_pdst;
  wire [6:0]  _slots_30_io_out_uop_prs1;
  wire [6:0]  _slots_30_io_out_uop_prs2;
  wire [6:0]  _slots_30_io_out_uop_prs3;
  wire        _slots_30_io_out_uop_prs1_busy;
  wire        _slots_30_io_out_uop_prs2_busy;
  wire        _slots_30_io_out_uop_prs3_busy;
  wire        _slots_30_io_out_uop_ppred_busy;
  wire        _slots_30_io_out_uop_bypassable;
  wire [4:0]  _slots_30_io_out_uop_mem_cmd;
  wire [1:0]  _slots_30_io_out_uop_mem_size;
  wire        _slots_30_io_out_uop_mem_signed;
  wire        _slots_30_io_out_uop_is_fence;
  wire        _slots_30_io_out_uop_is_amo;
  wire        _slots_30_io_out_uop_uses_ldq;
  wire        _slots_30_io_out_uop_uses_stq;
  wire        _slots_30_io_out_uop_ldst_val;
  wire [1:0]  _slots_30_io_out_uop_dst_rtype;
  wire [1:0]  _slots_30_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_30_io_out_uop_lrs2_rtype;
  wire        _slots_30_io_out_uop_fp_val;
  wire [6:0]  _slots_30_io_uop_uopc;
  wire        _slots_30_io_uop_is_rvc;
  wire [9:0]  _slots_30_io_uop_fu_code;
  wire        _slots_30_io_uop_iw_p1_poisoned;
  wire        _slots_30_io_uop_iw_p2_poisoned;
  wire        _slots_30_io_uop_is_br;
  wire        _slots_30_io_uop_is_jalr;
  wire        _slots_30_io_uop_is_jal;
  wire        _slots_30_io_uop_is_sfb;
  wire [19:0] _slots_30_io_uop_br_mask;
  wire [4:0]  _slots_30_io_uop_br_tag;
  wire [5:0]  _slots_30_io_uop_ftq_idx;
  wire        _slots_30_io_uop_edge_inst;
  wire [5:0]  _slots_30_io_uop_pc_lob;
  wire        _slots_30_io_uop_taken;
  wire [19:0] _slots_30_io_uop_imm_packed;
  wire [6:0]  _slots_30_io_uop_rob_idx;
  wire [4:0]  _slots_30_io_uop_ldq_idx;
  wire [4:0]  _slots_30_io_uop_stq_idx;
  wire [6:0]  _slots_30_io_uop_pdst;
  wire [6:0]  _slots_30_io_uop_prs1;
  wire [6:0]  _slots_30_io_uop_prs2;
  wire        _slots_30_io_uop_bypassable;
  wire [4:0]  _slots_30_io_uop_mem_cmd;
  wire        _slots_30_io_uop_is_amo;
  wire        _slots_30_io_uop_uses_stq;
  wire        _slots_30_io_uop_ldst_val;
  wire [1:0]  _slots_30_io_uop_dst_rtype;
  wire [1:0]  _slots_30_io_uop_lrs1_rtype;
  wire [1:0]  _slots_30_io_uop_lrs2_rtype;
  wire        _slots_30_io_uop_fp_val;
  wire        _slots_29_io_valid;
  wire        _slots_29_io_will_be_valid;
  wire        _slots_29_io_request;
  wire [6:0]  _slots_29_io_out_uop_uopc;
  wire        _slots_29_io_out_uop_is_rvc;
  wire [9:0]  _slots_29_io_out_uop_fu_code;
  wire [1:0]  _slots_29_io_out_uop_iw_state;
  wire        _slots_29_io_out_uop_iw_p1_poisoned;
  wire        _slots_29_io_out_uop_iw_p2_poisoned;
  wire        _slots_29_io_out_uop_is_br;
  wire        _slots_29_io_out_uop_is_jalr;
  wire        _slots_29_io_out_uop_is_jal;
  wire        _slots_29_io_out_uop_is_sfb;
  wire [19:0] _slots_29_io_out_uop_br_mask;
  wire [4:0]  _slots_29_io_out_uop_br_tag;
  wire [5:0]  _slots_29_io_out_uop_ftq_idx;
  wire        _slots_29_io_out_uop_edge_inst;
  wire [5:0]  _slots_29_io_out_uop_pc_lob;
  wire        _slots_29_io_out_uop_taken;
  wire [19:0] _slots_29_io_out_uop_imm_packed;
  wire [6:0]  _slots_29_io_out_uop_rob_idx;
  wire [4:0]  _slots_29_io_out_uop_ldq_idx;
  wire [4:0]  _slots_29_io_out_uop_stq_idx;
  wire [6:0]  _slots_29_io_out_uop_pdst;
  wire [6:0]  _slots_29_io_out_uop_prs1;
  wire [6:0]  _slots_29_io_out_uop_prs2;
  wire [6:0]  _slots_29_io_out_uop_prs3;
  wire        _slots_29_io_out_uop_prs1_busy;
  wire        _slots_29_io_out_uop_prs2_busy;
  wire        _slots_29_io_out_uop_prs3_busy;
  wire        _slots_29_io_out_uop_ppred_busy;
  wire        _slots_29_io_out_uop_bypassable;
  wire [4:0]  _slots_29_io_out_uop_mem_cmd;
  wire [1:0]  _slots_29_io_out_uop_mem_size;
  wire        _slots_29_io_out_uop_mem_signed;
  wire        _slots_29_io_out_uop_is_fence;
  wire        _slots_29_io_out_uop_is_amo;
  wire        _slots_29_io_out_uop_uses_ldq;
  wire        _slots_29_io_out_uop_uses_stq;
  wire        _slots_29_io_out_uop_ldst_val;
  wire [1:0]  _slots_29_io_out_uop_dst_rtype;
  wire [1:0]  _slots_29_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_29_io_out_uop_lrs2_rtype;
  wire        _slots_29_io_out_uop_fp_val;
  wire [6:0]  _slots_29_io_uop_uopc;
  wire        _slots_29_io_uop_is_rvc;
  wire [9:0]  _slots_29_io_uop_fu_code;
  wire        _slots_29_io_uop_iw_p1_poisoned;
  wire        _slots_29_io_uop_iw_p2_poisoned;
  wire        _slots_29_io_uop_is_br;
  wire        _slots_29_io_uop_is_jalr;
  wire        _slots_29_io_uop_is_jal;
  wire        _slots_29_io_uop_is_sfb;
  wire [19:0] _slots_29_io_uop_br_mask;
  wire [4:0]  _slots_29_io_uop_br_tag;
  wire [5:0]  _slots_29_io_uop_ftq_idx;
  wire        _slots_29_io_uop_edge_inst;
  wire [5:0]  _slots_29_io_uop_pc_lob;
  wire        _slots_29_io_uop_taken;
  wire [19:0] _slots_29_io_uop_imm_packed;
  wire [6:0]  _slots_29_io_uop_rob_idx;
  wire [4:0]  _slots_29_io_uop_ldq_idx;
  wire [4:0]  _slots_29_io_uop_stq_idx;
  wire [6:0]  _slots_29_io_uop_pdst;
  wire [6:0]  _slots_29_io_uop_prs1;
  wire [6:0]  _slots_29_io_uop_prs2;
  wire        _slots_29_io_uop_bypassable;
  wire [4:0]  _slots_29_io_uop_mem_cmd;
  wire        _slots_29_io_uop_is_amo;
  wire        _slots_29_io_uop_uses_stq;
  wire        _slots_29_io_uop_ldst_val;
  wire [1:0]  _slots_29_io_uop_dst_rtype;
  wire [1:0]  _slots_29_io_uop_lrs1_rtype;
  wire [1:0]  _slots_29_io_uop_lrs2_rtype;
  wire        _slots_29_io_uop_fp_val;
  wire        _slots_28_io_valid;
  wire        _slots_28_io_will_be_valid;
  wire        _slots_28_io_request;
  wire [6:0]  _slots_28_io_out_uop_uopc;
  wire        _slots_28_io_out_uop_is_rvc;
  wire [9:0]  _slots_28_io_out_uop_fu_code;
  wire [1:0]  _slots_28_io_out_uop_iw_state;
  wire        _slots_28_io_out_uop_iw_p1_poisoned;
  wire        _slots_28_io_out_uop_iw_p2_poisoned;
  wire        _slots_28_io_out_uop_is_br;
  wire        _slots_28_io_out_uop_is_jalr;
  wire        _slots_28_io_out_uop_is_jal;
  wire        _slots_28_io_out_uop_is_sfb;
  wire [19:0] _slots_28_io_out_uop_br_mask;
  wire [4:0]  _slots_28_io_out_uop_br_tag;
  wire [5:0]  _slots_28_io_out_uop_ftq_idx;
  wire        _slots_28_io_out_uop_edge_inst;
  wire [5:0]  _slots_28_io_out_uop_pc_lob;
  wire        _slots_28_io_out_uop_taken;
  wire [19:0] _slots_28_io_out_uop_imm_packed;
  wire [6:0]  _slots_28_io_out_uop_rob_idx;
  wire [4:0]  _slots_28_io_out_uop_ldq_idx;
  wire [4:0]  _slots_28_io_out_uop_stq_idx;
  wire [6:0]  _slots_28_io_out_uop_pdst;
  wire [6:0]  _slots_28_io_out_uop_prs1;
  wire [6:0]  _slots_28_io_out_uop_prs2;
  wire [6:0]  _slots_28_io_out_uop_prs3;
  wire        _slots_28_io_out_uop_prs1_busy;
  wire        _slots_28_io_out_uop_prs2_busy;
  wire        _slots_28_io_out_uop_prs3_busy;
  wire        _slots_28_io_out_uop_ppred_busy;
  wire        _slots_28_io_out_uop_bypassable;
  wire [4:0]  _slots_28_io_out_uop_mem_cmd;
  wire [1:0]  _slots_28_io_out_uop_mem_size;
  wire        _slots_28_io_out_uop_mem_signed;
  wire        _slots_28_io_out_uop_is_fence;
  wire        _slots_28_io_out_uop_is_amo;
  wire        _slots_28_io_out_uop_uses_ldq;
  wire        _slots_28_io_out_uop_uses_stq;
  wire        _slots_28_io_out_uop_ldst_val;
  wire [1:0]  _slots_28_io_out_uop_dst_rtype;
  wire [1:0]  _slots_28_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_28_io_out_uop_lrs2_rtype;
  wire        _slots_28_io_out_uop_fp_val;
  wire [6:0]  _slots_28_io_uop_uopc;
  wire        _slots_28_io_uop_is_rvc;
  wire [9:0]  _slots_28_io_uop_fu_code;
  wire        _slots_28_io_uop_iw_p1_poisoned;
  wire        _slots_28_io_uop_iw_p2_poisoned;
  wire        _slots_28_io_uop_is_br;
  wire        _slots_28_io_uop_is_jalr;
  wire        _slots_28_io_uop_is_jal;
  wire        _slots_28_io_uop_is_sfb;
  wire [19:0] _slots_28_io_uop_br_mask;
  wire [4:0]  _slots_28_io_uop_br_tag;
  wire [5:0]  _slots_28_io_uop_ftq_idx;
  wire        _slots_28_io_uop_edge_inst;
  wire [5:0]  _slots_28_io_uop_pc_lob;
  wire        _slots_28_io_uop_taken;
  wire [19:0] _slots_28_io_uop_imm_packed;
  wire [6:0]  _slots_28_io_uop_rob_idx;
  wire [4:0]  _slots_28_io_uop_ldq_idx;
  wire [4:0]  _slots_28_io_uop_stq_idx;
  wire [6:0]  _slots_28_io_uop_pdst;
  wire [6:0]  _slots_28_io_uop_prs1;
  wire [6:0]  _slots_28_io_uop_prs2;
  wire        _slots_28_io_uop_bypassable;
  wire [4:0]  _slots_28_io_uop_mem_cmd;
  wire        _slots_28_io_uop_is_amo;
  wire        _slots_28_io_uop_uses_stq;
  wire        _slots_28_io_uop_ldst_val;
  wire [1:0]  _slots_28_io_uop_dst_rtype;
  wire [1:0]  _slots_28_io_uop_lrs1_rtype;
  wire [1:0]  _slots_28_io_uop_lrs2_rtype;
  wire        _slots_28_io_uop_fp_val;
  wire        _slots_27_io_valid;
  wire        _slots_27_io_will_be_valid;
  wire        _slots_27_io_request;
  wire [6:0]  _slots_27_io_out_uop_uopc;
  wire        _slots_27_io_out_uop_is_rvc;
  wire [9:0]  _slots_27_io_out_uop_fu_code;
  wire [1:0]  _slots_27_io_out_uop_iw_state;
  wire        _slots_27_io_out_uop_iw_p1_poisoned;
  wire        _slots_27_io_out_uop_iw_p2_poisoned;
  wire        _slots_27_io_out_uop_is_br;
  wire        _slots_27_io_out_uop_is_jalr;
  wire        _slots_27_io_out_uop_is_jal;
  wire        _slots_27_io_out_uop_is_sfb;
  wire [19:0] _slots_27_io_out_uop_br_mask;
  wire [4:0]  _slots_27_io_out_uop_br_tag;
  wire [5:0]  _slots_27_io_out_uop_ftq_idx;
  wire        _slots_27_io_out_uop_edge_inst;
  wire [5:0]  _slots_27_io_out_uop_pc_lob;
  wire        _slots_27_io_out_uop_taken;
  wire [19:0] _slots_27_io_out_uop_imm_packed;
  wire [6:0]  _slots_27_io_out_uop_rob_idx;
  wire [4:0]  _slots_27_io_out_uop_ldq_idx;
  wire [4:0]  _slots_27_io_out_uop_stq_idx;
  wire [6:0]  _slots_27_io_out_uop_pdst;
  wire [6:0]  _slots_27_io_out_uop_prs1;
  wire [6:0]  _slots_27_io_out_uop_prs2;
  wire [6:0]  _slots_27_io_out_uop_prs3;
  wire        _slots_27_io_out_uop_prs1_busy;
  wire        _slots_27_io_out_uop_prs2_busy;
  wire        _slots_27_io_out_uop_prs3_busy;
  wire        _slots_27_io_out_uop_ppred_busy;
  wire        _slots_27_io_out_uop_bypassable;
  wire [4:0]  _slots_27_io_out_uop_mem_cmd;
  wire [1:0]  _slots_27_io_out_uop_mem_size;
  wire        _slots_27_io_out_uop_mem_signed;
  wire        _slots_27_io_out_uop_is_fence;
  wire        _slots_27_io_out_uop_is_amo;
  wire        _slots_27_io_out_uop_uses_ldq;
  wire        _slots_27_io_out_uop_uses_stq;
  wire        _slots_27_io_out_uop_ldst_val;
  wire [1:0]  _slots_27_io_out_uop_dst_rtype;
  wire [1:0]  _slots_27_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_27_io_out_uop_lrs2_rtype;
  wire        _slots_27_io_out_uop_fp_val;
  wire [6:0]  _slots_27_io_uop_uopc;
  wire        _slots_27_io_uop_is_rvc;
  wire [9:0]  _slots_27_io_uop_fu_code;
  wire        _slots_27_io_uop_iw_p1_poisoned;
  wire        _slots_27_io_uop_iw_p2_poisoned;
  wire        _slots_27_io_uop_is_br;
  wire        _slots_27_io_uop_is_jalr;
  wire        _slots_27_io_uop_is_jal;
  wire        _slots_27_io_uop_is_sfb;
  wire [19:0] _slots_27_io_uop_br_mask;
  wire [4:0]  _slots_27_io_uop_br_tag;
  wire [5:0]  _slots_27_io_uop_ftq_idx;
  wire        _slots_27_io_uop_edge_inst;
  wire [5:0]  _slots_27_io_uop_pc_lob;
  wire        _slots_27_io_uop_taken;
  wire [19:0] _slots_27_io_uop_imm_packed;
  wire [6:0]  _slots_27_io_uop_rob_idx;
  wire [4:0]  _slots_27_io_uop_ldq_idx;
  wire [4:0]  _slots_27_io_uop_stq_idx;
  wire [6:0]  _slots_27_io_uop_pdst;
  wire [6:0]  _slots_27_io_uop_prs1;
  wire [6:0]  _slots_27_io_uop_prs2;
  wire        _slots_27_io_uop_bypassable;
  wire [4:0]  _slots_27_io_uop_mem_cmd;
  wire        _slots_27_io_uop_is_amo;
  wire        _slots_27_io_uop_uses_stq;
  wire        _slots_27_io_uop_ldst_val;
  wire [1:0]  _slots_27_io_uop_dst_rtype;
  wire [1:0]  _slots_27_io_uop_lrs1_rtype;
  wire [1:0]  _slots_27_io_uop_lrs2_rtype;
  wire        _slots_27_io_uop_fp_val;
  wire        _slots_26_io_valid;
  wire        _slots_26_io_will_be_valid;
  wire        _slots_26_io_request;
  wire [6:0]  _slots_26_io_out_uop_uopc;
  wire        _slots_26_io_out_uop_is_rvc;
  wire [9:0]  _slots_26_io_out_uop_fu_code;
  wire [1:0]  _slots_26_io_out_uop_iw_state;
  wire        _slots_26_io_out_uop_iw_p1_poisoned;
  wire        _slots_26_io_out_uop_iw_p2_poisoned;
  wire        _slots_26_io_out_uop_is_br;
  wire        _slots_26_io_out_uop_is_jalr;
  wire        _slots_26_io_out_uop_is_jal;
  wire        _slots_26_io_out_uop_is_sfb;
  wire [19:0] _slots_26_io_out_uop_br_mask;
  wire [4:0]  _slots_26_io_out_uop_br_tag;
  wire [5:0]  _slots_26_io_out_uop_ftq_idx;
  wire        _slots_26_io_out_uop_edge_inst;
  wire [5:0]  _slots_26_io_out_uop_pc_lob;
  wire        _slots_26_io_out_uop_taken;
  wire [19:0] _slots_26_io_out_uop_imm_packed;
  wire [6:0]  _slots_26_io_out_uop_rob_idx;
  wire [4:0]  _slots_26_io_out_uop_ldq_idx;
  wire [4:0]  _slots_26_io_out_uop_stq_idx;
  wire [6:0]  _slots_26_io_out_uop_pdst;
  wire [6:0]  _slots_26_io_out_uop_prs1;
  wire [6:0]  _slots_26_io_out_uop_prs2;
  wire [6:0]  _slots_26_io_out_uop_prs3;
  wire        _slots_26_io_out_uop_prs1_busy;
  wire        _slots_26_io_out_uop_prs2_busy;
  wire        _slots_26_io_out_uop_prs3_busy;
  wire        _slots_26_io_out_uop_ppred_busy;
  wire        _slots_26_io_out_uop_bypassable;
  wire [4:0]  _slots_26_io_out_uop_mem_cmd;
  wire [1:0]  _slots_26_io_out_uop_mem_size;
  wire        _slots_26_io_out_uop_mem_signed;
  wire        _slots_26_io_out_uop_is_fence;
  wire        _slots_26_io_out_uop_is_amo;
  wire        _slots_26_io_out_uop_uses_ldq;
  wire        _slots_26_io_out_uop_uses_stq;
  wire        _slots_26_io_out_uop_ldst_val;
  wire [1:0]  _slots_26_io_out_uop_dst_rtype;
  wire [1:0]  _slots_26_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_26_io_out_uop_lrs2_rtype;
  wire        _slots_26_io_out_uop_fp_val;
  wire [6:0]  _slots_26_io_uop_uopc;
  wire        _slots_26_io_uop_is_rvc;
  wire [9:0]  _slots_26_io_uop_fu_code;
  wire        _slots_26_io_uop_iw_p1_poisoned;
  wire        _slots_26_io_uop_iw_p2_poisoned;
  wire        _slots_26_io_uop_is_br;
  wire        _slots_26_io_uop_is_jalr;
  wire        _slots_26_io_uop_is_jal;
  wire        _slots_26_io_uop_is_sfb;
  wire [19:0] _slots_26_io_uop_br_mask;
  wire [4:0]  _slots_26_io_uop_br_tag;
  wire [5:0]  _slots_26_io_uop_ftq_idx;
  wire        _slots_26_io_uop_edge_inst;
  wire [5:0]  _slots_26_io_uop_pc_lob;
  wire        _slots_26_io_uop_taken;
  wire [19:0] _slots_26_io_uop_imm_packed;
  wire [6:0]  _slots_26_io_uop_rob_idx;
  wire [4:0]  _slots_26_io_uop_ldq_idx;
  wire [4:0]  _slots_26_io_uop_stq_idx;
  wire [6:0]  _slots_26_io_uop_pdst;
  wire [6:0]  _slots_26_io_uop_prs1;
  wire [6:0]  _slots_26_io_uop_prs2;
  wire        _slots_26_io_uop_bypassable;
  wire [4:0]  _slots_26_io_uop_mem_cmd;
  wire        _slots_26_io_uop_is_amo;
  wire        _slots_26_io_uop_uses_stq;
  wire        _slots_26_io_uop_ldst_val;
  wire [1:0]  _slots_26_io_uop_dst_rtype;
  wire [1:0]  _slots_26_io_uop_lrs1_rtype;
  wire [1:0]  _slots_26_io_uop_lrs2_rtype;
  wire        _slots_26_io_uop_fp_val;
  wire        _slots_25_io_valid;
  wire        _slots_25_io_will_be_valid;
  wire        _slots_25_io_request;
  wire [6:0]  _slots_25_io_out_uop_uopc;
  wire        _slots_25_io_out_uop_is_rvc;
  wire [9:0]  _slots_25_io_out_uop_fu_code;
  wire [1:0]  _slots_25_io_out_uop_iw_state;
  wire        _slots_25_io_out_uop_iw_p1_poisoned;
  wire        _slots_25_io_out_uop_iw_p2_poisoned;
  wire        _slots_25_io_out_uop_is_br;
  wire        _slots_25_io_out_uop_is_jalr;
  wire        _slots_25_io_out_uop_is_jal;
  wire        _slots_25_io_out_uop_is_sfb;
  wire [19:0] _slots_25_io_out_uop_br_mask;
  wire [4:0]  _slots_25_io_out_uop_br_tag;
  wire [5:0]  _slots_25_io_out_uop_ftq_idx;
  wire        _slots_25_io_out_uop_edge_inst;
  wire [5:0]  _slots_25_io_out_uop_pc_lob;
  wire        _slots_25_io_out_uop_taken;
  wire [19:0] _slots_25_io_out_uop_imm_packed;
  wire [6:0]  _slots_25_io_out_uop_rob_idx;
  wire [4:0]  _slots_25_io_out_uop_ldq_idx;
  wire [4:0]  _slots_25_io_out_uop_stq_idx;
  wire [6:0]  _slots_25_io_out_uop_pdst;
  wire [6:0]  _slots_25_io_out_uop_prs1;
  wire [6:0]  _slots_25_io_out_uop_prs2;
  wire [6:0]  _slots_25_io_out_uop_prs3;
  wire        _slots_25_io_out_uop_prs1_busy;
  wire        _slots_25_io_out_uop_prs2_busy;
  wire        _slots_25_io_out_uop_prs3_busy;
  wire        _slots_25_io_out_uop_ppred_busy;
  wire        _slots_25_io_out_uop_bypassable;
  wire [4:0]  _slots_25_io_out_uop_mem_cmd;
  wire [1:0]  _slots_25_io_out_uop_mem_size;
  wire        _slots_25_io_out_uop_mem_signed;
  wire        _slots_25_io_out_uop_is_fence;
  wire        _slots_25_io_out_uop_is_amo;
  wire        _slots_25_io_out_uop_uses_ldq;
  wire        _slots_25_io_out_uop_uses_stq;
  wire        _slots_25_io_out_uop_ldst_val;
  wire [1:0]  _slots_25_io_out_uop_dst_rtype;
  wire [1:0]  _slots_25_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_25_io_out_uop_lrs2_rtype;
  wire        _slots_25_io_out_uop_fp_val;
  wire [6:0]  _slots_25_io_uop_uopc;
  wire        _slots_25_io_uop_is_rvc;
  wire [9:0]  _slots_25_io_uop_fu_code;
  wire        _slots_25_io_uop_iw_p1_poisoned;
  wire        _slots_25_io_uop_iw_p2_poisoned;
  wire        _slots_25_io_uop_is_br;
  wire        _slots_25_io_uop_is_jalr;
  wire        _slots_25_io_uop_is_jal;
  wire        _slots_25_io_uop_is_sfb;
  wire [19:0] _slots_25_io_uop_br_mask;
  wire [4:0]  _slots_25_io_uop_br_tag;
  wire [5:0]  _slots_25_io_uop_ftq_idx;
  wire        _slots_25_io_uop_edge_inst;
  wire [5:0]  _slots_25_io_uop_pc_lob;
  wire        _slots_25_io_uop_taken;
  wire [19:0] _slots_25_io_uop_imm_packed;
  wire [6:0]  _slots_25_io_uop_rob_idx;
  wire [4:0]  _slots_25_io_uop_ldq_idx;
  wire [4:0]  _slots_25_io_uop_stq_idx;
  wire [6:0]  _slots_25_io_uop_pdst;
  wire [6:0]  _slots_25_io_uop_prs1;
  wire [6:0]  _slots_25_io_uop_prs2;
  wire        _slots_25_io_uop_bypassable;
  wire [4:0]  _slots_25_io_uop_mem_cmd;
  wire        _slots_25_io_uop_is_amo;
  wire        _slots_25_io_uop_uses_stq;
  wire        _slots_25_io_uop_ldst_val;
  wire [1:0]  _slots_25_io_uop_dst_rtype;
  wire [1:0]  _slots_25_io_uop_lrs1_rtype;
  wire [1:0]  _slots_25_io_uop_lrs2_rtype;
  wire        _slots_25_io_uop_fp_val;
  wire        _slots_24_io_valid;
  wire        _slots_24_io_will_be_valid;
  wire        _slots_24_io_request;
  wire [6:0]  _slots_24_io_out_uop_uopc;
  wire        _slots_24_io_out_uop_is_rvc;
  wire [9:0]  _slots_24_io_out_uop_fu_code;
  wire [1:0]  _slots_24_io_out_uop_iw_state;
  wire        _slots_24_io_out_uop_iw_p1_poisoned;
  wire        _slots_24_io_out_uop_iw_p2_poisoned;
  wire        _slots_24_io_out_uop_is_br;
  wire        _slots_24_io_out_uop_is_jalr;
  wire        _slots_24_io_out_uop_is_jal;
  wire        _slots_24_io_out_uop_is_sfb;
  wire [19:0] _slots_24_io_out_uop_br_mask;
  wire [4:0]  _slots_24_io_out_uop_br_tag;
  wire [5:0]  _slots_24_io_out_uop_ftq_idx;
  wire        _slots_24_io_out_uop_edge_inst;
  wire [5:0]  _slots_24_io_out_uop_pc_lob;
  wire        _slots_24_io_out_uop_taken;
  wire [19:0] _slots_24_io_out_uop_imm_packed;
  wire [6:0]  _slots_24_io_out_uop_rob_idx;
  wire [4:0]  _slots_24_io_out_uop_ldq_idx;
  wire [4:0]  _slots_24_io_out_uop_stq_idx;
  wire [6:0]  _slots_24_io_out_uop_pdst;
  wire [6:0]  _slots_24_io_out_uop_prs1;
  wire [6:0]  _slots_24_io_out_uop_prs2;
  wire [6:0]  _slots_24_io_out_uop_prs3;
  wire        _slots_24_io_out_uop_prs1_busy;
  wire        _slots_24_io_out_uop_prs2_busy;
  wire        _slots_24_io_out_uop_prs3_busy;
  wire        _slots_24_io_out_uop_ppred_busy;
  wire        _slots_24_io_out_uop_bypassable;
  wire [4:0]  _slots_24_io_out_uop_mem_cmd;
  wire [1:0]  _slots_24_io_out_uop_mem_size;
  wire        _slots_24_io_out_uop_mem_signed;
  wire        _slots_24_io_out_uop_is_fence;
  wire        _slots_24_io_out_uop_is_amo;
  wire        _slots_24_io_out_uop_uses_ldq;
  wire        _slots_24_io_out_uop_uses_stq;
  wire        _slots_24_io_out_uop_ldst_val;
  wire [1:0]  _slots_24_io_out_uop_dst_rtype;
  wire [1:0]  _slots_24_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_24_io_out_uop_lrs2_rtype;
  wire        _slots_24_io_out_uop_fp_val;
  wire [6:0]  _slots_24_io_uop_uopc;
  wire        _slots_24_io_uop_is_rvc;
  wire [9:0]  _slots_24_io_uop_fu_code;
  wire        _slots_24_io_uop_iw_p1_poisoned;
  wire        _slots_24_io_uop_iw_p2_poisoned;
  wire        _slots_24_io_uop_is_br;
  wire        _slots_24_io_uop_is_jalr;
  wire        _slots_24_io_uop_is_jal;
  wire        _slots_24_io_uop_is_sfb;
  wire [19:0] _slots_24_io_uop_br_mask;
  wire [4:0]  _slots_24_io_uop_br_tag;
  wire [5:0]  _slots_24_io_uop_ftq_idx;
  wire        _slots_24_io_uop_edge_inst;
  wire [5:0]  _slots_24_io_uop_pc_lob;
  wire        _slots_24_io_uop_taken;
  wire [19:0] _slots_24_io_uop_imm_packed;
  wire [6:0]  _slots_24_io_uop_rob_idx;
  wire [4:0]  _slots_24_io_uop_ldq_idx;
  wire [4:0]  _slots_24_io_uop_stq_idx;
  wire [6:0]  _slots_24_io_uop_pdst;
  wire [6:0]  _slots_24_io_uop_prs1;
  wire [6:0]  _slots_24_io_uop_prs2;
  wire        _slots_24_io_uop_bypassable;
  wire [4:0]  _slots_24_io_uop_mem_cmd;
  wire        _slots_24_io_uop_is_amo;
  wire        _slots_24_io_uop_uses_stq;
  wire        _slots_24_io_uop_ldst_val;
  wire [1:0]  _slots_24_io_uop_dst_rtype;
  wire [1:0]  _slots_24_io_uop_lrs1_rtype;
  wire [1:0]  _slots_24_io_uop_lrs2_rtype;
  wire        _slots_24_io_uop_fp_val;
  wire        _slots_23_io_valid;
  wire        _slots_23_io_will_be_valid;
  wire        _slots_23_io_request;
  wire [6:0]  _slots_23_io_out_uop_uopc;
  wire        _slots_23_io_out_uop_is_rvc;
  wire [9:0]  _slots_23_io_out_uop_fu_code;
  wire [1:0]  _slots_23_io_out_uop_iw_state;
  wire        _slots_23_io_out_uop_iw_p1_poisoned;
  wire        _slots_23_io_out_uop_iw_p2_poisoned;
  wire        _slots_23_io_out_uop_is_br;
  wire        _slots_23_io_out_uop_is_jalr;
  wire        _slots_23_io_out_uop_is_jal;
  wire        _slots_23_io_out_uop_is_sfb;
  wire [19:0] _slots_23_io_out_uop_br_mask;
  wire [4:0]  _slots_23_io_out_uop_br_tag;
  wire [5:0]  _slots_23_io_out_uop_ftq_idx;
  wire        _slots_23_io_out_uop_edge_inst;
  wire [5:0]  _slots_23_io_out_uop_pc_lob;
  wire        _slots_23_io_out_uop_taken;
  wire [19:0] _slots_23_io_out_uop_imm_packed;
  wire [6:0]  _slots_23_io_out_uop_rob_idx;
  wire [4:0]  _slots_23_io_out_uop_ldq_idx;
  wire [4:0]  _slots_23_io_out_uop_stq_idx;
  wire [6:0]  _slots_23_io_out_uop_pdst;
  wire [6:0]  _slots_23_io_out_uop_prs1;
  wire [6:0]  _slots_23_io_out_uop_prs2;
  wire [6:0]  _slots_23_io_out_uop_prs3;
  wire        _slots_23_io_out_uop_prs1_busy;
  wire        _slots_23_io_out_uop_prs2_busy;
  wire        _slots_23_io_out_uop_prs3_busy;
  wire        _slots_23_io_out_uop_ppred_busy;
  wire        _slots_23_io_out_uop_bypassable;
  wire [4:0]  _slots_23_io_out_uop_mem_cmd;
  wire [1:0]  _slots_23_io_out_uop_mem_size;
  wire        _slots_23_io_out_uop_mem_signed;
  wire        _slots_23_io_out_uop_is_fence;
  wire        _slots_23_io_out_uop_is_amo;
  wire        _slots_23_io_out_uop_uses_ldq;
  wire        _slots_23_io_out_uop_uses_stq;
  wire        _slots_23_io_out_uop_ldst_val;
  wire [1:0]  _slots_23_io_out_uop_dst_rtype;
  wire [1:0]  _slots_23_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_23_io_out_uop_lrs2_rtype;
  wire        _slots_23_io_out_uop_fp_val;
  wire [6:0]  _slots_23_io_uop_uopc;
  wire        _slots_23_io_uop_is_rvc;
  wire [9:0]  _slots_23_io_uop_fu_code;
  wire        _slots_23_io_uop_iw_p1_poisoned;
  wire        _slots_23_io_uop_iw_p2_poisoned;
  wire        _slots_23_io_uop_is_br;
  wire        _slots_23_io_uop_is_jalr;
  wire        _slots_23_io_uop_is_jal;
  wire        _slots_23_io_uop_is_sfb;
  wire [19:0] _slots_23_io_uop_br_mask;
  wire [4:0]  _slots_23_io_uop_br_tag;
  wire [5:0]  _slots_23_io_uop_ftq_idx;
  wire        _slots_23_io_uop_edge_inst;
  wire [5:0]  _slots_23_io_uop_pc_lob;
  wire        _slots_23_io_uop_taken;
  wire [19:0] _slots_23_io_uop_imm_packed;
  wire [6:0]  _slots_23_io_uop_rob_idx;
  wire [4:0]  _slots_23_io_uop_ldq_idx;
  wire [4:0]  _slots_23_io_uop_stq_idx;
  wire [6:0]  _slots_23_io_uop_pdst;
  wire [6:0]  _slots_23_io_uop_prs1;
  wire [6:0]  _slots_23_io_uop_prs2;
  wire        _slots_23_io_uop_bypassable;
  wire [4:0]  _slots_23_io_uop_mem_cmd;
  wire        _slots_23_io_uop_is_amo;
  wire        _slots_23_io_uop_uses_stq;
  wire        _slots_23_io_uop_ldst_val;
  wire [1:0]  _slots_23_io_uop_dst_rtype;
  wire [1:0]  _slots_23_io_uop_lrs1_rtype;
  wire [1:0]  _slots_23_io_uop_lrs2_rtype;
  wire        _slots_23_io_uop_fp_val;
  wire        _slots_22_io_valid;
  wire        _slots_22_io_will_be_valid;
  wire        _slots_22_io_request;
  wire [6:0]  _slots_22_io_out_uop_uopc;
  wire        _slots_22_io_out_uop_is_rvc;
  wire [9:0]  _slots_22_io_out_uop_fu_code;
  wire [1:0]  _slots_22_io_out_uop_iw_state;
  wire        _slots_22_io_out_uop_iw_p1_poisoned;
  wire        _slots_22_io_out_uop_iw_p2_poisoned;
  wire        _slots_22_io_out_uop_is_br;
  wire        _slots_22_io_out_uop_is_jalr;
  wire        _slots_22_io_out_uop_is_jal;
  wire        _slots_22_io_out_uop_is_sfb;
  wire [19:0] _slots_22_io_out_uop_br_mask;
  wire [4:0]  _slots_22_io_out_uop_br_tag;
  wire [5:0]  _slots_22_io_out_uop_ftq_idx;
  wire        _slots_22_io_out_uop_edge_inst;
  wire [5:0]  _slots_22_io_out_uop_pc_lob;
  wire        _slots_22_io_out_uop_taken;
  wire [19:0] _slots_22_io_out_uop_imm_packed;
  wire [6:0]  _slots_22_io_out_uop_rob_idx;
  wire [4:0]  _slots_22_io_out_uop_ldq_idx;
  wire [4:0]  _slots_22_io_out_uop_stq_idx;
  wire [6:0]  _slots_22_io_out_uop_pdst;
  wire [6:0]  _slots_22_io_out_uop_prs1;
  wire [6:0]  _slots_22_io_out_uop_prs2;
  wire [6:0]  _slots_22_io_out_uop_prs3;
  wire        _slots_22_io_out_uop_prs1_busy;
  wire        _slots_22_io_out_uop_prs2_busy;
  wire        _slots_22_io_out_uop_prs3_busy;
  wire        _slots_22_io_out_uop_ppred_busy;
  wire        _slots_22_io_out_uop_bypassable;
  wire [4:0]  _slots_22_io_out_uop_mem_cmd;
  wire [1:0]  _slots_22_io_out_uop_mem_size;
  wire        _slots_22_io_out_uop_mem_signed;
  wire        _slots_22_io_out_uop_is_fence;
  wire        _slots_22_io_out_uop_is_amo;
  wire        _slots_22_io_out_uop_uses_ldq;
  wire        _slots_22_io_out_uop_uses_stq;
  wire        _slots_22_io_out_uop_ldst_val;
  wire [1:0]  _slots_22_io_out_uop_dst_rtype;
  wire [1:0]  _slots_22_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_22_io_out_uop_lrs2_rtype;
  wire        _slots_22_io_out_uop_fp_val;
  wire [6:0]  _slots_22_io_uop_uopc;
  wire        _slots_22_io_uop_is_rvc;
  wire [9:0]  _slots_22_io_uop_fu_code;
  wire        _slots_22_io_uop_iw_p1_poisoned;
  wire        _slots_22_io_uop_iw_p2_poisoned;
  wire        _slots_22_io_uop_is_br;
  wire        _slots_22_io_uop_is_jalr;
  wire        _slots_22_io_uop_is_jal;
  wire        _slots_22_io_uop_is_sfb;
  wire [19:0] _slots_22_io_uop_br_mask;
  wire [4:0]  _slots_22_io_uop_br_tag;
  wire [5:0]  _slots_22_io_uop_ftq_idx;
  wire        _slots_22_io_uop_edge_inst;
  wire [5:0]  _slots_22_io_uop_pc_lob;
  wire        _slots_22_io_uop_taken;
  wire [19:0] _slots_22_io_uop_imm_packed;
  wire [6:0]  _slots_22_io_uop_rob_idx;
  wire [4:0]  _slots_22_io_uop_ldq_idx;
  wire [4:0]  _slots_22_io_uop_stq_idx;
  wire [6:0]  _slots_22_io_uop_pdst;
  wire [6:0]  _slots_22_io_uop_prs1;
  wire [6:0]  _slots_22_io_uop_prs2;
  wire        _slots_22_io_uop_bypassable;
  wire [4:0]  _slots_22_io_uop_mem_cmd;
  wire        _slots_22_io_uop_is_amo;
  wire        _slots_22_io_uop_uses_stq;
  wire        _slots_22_io_uop_ldst_val;
  wire [1:0]  _slots_22_io_uop_dst_rtype;
  wire [1:0]  _slots_22_io_uop_lrs1_rtype;
  wire [1:0]  _slots_22_io_uop_lrs2_rtype;
  wire        _slots_22_io_uop_fp_val;
  wire        _slots_21_io_valid;
  wire        _slots_21_io_will_be_valid;
  wire        _slots_21_io_request;
  wire [6:0]  _slots_21_io_out_uop_uopc;
  wire        _slots_21_io_out_uop_is_rvc;
  wire [9:0]  _slots_21_io_out_uop_fu_code;
  wire [1:0]  _slots_21_io_out_uop_iw_state;
  wire        _slots_21_io_out_uop_iw_p1_poisoned;
  wire        _slots_21_io_out_uop_iw_p2_poisoned;
  wire        _slots_21_io_out_uop_is_br;
  wire        _slots_21_io_out_uop_is_jalr;
  wire        _slots_21_io_out_uop_is_jal;
  wire        _slots_21_io_out_uop_is_sfb;
  wire [19:0] _slots_21_io_out_uop_br_mask;
  wire [4:0]  _slots_21_io_out_uop_br_tag;
  wire [5:0]  _slots_21_io_out_uop_ftq_idx;
  wire        _slots_21_io_out_uop_edge_inst;
  wire [5:0]  _slots_21_io_out_uop_pc_lob;
  wire        _slots_21_io_out_uop_taken;
  wire [19:0] _slots_21_io_out_uop_imm_packed;
  wire [6:0]  _slots_21_io_out_uop_rob_idx;
  wire [4:0]  _slots_21_io_out_uop_ldq_idx;
  wire [4:0]  _slots_21_io_out_uop_stq_idx;
  wire [6:0]  _slots_21_io_out_uop_pdst;
  wire [6:0]  _slots_21_io_out_uop_prs1;
  wire [6:0]  _slots_21_io_out_uop_prs2;
  wire [6:0]  _slots_21_io_out_uop_prs3;
  wire        _slots_21_io_out_uop_prs1_busy;
  wire        _slots_21_io_out_uop_prs2_busy;
  wire        _slots_21_io_out_uop_prs3_busy;
  wire        _slots_21_io_out_uop_ppred_busy;
  wire        _slots_21_io_out_uop_bypassable;
  wire [4:0]  _slots_21_io_out_uop_mem_cmd;
  wire [1:0]  _slots_21_io_out_uop_mem_size;
  wire        _slots_21_io_out_uop_mem_signed;
  wire        _slots_21_io_out_uop_is_fence;
  wire        _slots_21_io_out_uop_is_amo;
  wire        _slots_21_io_out_uop_uses_ldq;
  wire        _slots_21_io_out_uop_uses_stq;
  wire        _slots_21_io_out_uop_ldst_val;
  wire [1:0]  _slots_21_io_out_uop_dst_rtype;
  wire [1:0]  _slots_21_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_21_io_out_uop_lrs2_rtype;
  wire        _slots_21_io_out_uop_fp_val;
  wire [6:0]  _slots_21_io_uop_uopc;
  wire        _slots_21_io_uop_is_rvc;
  wire [9:0]  _slots_21_io_uop_fu_code;
  wire        _slots_21_io_uop_iw_p1_poisoned;
  wire        _slots_21_io_uop_iw_p2_poisoned;
  wire        _slots_21_io_uop_is_br;
  wire        _slots_21_io_uop_is_jalr;
  wire        _slots_21_io_uop_is_jal;
  wire        _slots_21_io_uop_is_sfb;
  wire [19:0] _slots_21_io_uop_br_mask;
  wire [4:0]  _slots_21_io_uop_br_tag;
  wire [5:0]  _slots_21_io_uop_ftq_idx;
  wire        _slots_21_io_uop_edge_inst;
  wire [5:0]  _slots_21_io_uop_pc_lob;
  wire        _slots_21_io_uop_taken;
  wire [19:0] _slots_21_io_uop_imm_packed;
  wire [6:0]  _slots_21_io_uop_rob_idx;
  wire [4:0]  _slots_21_io_uop_ldq_idx;
  wire [4:0]  _slots_21_io_uop_stq_idx;
  wire [6:0]  _slots_21_io_uop_pdst;
  wire [6:0]  _slots_21_io_uop_prs1;
  wire [6:0]  _slots_21_io_uop_prs2;
  wire        _slots_21_io_uop_bypassable;
  wire [4:0]  _slots_21_io_uop_mem_cmd;
  wire        _slots_21_io_uop_is_amo;
  wire        _slots_21_io_uop_uses_stq;
  wire        _slots_21_io_uop_ldst_val;
  wire [1:0]  _slots_21_io_uop_dst_rtype;
  wire [1:0]  _slots_21_io_uop_lrs1_rtype;
  wire [1:0]  _slots_21_io_uop_lrs2_rtype;
  wire        _slots_21_io_uop_fp_val;
  wire        _slots_20_io_valid;
  wire        _slots_20_io_will_be_valid;
  wire        _slots_20_io_request;
  wire [6:0]  _slots_20_io_out_uop_uopc;
  wire        _slots_20_io_out_uop_is_rvc;
  wire [9:0]  _slots_20_io_out_uop_fu_code;
  wire [1:0]  _slots_20_io_out_uop_iw_state;
  wire        _slots_20_io_out_uop_iw_p1_poisoned;
  wire        _slots_20_io_out_uop_iw_p2_poisoned;
  wire        _slots_20_io_out_uop_is_br;
  wire        _slots_20_io_out_uop_is_jalr;
  wire        _slots_20_io_out_uop_is_jal;
  wire        _slots_20_io_out_uop_is_sfb;
  wire [19:0] _slots_20_io_out_uop_br_mask;
  wire [4:0]  _slots_20_io_out_uop_br_tag;
  wire [5:0]  _slots_20_io_out_uop_ftq_idx;
  wire        _slots_20_io_out_uop_edge_inst;
  wire [5:0]  _slots_20_io_out_uop_pc_lob;
  wire        _slots_20_io_out_uop_taken;
  wire [19:0] _slots_20_io_out_uop_imm_packed;
  wire [6:0]  _slots_20_io_out_uop_rob_idx;
  wire [4:0]  _slots_20_io_out_uop_ldq_idx;
  wire [4:0]  _slots_20_io_out_uop_stq_idx;
  wire [6:0]  _slots_20_io_out_uop_pdst;
  wire [6:0]  _slots_20_io_out_uop_prs1;
  wire [6:0]  _slots_20_io_out_uop_prs2;
  wire [6:0]  _slots_20_io_out_uop_prs3;
  wire        _slots_20_io_out_uop_prs1_busy;
  wire        _slots_20_io_out_uop_prs2_busy;
  wire        _slots_20_io_out_uop_prs3_busy;
  wire        _slots_20_io_out_uop_ppred_busy;
  wire        _slots_20_io_out_uop_bypassable;
  wire [4:0]  _slots_20_io_out_uop_mem_cmd;
  wire [1:0]  _slots_20_io_out_uop_mem_size;
  wire        _slots_20_io_out_uop_mem_signed;
  wire        _slots_20_io_out_uop_is_fence;
  wire        _slots_20_io_out_uop_is_amo;
  wire        _slots_20_io_out_uop_uses_ldq;
  wire        _slots_20_io_out_uop_uses_stq;
  wire        _slots_20_io_out_uop_ldst_val;
  wire [1:0]  _slots_20_io_out_uop_dst_rtype;
  wire [1:0]  _slots_20_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_20_io_out_uop_lrs2_rtype;
  wire        _slots_20_io_out_uop_fp_val;
  wire [6:0]  _slots_20_io_uop_uopc;
  wire        _slots_20_io_uop_is_rvc;
  wire [9:0]  _slots_20_io_uop_fu_code;
  wire        _slots_20_io_uop_iw_p1_poisoned;
  wire        _slots_20_io_uop_iw_p2_poisoned;
  wire        _slots_20_io_uop_is_br;
  wire        _slots_20_io_uop_is_jalr;
  wire        _slots_20_io_uop_is_jal;
  wire        _slots_20_io_uop_is_sfb;
  wire [19:0] _slots_20_io_uop_br_mask;
  wire [4:0]  _slots_20_io_uop_br_tag;
  wire [5:0]  _slots_20_io_uop_ftq_idx;
  wire        _slots_20_io_uop_edge_inst;
  wire [5:0]  _slots_20_io_uop_pc_lob;
  wire        _slots_20_io_uop_taken;
  wire [19:0] _slots_20_io_uop_imm_packed;
  wire [6:0]  _slots_20_io_uop_rob_idx;
  wire [4:0]  _slots_20_io_uop_ldq_idx;
  wire [4:0]  _slots_20_io_uop_stq_idx;
  wire [6:0]  _slots_20_io_uop_pdst;
  wire [6:0]  _slots_20_io_uop_prs1;
  wire [6:0]  _slots_20_io_uop_prs2;
  wire        _slots_20_io_uop_bypassable;
  wire [4:0]  _slots_20_io_uop_mem_cmd;
  wire        _slots_20_io_uop_is_amo;
  wire        _slots_20_io_uop_uses_stq;
  wire        _slots_20_io_uop_ldst_val;
  wire [1:0]  _slots_20_io_uop_dst_rtype;
  wire [1:0]  _slots_20_io_uop_lrs1_rtype;
  wire [1:0]  _slots_20_io_uop_lrs2_rtype;
  wire        _slots_20_io_uop_fp_val;
  wire        _slots_19_io_valid;
  wire        _slots_19_io_will_be_valid;
  wire        _slots_19_io_request;
  wire [6:0]  _slots_19_io_out_uop_uopc;
  wire        _slots_19_io_out_uop_is_rvc;
  wire [9:0]  _slots_19_io_out_uop_fu_code;
  wire [1:0]  _slots_19_io_out_uop_iw_state;
  wire        _slots_19_io_out_uop_iw_p1_poisoned;
  wire        _slots_19_io_out_uop_iw_p2_poisoned;
  wire        _slots_19_io_out_uop_is_br;
  wire        _slots_19_io_out_uop_is_jalr;
  wire        _slots_19_io_out_uop_is_jal;
  wire        _slots_19_io_out_uop_is_sfb;
  wire [19:0] _slots_19_io_out_uop_br_mask;
  wire [4:0]  _slots_19_io_out_uop_br_tag;
  wire [5:0]  _slots_19_io_out_uop_ftq_idx;
  wire        _slots_19_io_out_uop_edge_inst;
  wire [5:0]  _slots_19_io_out_uop_pc_lob;
  wire        _slots_19_io_out_uop_taken;
  wire [19:0] _slots_19_io_out_uop_imm_packed;
  wire [6:0]  _slots_19_io_out_uop_rob_idx;
  wire [4:0]  _slots_19_io_out_uop_ldq_idx;
  wire [4:0]  _slots_19_io_out_uop_stq_idx;
  wire [6:0]  _slots_19_io_out_uop_pdst;
  wire [6:0]  _slots_19_io_out_uop_prs1;
  wire [6:0]  _slots_19_io_out_uop_prs2;
  wire [6:0]  _slots_19_io_out_uop_prs3;
  wire        _slots_19_io_out_uop_prs1_busy;
  wire        _slots_19_io_out_uop_prs2_busy;
  wire        _slots_19_io_out_uop_prs3_busy;
  wire        _slots_19_io_out_uop_ppred_busy;
  wire        _slots_19_io_out_uop_bypassable;
  wire [4:0]  _slots_19_io_out_uop_mem_cmd;
  wire [1:0]  _slots_19_io_out_uop_mem_size;
  wire        _slots_19_io_out_uop_mem_signed;
  wire        _slots_19_io_out_uop_is_fence;
  wire        _slots_19_io_out_uop_is_amo;
  wire        _slots_19_io_out_uop_uses_ldq;
  wire        _slots_19_io_out_uop_uses_stq;
  wire        _slots_19_io_out_uop_ldst_val;
  wire [1:0]  _slots_19_io_out_uop_dst_rtype;
  wire [1:0]  _slots_19_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_19_io_out_uop_lrs2_rtype;
  wire        _slots_19_io_out_uop_fp_val;
  wire [6:0]  _slots_19_io_uop_uopc;
  wire        _slots_19_io_uop_is_rvc;
  wire [9:0]  _slots_19_io_uop_fu_code;
  wire        _slots_19_io_uop_iw_p1_poisoned;
  wire        _slots_19_io_uop_iw_p2_poisoned;
  wire        _slots_19_io_uop_is_br;
  wire        _slots_19_io_uop_is_jalr;
  wire        _slots_19_io_uop_is_jal;
  wire        _slots_19_io_uop_is_sfb;
  wire [19:0] _slots_19_io_uop_br_mask;
  wire [4:0]  _slots_19_io_uop_br_tag;
  wire [5:0]  _slots_19_io_uop_ftq_idx;
  wire        _slots_19_io_uop_edge_inst;
  wire [5:0]  _slots_19_io_uop_pc_lob;
  wire        _slots_19_io_uop_taken;
  wire [19:0] _slots_19_io_uop_imm_packed;
  wire [6:0]  _slots_19_io_uop_rob_idx;
  wire [4:0]  _slots_19_io_uop_ldq_idx;
  wire [4:0]  _slots_19_io_uop_stq_idx;
  wire [6:0]  _slots_19_io_uop_pdst;
  wire [6:0]  _slots_19_io_uop_prs1;
  wire [6:0]  _slots_19_io_uop_prs2;
  wire        _slots_19_io_uop_bypassable;
  wire [4:0]  _slots_19_io_uop_mem_cmd;
  wire        _slots_19_io_uop_is_amo;
  wire        _slots_19_io_uop_uses_stq;
  wire        _slots_19_io_uop_ldst_val;
  wire [1:0]  _slots_19_io_uop_dst_rtype;
  wire [1:0]  _slots_19_io_uop_lrs1_rtype;
  wire [1:0]  _slots_19_io_uop_lrs2_rtype;
  wire        _slots_19_io_uop_fp_val;
  wire        _slots_18_io_valid;
  wire        _slots_18_io_will_be_valid;
  wire        _slots_18_io_request;
  wire [6:0]  _slots_18_io_out_uop_uopc;
  wire        _slots_18_io_out_uop_is_rvc;
  wire [9:0]  _slots_18_io_out_uop_fu_code;
  wire [1:0]  _slots_18_io_out_uop_iw_state;
  wire        _slots_18_io_out_uop_iw_p1_poisoned;
  wire        _slots_18_io_out_uop_iw_p2_poisoned;
  wire        _slots_18_io_out_uop_is_br;
  wire        _slots_18_io_out_uop_is_jalr;
  wire        _slots_18_io_out_uop_is_jal;
  wire        _slots_18_io_out_uop_is_sfb;
  wire [19:0] _slots_18_io_out_uop_br_mask;
  wire [4:0]  _slots_18_io_out_uop_br_tag;
  wire [5:0]  _slots_18_io_out_uop_ftq_idx;
  wire        _slots_18_io_out_uop_edge_inst;
  wire [5:0]  _slots_18_io_out_uop_pc_lob;
  wire        _slots_18_io_out_uop_taken;
  wire [19:0] _slots_18_io_out_uop_imm_packed;
  wire [6:0]  _slots_18_io_out_uop_rob_idx;
  wire [4:0]  _slots_18_io_out_uop_ldq_idx;
  wire [4:0]  _slots_18_io_out_uop_stq_idx;
  wire [6:0]  _slots_18_io_out_uop_pdst;
  wire [6:0]  _slots_18_io_out_uop_prs1;
  wire [6:0]  _slots_18_io_out_uop_prs2;
  wire [6:0]  _slots_18_io_out_uop_prs3;
  wire        _slots_18_io_out_uop_prs1_busy;
  wire        _slots_18_io_out_uop_prs2_busy;
  wire        _slots_18_io_out_uop_prs3_busy;
  wire        _slots_18_io_out_uop_ppred_busy;
  wire        _slots_18_io_out_uop_bypassable;
  wire [4:0]  _slots_18_io_out_uop_mem_cmd;
  wire [1:0]  _slots_18_io_out_uop_mem_size;
  wire        _slots_18_io_out_uop_mem_signed;
  wire        _slots_18_io_out_uop_is_fence;
  wire        _slots_18_io_out_uop_is_amo;
  wire        _slots_18_io_out_uop_uses_ldq;
  wire        _slots_18_io_out_uop_uses_stq;
  wire        _slots_18_io_out_uop_ldst_val;
  wire [1:0]  _slots_18_io_out_uop_dst_rtype;
  wire [1:0]  _slots_18_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_18_io_out_uop_lrs2_rtype;
  wire        _slots_18_io_out_uop_fp_val;
  wire [6:0]  _slots_18_io_uop_uopc;
  wire        _slots_18_io_uop_is_rvc;
  wire [9:0]  _slots_18_io_uop_fu_code;
  wire        _slots_18_io_uop_iw_p1_poisoned;
  wire        _slots_18_io_uop_iw_p2_poisoned;
  wire        _slots_18_io_uop_is_br;
  wire        _slots_18_io_uop_is_jalr;
  wire        _slots_18_io_uop_is_jal;
  wire        _slots_18_io_uop_is_sfb;
  wire [19:0] _slots_18_io_uop_br_mask;
  wire [4:0]  _slots_18_io_uop_br_tag;
  wire [5:0]  _slots_18_io_uop_ftq_idx;
  wire        _slots_18_io_uop_edge_inst;
  wire [5:0]  _slots_18_io_uop_pc_lob;
  wire        _slots_18_io_uop_taken;
  wire [19:0] _slots_18_io_uop_imm_packed;
  wire [6:0]  _slots_18_io_uop_rob_idx;
  wire [4:0]  _slots_18_io_uop_ldq_idx;
  wire [4:0]  _slots_18_io_uop_stq_idx;
  wire [6:0]  _slots_18_io_uop_pdst;
  wire [6:0]  _slots_18_io_uop_prs1;
  wire [6:0]  _slots_18_io_uop_prs2;
  wire        _slots_18_io_uop_bypassable;
  wire [4:0]  _slots_18_io_uop_mem_cmd;
  wire        _slots_18_io_uop_is_amo;
  wire        _slots_18_io_uop_uses_stq;
  wire        _slots_18_io_uop_ldst_val;
  wire [1:0]  _slots_18_io_uop_dst_rtype;
  wire [1:0]  _slots_18_io_uop_lrs1_rtype;
  wire [1:0]  _slots_18_io_uop_lrs2_rtype;
  wire        _slots_18_io_uop_fp_val;
  wire        _slots_17_io_valid;
  wire        _slots_17_io_will_be_valid;
  wire        _slots_17_io_request;
  wire [6:0]  _slots_17_io_out_uop_uopc;
  wire        _slots_17_io_out_uop_is_rvc;
  wire [9:0]  _slots_17_io_out_uop_fu_code;
  wire [1:0]  _slots_17_io_out_uop_iw_state;
  wire        _slots_17_io_out_uop_iw_p1_poisoned;
  wire        _slots_17_io_out_uop_iw_p2_poisoned;
  wire        _slots_17_io_out_uop_is_br;
  wire        _slots_17_io_out_uop_is_jalr;
  wire        _slots_17_io_out_uop_is_jal;
  wire        _slots_17_io_out_uop_is_sfb;
  wire [19:0] _slots_17_io_out_uop_br_mask;
  wire [4:0]  _slots_17_io_out_uop_br_tag;
  wire [5:0]  _slots_17_io_out_uop_ftq_idx;
  wire        _slots_17_io_out_uop_edge_inst;
  wire [5:0]  _slots_17_io_out_uop_pc_lob;
  wire        _slots_17_io_out_uop_taken;
  wire [19:0] _slots_17_io_out_uop_imm_packed;
  wire [6:0]  _slots_17_io_out_uop_rob_idx;
  wire [4:0]  _slots_17_io_out_uop_ldq_idx;
  wire [4:0]  _slots_17_io_out_uop_stq_idx;
  wire [6:0]  _slots_17_io_out_uop_pdst;
  wire [6:0]  _slots_17_io_out_uop_prs1;
  wire [6:0]  _slots_17_io_out_uop_prs2;
  wire [6:0]  _slots_17_io_out_uop_prs3;
  wire        _slots_17_io_out_uop_prs1_busy;
  wire        _slots_17_io_out_uop_prs2_busy;
  wire        _slots_17_io_out_uop_prs3_busy;
  wire        _slots_17_io_out_uop_ppred_busy;
  wire        _slots_17_io_out_uop_bypassable;
  wire [4:0]  _slots_17_io_out_uop_mem_cmd;
  wire [1:0]  _slots_17_io_out_uop_mem_size;
  wire        _slots_17_io_out_uop_mem_signed;
  wire        _slots_17_io_out_uop_is_fence;
  wire        _slots_17_io_out_uop_is_amo;
  wire        _slots_17_io_out_uop_uses_ldq;
  wire        _slots_17_io_out_uop_uses_stq;
  wire        _slots_17_io_out_uop_ldst_val;
  wire [1:0]  _slots_17_io_out_uop_dst_rtype;
  wire [1:0]  _slots_17_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_17_io_out_uop_lrs2_rtype;
  wire        _slots_17_io_out_uop_fp_val;
  wire [6:0]  _slots_17_io_uop_uopc;
  wire        _slots_17_io_uop_is_rvc;
  wire [9:0]  _slots_17_io_uop_fu_code;
  wire        _slots_17_io_uop_iw_p1_poisoned;
  wire        _slots_17_io_uop_iw_p2_poisoned;
  wire        _slots_17_io_uop_is_br;
  wire        _slots_17_io_uop_is_jalr;
  wire        _slots_17_io_uop_is_jal;
  wire        _slots_17_io_uop_is_sfb;
  wire [19:0] _slots_17_io_uop_br_mask;
  wire [4:0]  _slots_17_io_uop_br_tag;
  wire [5:0]  _slots_17_io_uop_ftq_idx;
  wire        _slots_17_io_uop_edge_inst;
  wire [5:0]  _slots_17_io_uop_pc_lob;
  wire        _slots_17_io_uop_taken;
  wire [19:0] _slots_17_io_uop_imm_packed;
  wire [6:0]  _slots_17_io_uop_rob_idx;
  wire [4:0]  _slots_17_io_uop_ldq_idx;
  wire [4:0]  _slots_17_io_uop_stq_idx;
  wire [6:0]  _slots_17_io_uop_pdst;
  wire [6:0]  _slots_17_io_uop_prs1;
  wire [6:0]  _slots_17_io_uop_prs2;
  wire        _slots_17_io_uop_bypassable;
  wire [4:0]  _slots_17_io_uop_mem_cmd;
  wire        _slots_17_io_uop_is_amo;
  wire        _slots_17_io_uop_uses_stq;
  wire        _slots_17_io_uop_ldst_val;
  wire [1:0]  _slots_17_io_uop_dst_rtype;
  wire [1:0]  _slots_17_io_uop_lrs1_rtype;
  wire [1:0]  _slots_17_io_uop_lrs2_rtype;
  wire        _slots_17_io_uop_fp_val;
  wire        _slots_16_io_valid;
  wire        _slots_16_io_will_be_valid;
  wire        _slots_16_io_request;
  wire [6:0]  _slots_16_io_out_uop_uopc;
  wire        _slots_16_io_out_uop_is_rvc;
  wire [9:0]  _slots_16_io_out_uop_fu_code;
  wire [1:0]  _slots_16_io_out_uop_iw_state;
  wire        _slots_16_io_out_uop_iw_p1_poisoned;
  wire        _slots_16_io_out_uop_iw_p2_poisoned;
  wire        _slots_16_io_out_uop_is_br;
  wire        _slots_16_io_out_uop_is_jalr;
  wire        _slots_16_io_out_uop_is_jal;
  wire        _slots_16_io_out_uop_is_sfb;
  wire [19:0] _slots_16_io_out_uop_br_mask;
  wire [4:0]  _slots_16_io_out_uop_br_tag;
  wire [5:0]  _slots_16_io_out_uop_ftq_idx;
  wire        _slots_16_io_out_uop_edge_inst;
  wire [5:0]  _slots_16_io_out_uop_pc_lob;
  wire        _slots_16_io_out_uop_taken;
  wire [19:0] _slots_16_io_out_uop_imm_packed;
  wire [6:0]  _slots_16_io_out_uop_rob_idx;
  wire [4:0]  _slots_16_io_out_uop_ldq_idx;
  wire [4:0]  _slots_16_io_out_uop_stq_idx;
  wire [6:0]  _slots_16_io_out_uop_pdst;
  wire [6:0]  _slots_16_io_out_uop_prs1;
  wire [6:0]  _slots_16_io_out_uop_prs2;
  wire [6:0]  _slots_16_io_out_uop_prs3;
  wire        _slots_16_io_out_uop_prs1_busy;
  wire        _slots_16_io_out_uop_prs2_busy;
  wire        _slots_16_io_out_uop_prs3_busy;
  wire        _slots_16_io_out_uop_ppred_busy;
  wire        _slots_16_io_out_uop_bypassable;
  wire [4:0]  _slots_16_io_out_uop_mem_cmd;
  wire [1:0]  _slots_16_io_out_uop_mem_size;
  wire        _slots_16_io_out_uop_mem_signed;
  wire        _slots_16_io_out_uop_is_fence;
  wire        _slots_16_io_out_uop_is_amo;
  wire        _slots_16_io_out_uop_uses_ldq;
  wire        _slots_16_io_out_uop_uses_stq;
  wire        _slots_16_io_out_uop_ldst_val;
  wire [1:0]  _slots_16_io_out_uop_dst_rtype;
  wire [1:0]  _slots_16_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_16_io_out_uop_lrs2_rtype;
  wire        _slots_16_io_out_uop_fp_val;
  wire [6:0]  _slots_16_io_uop_uopc;
  wire        _slots_16_io_uop_is_rvc;
  wire [9:0]  _slots_16_io_uop_fu_code;
  wire        _slots_16_io_uop_iw_p1_poisoned;
  wire        _slots_16_io_uop_iw_p2_poisoned;
  wire        _slots_16_io_uop_is_br;
  wire        _slots_16_io_uop_is_jalr;
  wire        _slots_16_io_uop_is_jal;
  wire        _slots_16_io_uop_is_sfb;
  wire [19:0] _slots_16_io_uop_br_mask;
  wire [4:0]  _slots_16_io_uop_br_tag;
  wire [5:0]  _slots_16_io_uop_ftq_idx;
  wire        _slots_16_io_uop_edge_inst;
  wire [5:0]  _slots_16_io_uop_pc_lob;
  wire        _slots_16_io_uop_taken;
  wire [19:0] _slots_16_io_uop_imm_packed;
  wire [6:0]  _slots_16_io_uop_rob_idx;
  wire [4:0]  _slots_16_io_uop_ldq_idx;
  wire [4:0]  _slots_16_io_uop_stq_idx;
  wire [6:0]  _slots_16_io_uop_pdst;
  wire [6:0]  _slots_16_io_uop_prs1;
  wire [6:0]  _slots_16_io_uop_prs2;
  wire        _slots_16_io_uop_bypassable;
  wire [4:0]  _slots_16_io_uop_mem_cmd;
  wire        _slots_16_io_uop_is_amo;
  wire        _slots_16_io_uop_uses_stq;
  wire        _slots_16_io_uop_ldst_val;
  wire [1:0]  _slots_16_io_uop_dst_rtype;
  wire [1:0]  _slots_16_io_uop_lrs1_rtype;
  wire [1:0]  _slots_16_io_uop_lrs2_rtype;
  wire        _slots_16_io_uop_fp_val;
  wire        _slots_15_io_valid;
  wire        _slots_15_io_will_be_valid;
  wire        _slots_15_io_request;
  wire [6:0]  _slots_15_io_out_uop_uopc;
  wire        _slots_15_io_out_uop_is_rvc;
  wire [9:0]  _slots_15_io_out_uop_fu_code;
  wire [1:0]  _slots_15_io_out_uop_iw_state;
  wire        _slots_15_io_out_uop_iw_p1_poisoned;
  wire        _slots_15_io_out_uop_iw_p2_poisoned;
  wire        _slots_15_io_out_uop_is_br;
  wire        _slots_15_io_out_uop_is_jalr;
  wire        _slots_15_io_out_uop_is_jal;
  wire        _slots_15_io_out_uop_is_sfb;
  wire [19:0] _slots_15_io_out_uop_br_mask;
  wire [4:0]  _slots_15_io_out_uop_br_tag;
  wire [5:0]  _slots_15_io_out_uop_ftq_idx;
  wire        _slots_15_io_out_uop_edge_inst;
  wire [5:0]  _slots_15_io_out_uop_pc_lob;
  wire        _slots_15_io_out_uop_taken;
  wire [19:0] _slots_15_io_out_uop_imm_packed;
  wire [6:0]  _slots_15_io_out_uop_rob_idx;
  wire [4:0]  _slots_15_io_out_uop_ldq_idx;
  wire [4:0]  _slots_15_io_out_uop_stq_idx;
  wire [6:0]  _slots_15_io_out_uop_pdst;
  wire [6:0]  _slots_15_io_out_uop_prs1;
  wire [6:0]  _slots_15_io_out_uop_prs2;
  wire [6:0]  _slots_15_io_out_uop_prs3;
  wire        _slots_15_io_out_uop_prs1_busy;
  wire        _slots_15_io_out_uop_prs2_busy;
  wire        _slots_15_io_out_uop_prs3_busy;
  wire        _slots_15_io_out_uop_ppred_busy;
  wire        _slots_15_io_out_uop_bypassable;
  wire [4:0]  _slots_15_io_out_uop_mem_cmd;
  wire [1:0]  _slots_15_io_out_uop_mem_size;
  wire        _slots_15_io_out_uop_mem_signed;
  wire        _slots_15_io_out_uop_is_fence;
  wire        _slots_15_io_out_uop_is_amo;
  wire        _slots_15_io_out_uop_uses_ldq;
  wire        _slots_15_io_out_uop_uses_stq;
  wire        _slots_15_io_out_uop_ldst_val;
  wire [1:0]  _slots_15_io_out_uop_dst_rtype;
  wire [1:0]  _slots_15_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_15_io_out_uop_lrs2_rtype;
  wire        _slots_15_io_out_uop_fp_val;
  wire [6:0]  _slots_15_io_uop_uopc;
  wire        _slots_15_io_uop_is_rvc;
  wire [9:0]  _slots_15_io_uop_fu_code;
  wire        _slots_15_io_uop_iw_p1_poisoned;
  wire        _slots_15_io_uop_iw_p2_poisoned;
  wire        _slots_15_io_uop_is_br;
  wire        _slots_15_io_uop_is_jalr;
  wire        _slots_15_io_uop_is_jal;
  wire        _slots_15_io_uop_is_sfb;
  wire [19:0] _slots_15_io_uop_br_mask;
  wire [4:0]  _slots_15_io_uop_br_tag;
  wire [5:0]  _slots_15_io_uop_ftq_idx;
  wire        _slots_15_io_uop_edge_inst;
  wire [5:0]  _slots_15_io_uop_pc_lob;
  wire        _slots_15_io_uop_taken;
  wire [19:0] _slots_15_io_uop_imm_packed;
  wire [6:0]  _slots_15_io_uop_rob_idx;
  wire [4:0]  _slots_15_io_uop_ldq_idx;
  wire [4:0]  _slots_15_io_uop_stq_idx;
  wire [6:0]  _slots_15_io_uop_pdst;
  wire [6:0]  _slots_15_io_uop_prs1;
  wire [6:0]  _slots_15_io_uop_prs2;
  wire        _slots_15_io_uop_bypassable;
  wire [4:0]  _slots_15_io_uop_mem_cmd;
  wire        _slots_15_io_uop_is_amo;
  wire        _slots_15_io_uop_uses_stq;
  wire        _slots_15_io_uop_ldst_val;
  wire [1:0]  _slots_15_io_uop_dst_rtype;
  wire [1:0]  _slots_15_io_uop_lrs1_rtype;
  wire [1:0]  _slots_15_io_uop_lrs2_rtype;
  wire        _slots_15_io_uop_fp_val;
  wire        _slots_14_io_valid;
  wire        _slots_14_io_will_be_valid;
  wire        _slots_14_io_request;
  wire [6:0]  _slots_14_io_out_uop_uopc;
  wire        _slots_14_io_out_uop_is_rvc;
  wire [9:0]  _slots_14_io_out_uop_fu_code;
  wire [1:0]  _slots_14_io_out_uop_iw_state;
  wire        _slots_14_io_out_uop_iw_p1_poisoned;
  wire        _slots_14_io_out_uop_iw_p2_poisoned;
  wire        _slots_14_io_out_uop_is_br;
  wire        _slots_14_io_out_uop_is_jalr;
  wire        _slots_14_io_out_uop_is_jal;
  wire        _slots_14_io_out_uop_is_sfb;
  wire [19:0] _slots_14_io_out_uop_br_mask;
  wire [4:0]  _slots_14_io_out_uop_br_tag;
  wire [5:0]  _slots_14_io_out_uop_ftq_idx;
  wire        _slots_14_io_out_uop_edge_inst;
  wire [5:0]  _slots_14_io_out_uop_pc_lob;
  wire        _slots_14_io_out_uop_taken;
  wire [19:0] _slots_14_io_out_uop_imm_packed;
  wire [6:0]  _slots_14_io_out_uop_rob_idx;
  wire [4:0]  _slots_14_io_out_uop_ldq_idx;
  wire [4:0]  _slots_14_io_out_uop_stq_idx;
  wire [6:0]  _slots_14_io_out_uop_pdst;
  wire [6:0]  _slots_14_io_out_uop_prs1;
  wire [6:0]  _slots_14_io_out_uop_prs2;
  wire [6:0]  _slots_14_io_out_uop_prs3;
  wire        _slots_14_io_out_uop_prs1_busy;
  wire        _slots_14_io_out_uop_prs2_busy;
  wire        _slots_14_io_out_uop_prs3_busy;
  wire        _slots_14_io_out_uop_ppred_busy;
  wire        _slots_14_io_out_uop_bypassable;
  wire [4:0]  _slots_14_io_out_uop_mem_cmd;
  wire [1:0]  _slots_14_io_out_uop_mem_size;
  wire        _slots_14_io_out_uop_mem_signed;
  wire        _slots_14_io_out_uop_is_fence;
  wire        _slots_14_io_out_uop_is_amo;
  wire        _slots_14_io_out_uop_uses_ldq;
  wire        _slots_14_io_out_uop_uses_stq;
  wire        _slots_14_io_out_uop_ldst_val;
  wire [1:0]  _slots_14_io_out_uop_dst_rtype;
  wire [1:0]  _slots_14_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_14_io_out_uop_lrs2_rtype;
  wire        _slots_14_io_out_uop_fp_val;
  wire [6:0]  _slots_14_io_uop_uopc;
  wire        _slots_14_io_uop_is_rvc;
  wire [9:0]  _slots_14_io_uop_fu_code;
  wire        _slots_14_io_uop_iw_p1_poisoned;
  wire        _slots_14_io_uop_iw_p2_poisoned;
  wire        _slots_14_io_uop_is_br;
  wire        _slots_14_io_uop_is_jalr;
  wire        _slots_14_io_uop_is_jal;
  wire        _slots_14_io_uop_is_sfb;
  wire [19:0] _slots_14_io_uop_br_mask;
  wire [4:0]  _slots_14_io_uop_br_tag;
  wire [5:0]  _slots_14_io_uop_ftq_idx;
  wire        _slots_14_io_uop_edge_inst;
  wire [5:0]  _slots_14_io_uop_pc_lob;
  wire        _slots_14_io_uop_taken;
  wire [19:0] _slots_14_io_uop_imm_packed;
  wire [6:0]  _slots_14_io_uop_rob_idx;
  wire [4:0]  _slots_14_io_uop_ldq_idx;
  wire [4:0]  _slots_14_io_uop_stq_idx;
  wire [6:0]  _slots_14_io_uop_pdst;
  wire [6:0]  _slots_14_io_uop_prs1;
  wire [6:0]  _slots_14_io_uop_prs2;
  wire        _slots_14_io_uop_bypassable;
  wire [4:0]  _slots_14_io_uop_mem_cmd;
  wire        _slots_14_io_uop_is_amo;
  wire        _slots_14_io_uop_uses_stq;
  wire        _slots_14_io_uop_ldst_val;
  wire [1:0]  _slots_14_io_uop_dst_rtype;
  wire [1:0]  _slots_14_io_uop_lrs1_rtype;
  wire [1:0]  _slots_14_io_uop_lrs2_rtype;
  wire        _slots_14_io_uop_fp_val;
  wire        _slots_13_io_valid;
  wire        _slots_13_io_will_be_valid;
  wire        _slots_13_io_request;
  wire [6:0]  _slots_13_io_out_uop_uopc;
  wire        _slots_13_io_out_uop_is_rvc;
  wire [9:0]  _slots_13_io_out_uop_fu_code;
  wire [1:0]  _slots_13_io_out_uop_iw_state;
  wire        _slots_13_io_out_uop_iw_p1_poisoned;
  wire        _slots_13_io_out_uop_iw_p2_poisoned;
  wire        _slots_13_io_out_uop_is_br;
  wire        _slots_13_io_out_uop_is_jalr;
  wire        _slots_13_io_out_uop_is_jal;
  wire        _slots_13_io_out_uop_is_sfb;
  wire [19:0] _slots_13_io_out_uop_br_mask;
  wire [4:0]  _slots_13_io_out_uop_br_tag;
  wire [5:0]  _slots_13_io_out_uop_ftq_idx;
  wire        _slots_13_io_out_uop_edge_inst;
  wire [5:0]  _slots_13_io_out_uop_pc_lob;
  wire        _slots_13_io_out_uop_taken;
  wire [19:0] _slots_13_io_out_uop_imm_packed;
  wire [6:0]  _slots_13_io_out_uop_rob_idx;
  wire [4:0]  _slots_13_io_out_uop_ldq_idx;
  wire [4:0]  _slots_13_io_out_uop_stq_idx;
  wire [6:0]  _slots_13_io_out_uop_pdst;
  wire [6:0]  _slots_13_io_out_uop_prs1;
  wire [6:0]  _slots_13_io_out_uop_prs2;
  wire [6:0]  _slots_13_io_out_uop_prs3;
  wire        _slots_13_io_out_uop_prs1_busy;
  wire        _slots_13_io_out_uop_prs2_busy;
  wire        _slots_13_io_out_uop_prs3_busy;
  wire        _slots_13_io_out_uop_ppred_busy;
  wire        _slots_13_io_out_uop_bypassable;
  wire [4:0]  _slots_13_io_out_uop_mem_cmd;
  wire [1:0]  _slots_13_io_out_uop_mem_size;
  wire        _slots_13_io_out_uop_mem_signed;
  wire        _slots_13_io_out_uop_is_fence;
  wire        _slots_13_io_out_uop_is_amo;
  wire        _slots_13_io_out_uop_uses_ldq;
  wire        _slots_13_io_out_uop_uses_stq;
  wire        _slots_13_io_out_uop_ldst_val;
  wire [1:0]  _slots_13_io_out_uop_dst_rtype;
  wire [1:0]  _slots_13_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_13_io_out_uop_lrs2_rtype;
  wire        _slots_13_io_out_uop_fp_val;
  wire [6:0]  _slots_13_io_uop_uopc;
  wire        _slots_13_io_uop_is_rvc;
  wire [9:0]  _slots_13_io_uop_fu_code;
  wire        _slots_13_io_uop_iw_p1_poisoned;
  wire        _slots_13_io_uop_iw_p2_poisoned;
  wire        _slots_13_io_uop_is_br;
  wire        _slots_13_io_uop_is_jalr;
  wire        _slots_13_io_uop_is_jal;
  wire        _slots_13_io_uop_is_sfb;
  wire [19:0] _slots_13_io_uop_br_mask;
  wire [4:0]  _slots_13_io_uop_br_tag;
  wire [5:0]  _slots_13_io_uop_ftq_idx;
  wire        _slots_13_io_uop_edge_inst;
  wire [5:0]  _slots_13_io_uop_pc_lob;
  wire        _slots_13_io_uop_taken;
  wire [19:0] _slots_13_io_uop_imm_packed;
  wire [6:0]  _slots_13_io_uop_rob_idx;
  wire [4:0]  _slots_13_io_uop_ldq_idx;
  wire [4:0]  _slots_13_io_uop_stq_idx;
  wire [6:0]  _slots_13_io_uop_pdst;
  wire [6:0]  _slots_13_io_uop_prs1;
  wire [6:0]  _slots_13_io_uop_prs2;
  wire        _slots_13_io_uop_bypassable;
  wire [4:0]  _slots_13_io_uop_mem_cmd;
  wire        _slots_13_io_uop_is_amo;
  wire        _slots_13_io_uop_uses_stq;
  wire        _slots_13_io_uop_ldst_val;
  wire [1:0]  _slots_13_io_uop_dst_rtype;
  wire [1:0]  _slots_13_io_uop_lrs1_rtype;
  wire [1:0]  _slots_13_io_uop_lrs2_rtype;
  wire        _slots_13_io_uop_fp_val;
  wire        _slots_12_io_valid;
  wire        _slots_12_io_will_be_valid;
  wire        _slots_12_io_request;
  wire [6:0]  _slots_12_io_out_uop_uopc;
  wire        _slots_12_io_out_uop_is_rvc;
  wire [9:0]  _slots_12_io_out_uop_fu_code;
  wire [1:0]  _slots_12_io_out_uop_iw_state;
  wire        _slots_12_io_out_uop_iw_p1_poisoned;
  wire        _slots_12_io_out_uop_iw_p2_poisoned;
  wire        _slots_12_io_out_uop_is_br;
  wire        _slots_12_io_out_uop_is_jalr;
  wire        _slots_12_io_out_uop_is_jal;
  wire        _slots_12_io_out_uop_is_sfb;
  wire [19:0] _slots_12_io_out_uop_br_mask;
  wire [4:0]  _slots_12_io_out_uop_br_tag;
  wire [5:0]  _slots_12_io_out_uop_ftq_idx;
  wire        _slots_12_io_out_uop_edge_inst;
  wire [5:0]  _slots_12_io_out_uop_pc_lob;
  wire        _slots_12_io_out_uop_taken;
  wire [19:0] _slots_12_io_out_uop_imm_packed;
  wire [6:0]  _slots_12_io_out_uop_rob_idx;
  wire [4:0]  _slots_12_io_out_uop_ldq_idx;
  wire [4:0]  _slots_12_io_out_uop_stq_idx;
  wire [6:0]  _slots_12_io_out_uop_pdst;
  wire [6:0]  _slots_12_io_out_uop_prs1;
  wire [6:0]  _slots_12_io_out_uop_prs2;
  wire [6:0]  _slots_12_io_out_uop_prs3;
  wire        _slots_12_io_out_uop_prs1_busy;
  wire        _slots_12_io_out_uop_prs2_busy;
  wire        _slots_12_io_out_uop_prs3_busy;
  wire        _slots_12_io_out_uop_ppred_busy;
  wire        _slots_12_io_out_uop_bypassable;
  wire [4:0]  _slots_12_io_out_uop_mem_cmd;
  wire [1:0]  _slots_12_io_out_uop_mem_size;
  wire        _slots_12_io_out_uop_mem_signed;
  wire        _slots_12_io_out_uop_is_fence;
  wire        _slots_12_io_out_uop_is_amo;
  wire        _slots_12_io_out_uop_uses_ldq;
  wire        _slots_12_io_out_uop_uses_stq;
  wire        _slots_12_io_out_uop_ldst_val;
  wire [1:0]  _slots_12_io_out_uop_dst_rtype;
  wire [1:0]  _slots_12_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_12_io_out_uop_lrs2_rtype;
  wire        _slots_12_io_out_uop_fp_val;
  wire [6:0]  _slots_12_io_uop_uopc;
  wire        _slots_12_io_uop_is_rvc;
  wire [9:0]  _slots_12_io_uop_fu_code;
  wire        _slots_12_io_uop_iw_p1_poisoned;
  wire        _slots_12_io_uop_iw_p2_poisoned;
  wire        _slots_12_io_uop_is_br;
  wire        _slots_12_io_uop_is_jalr;
  wire        _slots_12_io_uop_is_jal;
  wire        _slots_12_io_uop_is_sfb;
  wire [19:0] _slots_12_io_uop_br_mask;
  wire [4:0]  _slots_12_io_uop_br_tag;
  wire [5:0]  _slots_12_io_uop_ftq_idx;
  wire        _slots_12_io_uop_edge_inst;
  wire [5:0]  _slots_12_io_uop_pc_lob;
  wire        _slots_12_io_uop_taken;
  wire [19:0] _slots_12_io_uop_imm_packed;
  wire [6:0]  _slots_12_io_uop_rob_idx;
  wire [4:0]  _slots_12_io_uop_ldq_idx;
  wire [4:0]  _slots_12_io_uop_stq_idx;
  wire [6:0]  _slots_12_io_uop_pdst;
  wire [6:0]  _slots_12_io_uop_prs1;
  wire [6:0]  _slots_12_io_uop_prs2;
  wire        _slots_12_io_uop_bypassable;
  wire [4:0]  _slots_12_io_uop_mem_cmd;
  wire        _slots_12_io_uop_is_amo;
  wire        _slots_12_io_uop_uses_stq;
  wire        _slots_12_io_uop_ldst_val;
  wire [1:0]  _slots_12_io_uop_dst_rtype;
  wire [1:0]  _slots_12_io_uop_lrs1_rtype;
  wire [1:0]  _slots_12_io_uop_lrs2_rtype;
  wire        _slots_12_io_uop_fp_val;
  wire        _slots_11_io_valid;
  wire        _slots_11_io_will_be_valid;
  wire        _slots_11_io_request;
  wire [6:0]  _slots_11_io_out_uop_uopc;
  wire        _slots_11_io_out_uop_is_rvc;
  wire [9:0]  _slots_11_io_out_uop_fu_code;
  wire [1:0]  _slots_11_io_out_uop_iw_state;
  wire        _slots_11_io_out_uop_iw_p1_poisoned;
  wire        _slots_11_io_out_uop_iw_p2_poisoned;
  wire        _slots_11_io_out_uop_is_br;
  wire        _slots_11_io_out_uop_is_jalr;
  wire        _slots_11_io_out_uop_is_jal;
  wire        _slots_11_io_out_uop_is_sfb;
  wire [19:0] _slots_11_io_out_uop_br_mask;
  wire [4:0]  _slots_11_io_out_uop_br_tag;
  wire [5:0]  _slots_11_io_out_uop_ftq_idx;
  wire        _slots_11_io_out_uop_edge_inst;
  wire [5:0]  _slots_11_io_out_uop_pc_lob;
  wire        _slots_11_io_out_uop_taken;
  wire [19:0] _slots_11_io_out_uop_imm_packed;
  wire [6:0]  _slots_11_io_out_uop_rob_idx;
  wire [4:0]  _slots_11_io_out_uop_ldq_idx;
  wire [4:0]  _slots_11_io_out_uop_stq_idx;
  wire [6:0]  _slots_11_io_out_uop_pdst;
  wire [6:0]  _slots_11_io_out_uop_prs1;
  wire [6:0]  _slots_11_io_out_uop_prs2;
  wire [6:0]  _slots_11_io_out_uop_prs3;
  wire        _slots_11_io_out_uop_prs1_busy;
  wire        _slots_11_io_out_uop_prs2_busy;
  wire        _slots_11_io_out_uop_prs3_busy;
  wire        _slots_11_io_out_uop_ppred_busy;
  wire        _slots_11_io_out_uop_bypassable;
  wire [4:0]  _slots_11_io_out_uop_mem_cmd;
  wire [1:0]  _slots_11_io_out_uop_mem_size;
  wire        _slots_11_io_out_uop_mem_signed;
  wire        _slots_11_io_out_uop_is_fence;
  wire        _slots_11_io_out_uop_is_amo;
  wire        _slots_11_io_out_uop_uses_ldq;
  wire        _slots_11_io_out_uop_uses_stq;
  wire        _slots_11_io_out_uop_ldst_val;
  wire [1:0]  _slots_11_io_out_uop_dst_rtype;
  wire [1:0]  _slots_11_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_11_io_out_uop_lrs2_rtype;
  wire        _slots_11_io_out_uop_fp_val;
  wire [6:0]  _slots_11_io_uop_uopc;
  wire        _slots_11_io_uop_is_rvc;
  wire [9:0]  _slots_11_io_uop_fu_code;
  wire        _slots_11_io_uop_iw_p1_poisoned;
  wire        _slots_11_io_uop_iw_p2_poisoned;
  wire        _slots_11_io_uop_is_br;
  wire        _slots_11_io_uop_is_jalr;
  wire        _slots_11_io_uop_is_jal;
  wire        _slots_11_io_uop_is_sfb;
  wire [19:0] _slots_11_io_uop_br_mask;
  wire [4:0]  _slots_11_io_uop_br_tag;
  wire [5:0]  _slots_11_io_uop_ftq_idx;
  wire        _slots_11_io_uop_edge_inst;
  wire [5:0]  _slots_11_io_uop_pc_lob;
  wire        _slots_11_io_uop_taken;
  wire [19:0] _slots_11_io_uop_imm_packed;
  wire [6:0]  _slots_11_io_uop_rob_idx;
  wire [4:0]  _slots_11_io_uop_ldq_idx;
  wire [4:0]  _slots_11_io_uop_stq_idx;
  wire [6:0]  _slots_11_io_uop_pdst;
  wire [6:0]  _slots_11_io_uop_prs1;
  wire [6:0]  _slots_11_io_uop_prs2;
  wire        _slots_11_io_uop_bypassable;
  wire [4:0]  _slots_11_io_uop_mem_cmd;
  wire        _slots_11_io_uop_is_amo;
  wire        _slots_11_io_uop_uses_stq;
  wire        _slots_11_io_uop_ldst_val;
  wire [1:0]  _slots_11_io_uop_dst_rtype;
  wire [1:0]  _slots_11_io_uop_lrs1_rtype;
  wire [1:0]  _slots_11_io_uop_lrs2_rtype;
  wire        _slots_11_io_uop_fp_val;
  wire        _slots_10_io_valid;
  wire        _slots_10_io_will_be_valid;
  wire        _slots_10_io_request;
  wire [6:0]  _slots_10_io_out_uop_uopc;
  wire        _slots_10_io_out_uop_is_rvc;
  wire [9:0]  _slots_10_io_out_uop_fu_code;
  wire [1:0]  _slots_10_io_out_uop_iw_state;
  wire        _slots_10_io_out_uop_iw_p1_poisoned;
  wire        _slots_10_io_out_uop_iw_p2_poisoned;
  wire        _slots_10_io_out_uop_is_br;
  wire        _slots_10_io_out_uop_is_jalr;
  wire        _slots_10_io_out_uop_is_jal;
  wire        _slots_10_io_out_uop_is_sfb;
  wire [19:0] _slots_10_io_out_uop_br_mask;
  wire [4:0]  _slots_10_io_out_uop_br_tag;
  wire [5:0]  _slots_10_io_out_uop_ftq_idx;
  wire        _slots_10_io_out_uop_edge_inst;
  wire [5:0]  _slots_10_io_out_uop_pc_lob;
  wire        _slots_10_io_out_uop_taken;
  wire [19:0] _slots_10_io_out_uop_imm_packed;
  wire [6:0]  _slots_10_io_out_uop_rob_idx;
  wire [4:0]  _slots_10_io_out_uop_ldq_idx;
  wire [4:0]  _slots_10_io_out_uop_stq_idx;
  wire [6:0]  _slots_10_io_out_uop_pdst;
  wire [6:0]  _slots_10_io_out_uop_prs1;
  wire [6:0]  _slots_10_io_out_uop_prs2;
  wire [6:0]  _slots_10_io_out_uop_prs3;
  wire        _slots_10_io_out_uop_prs1_busy;
  wire        _slots_10_io_out_uop_prs2_busy;
  wire        _slots_10_io_out_uop_prs3_busy;
  wire        _slots_10_io_out_uop_ppred_busy;
  wire        _slots_10_io_out_uop_bypassable;
  wire [4:0]  _slots_10_io_out_uop_mem_cmd;
  wire [1:0]  _slots_10_io_out_uop_mem_size;
  wire        _slots_10_io_out_uop_mem_signed;
  wire        _slots_10_io_out_uop_is_fence;
  wire        _slots_10_io_out_uop_is_amo;
  wire        _slots_10_io_out_uop_uses_ldq;
  wire        _slots_10_io_out_uop_uses_stq;
  wire        _slots_10_io_out_uop_ldst_val;
  wire [1:0]  _slots_10_io_out_uop_dst_rtype;
  wire [1:0]  _slots_10_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_10_io_out_uop_lrs2_rtype;
  wire        _slots_10_io_out_uop_fp_val;
  wire [6:0]  _slots_10_io_uop_uopc;
  wire        _slots_10_io_uop_is_rvc;
  wire [9:0]  _slots_10_io_uop_fu_code;
  wire        _slots_10_io_uop_iw_p1_poisoned;
  wire        _slots_10_io_uop_iw_p2_poisoned;
  wire        _slots_10_io_uop_is_br;
  wire        _slots_10_io_uop_is_jalr;
  wire        _slots_10_io_uop_is_jal;
  wire        _slots_10_io_uop_is_sfb;
  wire [19:0] _slots_10_io_uop_br_mask;
  wire [4:0]  _slots_10_io_uop_br_tag;
  wire [5:0]  _slots_10_io_uop_ftq_idx;
  wire        _slots_10_io_uop_edge_inst;
  wire [5:0]  _slots_10_io_uop_pc_lob;
  wire        _slots_10_io_uop_taken;
  wire [19:0] _slots_10_io_uop_imm_packed;
  wire [6:0]  _slots_10_io_uop_rob_idx;
  wire [4:0]  _slots_10_io_uop_ldq_idx;
  wire [4:0]  _slots_10_io_uop_stq_idx;
  wire [6:0]  _slots_10_io_uop_pdst;
  wire [6:0]  _slots_10_io_uop_prs1;
  wire [6:0]  _slots_10_io_uop_prs2;
  wire        _slots_10_io_uop_bypassable;
  wire [4:0]  _slots_10_io_uop_mem_cmd;
  wire        _slots_10_io_uop_is_amo;
  wire        _slots_10_io_uop_uses_stq;
  wire        _slots_10_io_uop_ldst_val;
  wire [1:0]  _slots_10_io_uop_dst_rtype;
  wire [1:0]  _slots_10_io_uop_lrs1_rtype;
  wire [1:0]  _slots_10_io_uop_lrs2_rtype;
  wire        _slots_10_io_uop_fp_val;
  wire        _slots_9_io_valid;
  wire        _slots_9_io_will_be_valid;
  wire        _slots_9_io_request;
  wire [6:0]  _slots_9_io_out_uop_uopc;
  wire        _slots_9_io_out_uop_is_rvc;
  wire [9:0]  _slots_9_io_out_uop_fu_code;
  wire [1:0]  _slots_9_io_out_uop_iw_state;
  wire        _slots_9_io_out_uop_iw_p1_poisoned;
  wire        _slots_9_io_out_uop_iw_p2_poisoned;
  wire        _slots_9_io_out_uop_is_br;
  wire        _slots_9_io_out_uop_is_jalr;
  wire        _slots_9_io_out_uop_is_jal;
  wire        _slots_9_io_out_uop_is_sfb;
  wire [19:0] _slots_9_io_out_uop_br_mask;
  wire [4:0]  _slots_9_io_out_uop_br_tag;
  wire [5:0]  _slots_9_io_out_uop_ftq_idx;
  wire        _slots_9_io_out_uop_edge_inst;
  wire [5:0]  _slots_9_io_out_uop_pc_lob;
  wire        _slots_9_io_out_uop_taken;
  wire [19:0] _slots_9_io_out_uop_imm_packed;
  wire [6:0]  _slots_9_io_out_uop_rob_idx;
  wire [4:0]  _slots_9_io_out_uop_ldq_idx;
  wire [4:0]  _slots_9_io_out_uop_stq_idx;
  wire [6:0]  _slots_9_io_out_uop_pdst;
  wire [6:0]  _slots_9_io_out_uop_prs1;
  wire [6:0]  _slots_9_io_out_uop_prs2;
  wire [6:0]  _slots_9_io_out_uop_prs3;
  wire        _slots_9_io_out_uop_prs1_busy;
  wire        _slots_9_io_out_uop_prs2_busy;
  wire        _slots_9_io_out_uop_prs3_busy;
  wire        _slots_9_io_out_uop_ppred_busy;
  wire        _slots_9_io_out_uop_bypassable;
  wire [4:0]  _slots_9_io_out_uop_mem_cmd;
  wire [1:0]  _slots_9_io_out_uop_mem_size;
  wire        _slots_9_io_out_uop_mem_signed;
  wire        _slots_9_io_out_uop_is_fence;
  wire        _slots_9_io_out_uop_is_amo;
  wire        _slots_9_io_out_uop_uses_ldq;
  wire        _slots_9_io_out_uop_uses_stq;
  wire        _slots_9_io_out_uop_ldst_val;
  wire [1:0]  _slots_9_io_out_uop_dst_rtype;
  wire [1:0]  _slots_9_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_9_io_out_uop_lrs2_rtype;
  wire        _slots_9_io_out_uop_fp_val;
  wire [6:0]  _slots_9_io_uop_uopc;
  wire        _slots_9_io_uop_is_rvc;
  wire [9:0]  _slots_9_io_uop_fu_code;
  wire        _slots_9_io_uop_iw_p1_poisoned;
  wire        _slots_9_io_uop_iw_p2_poisoned;
  wire        _slots_9_io_uop_is_br;
  wire        _slots_9_io_uop_is_jalr;
  wire        _slots_9_io_uop_is_jal;
  wire        _slots_9_io_uop_is_sfb;
  wire [19:0] _slots_9_io_uop_br_mask;
  wire [4:0]  _slots_9_io_uop_br_tag;
  wire [5:0]  _slots_9_io_uop_ftq_idx;
  wire        _slots_9_io_uop_edge_inst;
  wire [5:0]  _slots_9_io_uop_pc_lob;
  wire        _slots_9_io_uop_taken;
  wire [19:0] _slots_9_io_uop_imm_packed;
  wire [6:0]  _slots_9_io_uop_rob_idx;
  wire [4:0]  _slots_9_io_uop_ldq_idx;
  wire [4:0]  _slots_9_io_uop_stq_idx;
  wire [6:0]  _slots_9_io_uop_pdst;
  wire [6:0]  _slots_9_io_uop_prs1;
  wire [6:0]  _slots_9_io_uop_prs2;
  wire        _slots_9_io_uop_bypassable;
  wire [4:0]  _slots_9_io_uop_mem_cmd;
  wire        _slots_9_io_uop_is_amo;
  wire        _slots_9_io_uop_uses_stq;
  wire        _slots_9_io_uop_ldst_val;
  wire [1:0]  _slots_9_io_uop_dst_rtype;
  wire [1:0]  _slots_9_io_uop_lrs1_rtype;
  wire [1:0]  _slots_9_io_uop_lrs2_rtype;
  wire        _slots_9_io_uop_fp_val;
  wire        _slots_8_io_valid;
  wire        _slots_8_io_will_be_valid;
  wire        _slots_8_io_request;
  wire [6:0]  _slots_8_io_out_uop_uopc;
  wire        _slots_8_io_out_uop_is_rvc;
  wire [9:0]  _slots_8_io_out_uop_fu_code;
  wire [1:0]  _slots_8_io_out_uop_iw_state;
  wire        _slots_8_io_out_uop_iw_p1_poisoned;
  wire        _slots_8_io_out_uop_iw_p2_poisoned;
  wire        _slots_8_io_out_uop_is_br;
  wire        _slots_8_io_out_uop_is_jalr;
  wire        _slots_8_io_out_uop_is_jal;
  wire        _slots_8_io_out_uop_is_sfb;
  wire [19:0] _slots_8_io_out_uop_br_mask;
  wire [4:0]  _slots_8_io_out_uop_br_tag;
  wire [5:0]  _slots_8_io_out_uop_ftq_idx;
  wire        _slots_8_io_out_uop_edge_inst;
  wire [5:0]  _slots_8_io_out_uop_pc_lob;
  wire        _slots_8_io_out_uop_taken;
  wire [19:0] _slots_8_io_out_uop_imm_packed;
  wire [6:0]  _slots_8_io_out_uop_rob_idx;
  wire [4:0]  _slots_8_io_out_uop_ldq_idx;
  wire [4:0]  _slots_8_io_out_uop_stq_idx;
  wire [6:0]  _slots_8_io_out_uop_pdst;
  wire [6:0]  _slots_8_io_out_uop_prs1;
  wire [6:0]  _slots_8_io_out_uop_prs2;
  wire [6:0]  _slots_8_io_out_uop_prs3;
  wire        _slots_8_io_out_uop_prs1_busy;
  wire        _slots_8_io_out_uop_prs2_busy;
  wire        _slots_8_io_out_uop_prs3_busy;
  wire        _slots_8_io_out_uop_ppred_busy;
  wire        _slots_8_io_out_uop_bypassable;
  wire [4:0]  _slots_8_io_out_uop_mem_cmd;
  wire [1:0]  _slots_8_io_out_uop_mem_size;
  wire        _slots_8_io_out_uop_mem_signed;
  wire        _slots_8_io_out_uop_is_fence;
  wire        _slots_8_io_out_uop_is_amo;
  wire        _slots_8_io_out_uop_uses_ldq;
  wire        _slots_8_io_out_uop_uses_stq;
  wire        _slots_8_io_out_uop_ldst_val;
  wire [1:0]  _slots_8_io_out_uop_dst_rtype;
  wire [1:0]  _slots_8_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_8_io_out_uop_lrs2_rtype;
  wire        _slots_8_io_out_uop_fp_val;
  wire [6:0]  _slots_8_io_uop_uopc;
  wire        _slots_8_io_uop_is_rvc;
  wire [9:0]  _slots_8_io_uop_fu_code;
  wire        _slots_8_io_uop_iw_p1_poisoned;
  wire        _slots_8_io_uop_iw_p2_poisoned;
  wire        _slots_8_io_uop_is_br;
  wire        _slots_8_io_uop_is_jalr;
  wire        _slots_8_io_uop_is_jal;
  wire        _slots_8_io_uop_is_sfb;
  wire [19:0] _slots_8_io_uop_br_mask;
  wire [4:0]  _slots_8_io_uop_br_tag;
  wire [5:0]  _slots_8_io_uop_ftq_idx;
  wire        _slots_8_io_uop_edge_inst;
  wire [5:0]  _slots_8_io_uop_pc_lob;
  wire        _slots_8_io_uop_taken;
  wire [19:0] _slots_8_io_uop_imm_packed;
  wire [6:0]  _slots_8_io_uop_rob_idx;
  wire [4:0]  _slots_8_io_uop_ldq_idx;
  wire [4:0]  _slots_8_io_uop_stq_idx;
  wire [6:0]  _slots_8_io_uop_pdst;
  wire [6:0]  _slots_8_io_uop_prs1;
  wire [6:0]  _slots_8_io_uop_prs2;
  wire        _slots_8_io_uop_bypassable;
  wire [4:0]  _slots_8_io_uop_mem_cmd;
  wire        _slots_8_io_uop_is_amo;
  wire        _slots_8_io_uop_uses_stq;
  wire        _slots_8_io_uop_ldst_val;
  wire [1:0]  _slots_8_io_uop_dst_rtype;
  wire [1:0]  _slots_8_io_uop_lrs1_rtype;
  wire [1:0]  _slots_8_io_uop_lrs2_rtype;
  wire        _slots_8_io_uop_fp_val;
  wire        _slots_7_io_valid;
  wire        _slots_7_io_will_be_valid;
  wire        _slots_7_io_request;
  wire [6:0]  _slots_7_io_out_uop_uopc;
  wire        _slots_7_io_out_uop_is_rvc;
  wire [9:0]  _slots_7_io_out_uop_fu_code;
  wire [1:0]  _slots_7_io_out_uop_iw_state;
  wire        _slots_7_io_out_uop_iw_p1_poisoned;
  wire        _slots_7_io_out_uop_iw_p2_poisoned;
  wire        _slots_7_io_out_uop_is_br;
  wire        _slots_7_io_out_uop_is_jalr;
  wire        _slots_7_io_out_uop_is_jal;
  wire        _slots_7_io_out_uop_is_sfb;
  wire [19:0] _slots_7_io_out_uop_br_mask;
  wire [4:0]  _slots_7_io_out_uop_br_tag;
  wire [5:0]  _slots_7_io_out_uop_ftq_idx;
  wire        _slots_7_io_out_uop_edge_inst;
  wire [5:0]  _slots_7_io_out_uop_pc_lob;
  wire        _slots_7_io_out_uop_taken;
  wire [19:0] _slots_7_io_out_uop_imm_packed;
  wire [6:0]  _slots_7_io_out_uop_rob_idx;
  wire [4:0]  _slots_7_io_out_uop_ldq_idx;
  wire [4:0]  _slots_7_io_out_uop_stq_idx;
  wire [6:0]  _slots_7_io_out_uop_pdst;
  wire [6:0]  _slots_7_io_out_uop_prs1;
  wire [6:0]  _slots_7_io_out_uop_prs2;
  wire [6:0]  _slots_7_io_out_uop_prs3;
  wire        _slots_7_io_out_uop_prs1_busy;
  wire        _slots_7_io_out_uop_prs2_busy;
  wire        _slots_7_io_out_uop_prs3_busy;
  wire        _slots_7_io_out_uop_ppred_busy;
  wire        _slots_7_io_out_uop_bypassable;
  wire [4:0]  _slots_7_io_out_uop_mem_cmd;
  wire [1:0]  _slots_7_io_out_uop_mem_size;
  wire        _slots_7_io_out_uop_mem_signed;
  wire        _slots_7_io_out_uop_is_fence;
  wire        _slots_7_io_out_uop_is_amo;
  wire        _slots_7_io_out_uop_uses_ldq;
  wire        _slots_7_io_out_uop_uses_stq;
  wire        _slots_7_io_out_uop_ldst_val;
  wire [1:0]  _slots_7_io_out_uop_dst_rtype;
  wire [1:0]  _slots_7_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_7_io_out_uop_lrs2_rtype;
  wire        _slots_7_io_out_uop_fp_val;
  wire [6:0]  _slots_7_io_uop_uopc;
  wire        _slots_7_io_uop_is_rvc;
  wire [9:0]  _slots_7_io_uop_fu_code;
  wire        _slots_7_io_uop_iw_p1_poisoned;
  wire        _slots_7_io_uop_iw_p2_poisoned;
  wire        _slots_7_io_uop_is_br;
  wire        _slots_7_io_uop_is_jalr;
  wire        _slots_7_io_uop_is_jal;
  wire        _slots_7_io_uop_is_sfb;
  wire [19:0] _slots_7_io_uop_br_mask;
  wire [4:0]  _slots_7_io_uop_br_tag;
  wire [5:0]  _slots_7_io_uop_ftq_idx;
  wire        _slots_7_io_uop_edge_inst;
  wire [5:0]  _slots_7_io_uop_pc_lob;
  wire        _slots_7_io_uop_taken;
  wire [19:0] _slots_7_io_uop_imm_packed;
  wire [6:0]  _slots_7_io_uop_rob_idx;
  wire [4:0]  _slots_7_io_uop_ldq_idx;
  wire [4:0]  _slots_7_io_uop_stq_idx;
  wire [6:0]  _slots_7_io_uop_pdst;
  wire [6:0]  _slots_7_io_uop_prs1;
  wire [6:0]  _slots_7_io_uop_prs2;
  wire        _slots_7_io_uop_bypassable;
  wire [4:0]  _slots_7_io_uop_mem_cmd;
  wire        _slots_7_io_uop_is_amo;
  wire        _slots_7_io_uop_uses_stq;
  wire        _slots_7_io_uop_ldst_val;
  wire [1:0]  _slots_7_io_uop_dst_rtype;
  wire [1:0]  _slots_7_io_uop_lrs1_rtype;
  wire [1:0]  _slots_7_io_uop_lrs2_rtype;
  wire        _slots_7_io_uop_fp_val;
  wire        _slots_6_io_valid;
  wire        _slots_6_io_will_be_valid;
  wire        _slots_6_io_request;
  wire [6:0]  _slots_6_io_out_uop_uopc;
  wire        _slots_6_io_out_uop_is_rvc;
  wire [9:0]  _slots_6_io_out_uop_fu_code;
  wire [1:0]  _slots_6_io_out_uop_iw_state;
  wire        _slots_6_io_out_uop_iw_p1_poisoned;
  wire        _slots_6_io_out_uop_iw_p2_poisoned;
  wire        _slots_6_io_out_uop_is_br;
  wire        _slots_6_io_out_uop_is_jalr;
  wire        _slots_6_io_out_uop_is_jal;
  wire        _slots_6_io_out_uop_is_sfb;
  wire [19:0] _slots_6_io_out_uop_br_mask;
  wire [4:0]  _slots_6_io_out_uop_br_tag;
  wire [5:0]  _slots_6_io_out_uop_ftq_idx;
  wire        _slots_6_io_out_uop_edge_inst;
  wire [5:0]  _slots_6_io_out_uop_pc_lob;
  wire        _slots_6_io_out_uop_taken;
  wire [19:0] _slots_6_io_out_uop_imm_packed;
  wire [6:0]  _slots_6_io_out_uop_rob_idx;
  wire [4:0]  _slots_6_io_out_uop_ldq_idx;
  wire [4:0]  _slots_6_io_out_uop_stq_idx;
  wire [6:0]  _slots_6_io_out_uop_pdst;
  wire [6:0]  _slots_6_io_out_uop_prs1;
  wire [6:0]  _slots_6_io_out_uop_prs2;
  wire [6:0]  _slots_6_io_out_uop_prs3;
  wire        _slots_6_io_out_uop_prs1_busy;
  wire        _slots_6_io_out_uop_prs2_busy;
  wire        _slots_6_io_out_uop_prs3_busy;
  wire        _slots_6_io_out_uop_ppred_busy;
  wire        _slots_6_io_out_uop_bypassable;
  wire [4:0]  _slots_6_io_out_uop_mem_cmd;
  wire [1:0]  _slots_6_io_out_uop_mem_size;
  wire        _slots_6_io_out_uop_mem_signed;
  wire        _slots_6_io_out_uop_is_fence;
  wire        _slots_6_io_out_uop_is_amo;
  wire        _slots_6_io_out_uop_uses_ldq;
  wire        _slots_6_io_out_uop_uses_stq;
  wire        _slots_6_io_out_uop_ldst_val;
  wire [1:0]  _slots_6_io_out_uop_dst_rtype;
  wire [1:0]  _slots_6_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_6_io_out_uop_lrs2_rtype;
  wire        _slots_6_io_out_uop_fp_val;
  wire [6:0]  _slots_6_io_uop_uopc;
  wire        _slots_6_io_uop_is_rvc;
  wire [9:0]  _slots_6_io_uop_fu_code;
  wire        _slots_6_io_uop_iw_p1_poisoned;
  wire        _slots_6_io_uop_iw_p2_poisoned;
  wire        _slots_6_io_uop_is_br;
  wire        _slots_6_io_uop_is_jalr;
  wire        _slots_6_io_uop_is_jal;
  wire        _slots_6_io_uop_is_sfb;
  wire [19:0] _slots_6_io_uop_br_mask;
  wire [4:0]  _slots_6_io_uop_br_tag;
  wire [5:0]  _slots_6_io_uop_ftq_idx;
  wire        _slots_6_io_uop_edge_inst;
  wire [5:0]  _slots_6_io_uop_pc_lob;
  wire        _slots_6_io_uop_taken;
  wire [19:0] _slots_6_io_uop_imm_packed;
  wire [6:0]  _slots_6_io_uop_rob_idx;
  wire [4:0]  _slots_6_io_uop_ldq_idx;
  wire [4:0]  _slots_6_io_uop_stq_idx;
  wire [6:0]  _slots_6_io_uop_pdst;
  wire [6:0]  _slots_6_io_uop_prs1;
  wire [6:0]  _slots_6_io_uop_prs2;
  wire        _slots_6_io_uop_bypassable;
  wire [4:0]  _slots_6_io_uop_mem_cmd;
  wire        _slots_6_io_uop_is_amo;
  wire        _slots_6_io_uop_uses_stq;
  wire        _slots_6_io_uop_ldst_val;
  wire [1:0]  _slots_6_io_uop_dst_rtype;
  wire [1:0]  _slots_6_io_uop_lrs1_rtype;
  wire [1:0]  _slots_6_io_uop_lrs2_rtype;
  wire        _slots_6_io_uop_fp_val;
  wire        _slots_5_io_valid;
  wire        _slots_5_io_will_be_valid;
  wire        _slots_5_io_request;
  wire [6:0]  _slots_5_io_out_uop_uopc;
  wire        _slots_5_io_out_uop_is_rvc;
  wire [9:0]  _slots_5_io_out_uop_fu_code;
  wire [1:0]  _slots_5_io_out_uop_iw_state;
  wire        _slots_5_io_out_uop_iw_p1_poisoned;
  wire        _slots_5_io_out_uop_iw_p2_poisoned;
  wire        _slots_5_io_out_uop_is_br;
  wire        _slots_5_io_out_uop_is_jalr;
  wire        _slots_5_io_out_uop_is_jal;
  wire        _slots_5_io_out_uop_is_sfb;
  wire [19:0] _slots_5_io_out_uop_br_mask;
  wire [4:0]  _slots_5_io_out_uop_br_tag;
  wire [5:0]  _slots_5_io_out_uop_ftq_idx;
  wire        _slots_5_io_out_uop_edge_inst;
  wire [5:0]  _slots_5_io_out_uop_pc_lob;
  wire        _slots_5_io_out_uop_taken;
  wire [19:0] _slots_5_io_out_uop_imm_packed;
  wire [6:0]  _slots_5_io_out_uop_rob_idx;
  wire [4:0]  _slots_5_io_out_uop_ldq_idx;
  wire [4:0]  _slots_5_io_out_uop_stq_idx;
  wire [6:0]  _slots_5_io_out_uop_pdst;
  wire [6:0]  _slots_5_io_out_uop_prs1;
  wire [6:0]  _slots_5_io_out_uop_prs2;
  wire [6:0]  _slots_5_io_out_uop_prs3;
  wire        _slots_5_io_out_uop_prs1_busy;
  wire        _slots_5_io_out_uop_prs2_busy;
  wire        _slots_5_io_out_uop_prs3_busy;
  wire        _slots_5_io_out_uop_ppred_busy;
  wire        _slots_5_io_out_uop_bypassable;
  wire [4:0]  _slots_5_io_out_uop_mem_cmd;
  wire [1:0]  _slots_5_io_out_uop_mem_size;
  wire        _slots_5_io_out_uop_mem_signed;
  wire        _slots_5_io_out_uop_is_fence;
  wire        _slots_5_io_out_uop_is_amo;
  wire        _slots_5_io_out_uop_uses_ldq;
  wire        _slots_5_io_out_uop_uses_stq;
  wire        _slots_5_io_out_uop_ldst_val;
  wire [1:0]  _slots_5_io_out_uop_dst_rtype;
  wire [1:0]  _slots_5_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_5_io_out_uop_lrs2_rtype;
  wire        _slots_5_io_out_uop_fp_val;
  wire [6:0]  _slots_5_io_uop_uopc;
  wire        _slots_5_io_uop_is_rvc;
  wire [9:0]  _slots_5_io_uop_fu_code;
  wire        _slots_5_io_uop_iw_p1_poisoned;
  wire        _slots_5_io_uop_iw_p2_poisoned;
  wire        _slots_5_io_uop_is_br;
  wire        _slots_5_io_uop_is_jalr;
  wire        _slots_5_io_uop_is_jal;
  wire        _slots_5_io_uop_is_sfb;
  wire [19:0] _slots_5_io_uop_br_mask;
  wire [4:0]  _slots_5_io_uop_br_tag;
  wire [5:0]  _slots_5_io_uop_ftq_idx;
  wire        _slots_5_io_uop_edge_inst;
  wire [5:0]  _slots_5_io_uop_pc_lob;
  wire        _slots_5_io_uop_taken;
  wire [19:0] _slots_5_io_uop_imm_packed;
  wire [6:0]  _slots_5_io_uop_rob_idx;
  wire [4:0]  _slots_5_io_uop_ldq_idx;
  wire [4:0]  _slots_5_io_uop_stq_idx;
  wire [6:0]  _slots_5_io_uop_pdst;
  wire [6:0]  _slots_5_io_uop_prs1;
  wire [6:0]  _slots_5_io_uop_prs2;
  wire        _slots_5_io_uop_bypassable;
  wire [4:0]  _slots_5_io_uop_mem_cmd;
  wire        _slots_5_io_uop_is_amo;
  wire        _slots_5_io_uop_uses_stq;
  wire        _slots_5_io_uop_ldst_val;
  wire [1:0]  _slots_5_io_uop_dst_rtype;
  wire [1:0]  _slots_5_io_uop_lrs1_rtype;
  wire [1:0]  _slots_5_io_uop_lrs2_rtype;
  wire        _slots_5_io_uop_fp_val;
  wire        _slots_4_io_valid;
  wire        _slots_4_io_will_be_valid;
  wire        _slots_4_io_request;
  wire [6:0]  _slots_4_io_out_uop_uopc;
  wire        _slots_4_io_out_uop_is_rvc;
  wire [9:0]  _slots_4_io_out_uop_fu_code;
  wire [1:0]  _slots_4_io_out_uop_iw_state;
  wire        _slots_4_io_out_uop_iw_p1_poisoned;
  wire        _slots_4_io_out_uop_iw_p2_poisoned;
  wire        _slots_4_io_out_uop_is_br;
  wire        _slots_4_io_out_uop_is_jalr;
  wire        _slots_4_io_out_uop_is_jal;
  wire        _slots_4_io_out_uop_is_sfb;
  wire [19:0] _slots_4_io_out_uop_br_mask;
  wire [4:0]  _slots_4_io_out_uop_br_tag;
  wire [5:0]  _slots_4_io_out_uop_ftq_idx;
  wire        _slots_4_io_out_uop_edge_inst;
  wire [5:0]  _slots_4_io_out_uop_pc_lob;
  wire        _slots_4_io_out_uop_taken;
  wire [19:0] _slots_4_io_out_uop_imm_packed;
  wire [6:0]  _slots_4_io_out_uop_rob_idx;
  wire [4:0]  _slots_4_io_out_uop_ldq_idx;
  wire [4:0]  _slots_4_io_out_uop_stq_idx;
  wire [6:0]  _slots_4_io_out_uop_pdst;
  wire [6:0]  _slots_4_io_out_uop_prs1;
  wire [6:0]  _slots_4_io_out_uop_prs2;
  wire [6:0]  _slots_4_io_out_uop_prs3;
  wire        _slots_4_io_out_uop_prs1_busy;
  wire        _slots_4_io_out_uop_prs2_busy;
  wire        _slots_4_io_out_uop_prs3_busy;
  wire        _slots_4_io_out_uop_ppred_busy;
  wire        _slots_4_io_out_uop_bypassable;
  wire [4:0]  _slots_4_io_out_uop_mem_cmd;
  wire [1:0]  _slots_4_io_out_uop_mem_size;
  wire        _slots_4_io_out_uop_mem_signed;
  wire        _slots_4_io_out_uop_is_fence;
  wire        _slots_4_io_out_uop_is_amo;
  wire        _slots_4_io_out_uop_uses_ldq;
  wire        _slots_4_io_out_uop_uses_stq;
  wire        _slots_4_io_out_uop_ldst_val;
  wire [1:0]  _slots_4_io_out_uop_dst_rtype;
  wire [1:0]  _slots_4_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_4_io_out_uop_lrs2_rtype;
  wire        _slots_4_io_out_uop_fp_val;
  wire [6:0]  _slots_4_io_uop_uopc;
  wire        _slots_4_io_uop_is_rvc;
  wire [9:0]  _slots_4_io_uop_fu_code;
  wire        _slots_4_io_uop_iw_p1_poisoned;
  wire        _slots_4_io_uop_iw_p2_poisoned;
  wire        _slots_4_io_uop_is_br;
  wire        _slots_4_io_uop_is_jalr;
  wire        _slots_4_io_uop_is_jal;
  wire        _slots_4_io_uop_is_sfb;
  wire [19:0] _slots_4_io_uop_br_mask;
  wire [4:0]  _slots_4_io_uop_br_tag;
  wire [5:0]  _slots_4_io_uop_ftq_idx;
  wire        _slots_4_io_uop_edge_inst;
  wire [5:0]  _slots_4_io_uop_pc_lob;
  wire        _slots_4_io_uop_taken;
  wire [19:0] _slots_4_io_uop_imm_packed;
  wire [6:0]  _slots_4_io_uop_rob_idx;
  wire [4:0]  _slots_4_io_uop_ldq_idx;
  wire [4:0]  _slots_4_io_uop_stq_idx;
  wire [6:0]  _slots_4_io_uop_pdst;
  wire [6:0]  _slots_4_io_uop_prs1;
  wire [6:0]  _slots_4_io_uop_prs2;
  wire        _slots_4_io_uop_bypassable;
  wire [4:0]  _slots_4_io_uop_mem_cmd;
  wire        _slots_4_io_uop_is_amo;
  wire        _slots_4_io_uop_uses_stq;
  wire        _slots_4_io_uop_ldst_val;
  wire [1:0]  _slots_4_io_uop_dst_rtype;
  wire [1:0]  _slots_4_io_uop_lrs1_rtype;
  wire [1:0]  _slots_4_io_uop_lrs2_rtype;
  wire        _slots_4_io_uop_fp_val;
  wire        _slots_3_io_valid;
  wire        _slots_3_io_will_be_valid;
  wire        _slots_3_io_request;
  wire [6:0]  _slots_3_io_out_uop_uopc;
  wire        _slots_3_io_out_uop_is_rvc;
  wire [9:0]  _slots_3_io_out_uop_fu_code;
  wire [1:0]  _slots_3_io_out_uop_iw_state;
  wire        _slots_3_io_out_uop_iw_p1_poisoned;
  wire        _slots_3_io_out_uop_iw_p2_poisoned;
  wire        _slots_3_io_out_uop_is_br;
  wire        _slots_3_io_out_uop_is_jalr;
  wire        _slots_3_io_out_uop_is_jal;
  wire        _slots_3_io_out_uop_is_sfb;
  wire [19:0] _slots_3_io_out_uop_br_mask;
  wire [4:0]  _slots_3_io_out_uop_br_tag;
  wire [5:0]  _slots_3_io_out_uop_ftq_idx;
  wire        _slots_3_io_out_uop_edge_inst;
  wire [5:0]  _slots_3_io_out_uop_pc_lob;
  wire        _slots_3_io_out_uop_taken;
  wire [19:0] _slots_3_io_out_uop_imm_packed;
  wire [6:0]  _slots_3_io_out_uop_rob_idx;
  wire [4:0]  _slots_3_io_out_uop_ldq_idx;
  wire [4:0]  _slots_3_io_out_uop_stq_idx;
  wire [6:0]  _slots_3_io_out_uop_pdst;
  wire [6:0]  _slots_3_io_out_uop_prs1;
  wire [6:0]  _slots_3_io_out_uop_prs2;
  wire [6:0]  _slots_3_io_out_uop_prs3;
  wire        _slots_3_io_out_uop_prs1_busy;
  wire        _slots_3_io_out_uop_prs2_busy;
  wire        _slots_3_io_out_uop_prs3_busy;
  wire        _slots_3_io_out_uop_ppred_busy;
  wire        _slots_3_io_out_uop_bypassable;
  wire [4:0]  _slots_3_io_out_uop_mem_cmd;
  wire [1:0]  _slots_3_io_out_uop_mem_size;
  wire        _slots_3_io_out_uop_mem_signed;
  wire        _slots_3_io_out_uop_is_fence;
  wire        _slots_3_io_out_uop_is_amo;
  wire        _slots_3_io_out_uop_uses_ldq;
  wire        _slots_3_io_out_uop_uses_stq;
  wire        _slots_3_io_out_uop_ldst_val;
  wire [1:0]  _slots_3_io_out_uop_dst_rtype;
  wire [1:0]  _slots_3_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_3_io_out_uop_lrs2_rtype;
  wire        _slots_3_io_out_uop_fp_val;
  wire [6:0]  _slots_3_io_uop_uopc;
  wire        _slots_3_io_uop_is_rvc;
  wire [9:0]  _slots_3_io_uop_fu_code;
  wire        _slots_3_io_uop_iw_p1_poisoned;
  wire        _slots_3_io_uop_iw_p2_poisoned;
  wire        _slots_3_io_uop_is_br;
  wire        _slots_3_io_uop_is_jalr;
  wire        _slots_3_io_uop_is_jal;
  wire        _slots_3_io_uop_is_sfb;
  wire [19:0] _slots_3_io_uop_br_mask;
  wire [4:0]  _slots_3_io_uop_br_tag;
  wire [5:0]  _slots_3_io_uop_ftq_idx;
  wire        _slots_3_io_uop_edge_inst;
  wire [5:0]  _slots_3_io_uop_pc_lob;
  wire        _slots_3_io_uop_taken;
  wire [19:0] _slots_3_io_uop_imm_packed;
  wire [6:0]  _slots_3_io_uop_rob_idx;
  wire [4:0]  _slots_3_io_uop_ldq_idx;
  wire [4:0]  _slots_3_io_uop_stq_idx;
  wire [6:0]  _slots_3_io_uop_pdst;
  wire [6:0]  _slots_3_io_uop_prs1;
  wire [6:0]  _slots_3_io_uop_prs2;
  wire        _slots_3_io_uop_bypassable;
  wire [4:0]  _slots_3_io_uop_mem_cmd;
  wire        _slots_3_io_uop_is_amo;
  wire        _slots_3_io_uop_uses_stq;
  wire        _slots_3_io_uop_ldst_val;
  wire [1:0]  _slots_3_io_uop_dst_rtype;
  wire [1:0]  _slots_3_io_uop_lrs1_rtype;
  wire [1:0]  _slots_3_io_uop_lrs2_rtype;
  wire        _slots_3_io_uop_fp_val;
  wire        _slots_2_io_valid;
  wire        _slots_2_io_will_be_valid;
  wire        _slots_2_io_request;
  wire [6:0]  _slots_2_io_out_uop_uopc;
  wire        _slots_2_io_out_uop_is_rvc;
  wire [9:0]  _slots_2_io_out_uop_fu_code;
  wire [1:0]  _slots_2_io_out_uop_iw_state;
  wire        _slots_2_io_out_uop_iw_p1_poisoned;
  wire        _slots_2_io_out_uop_iw_p2_poisoned;
  wire        _slots_2_io_out_uop_is_br;
  wire        _slots_2_io_out_uop_is_jalr;
  wire        _slots_2_io_out_uop_is_jal;
  wire        _slots_2_io_out_uop_is_sfb;
  wire [19:0] _slots_2_io_out_uop_br_mask;
  wire [4:0]  _slots_2_io_out_uop_br_tag;
  wire [5:0]  _slots_2_io_out_uop_ftq_idx;
  wire        _slots_2_io_out_uop_edge_inst;
  wire [5:0]  _slots_2_io_out_uop_pc_lob;
  wire        _slots_2_io_out_uop_taken;
  wire [19:0] _slots_2_io_out_uop_imm_packed;
  wire [6:0]  _slots_2_io_out_uop_rob_idx;
  wire [4:0]  _slots_2_io_out_uop_ldq_idx;
  wire [4:0]  _slots_2_io_out_uop_stq_idx;
  wire [6:0]  _slots_2_io_out_uop_pdst;
  wire [6:0]  _slots_2_io_out_uop_prs1;
  wire [6:0]  _slots_2_io_out_uop_prs2;
  wire [6:0]  _slots_2_io_out_uop_prs3;
  wire        _slots_2_io_out_uop_prs1_busy;
  wire        _slots_2_io_out_uop_prs2_busy;
  wire        _slots_2_io_out_uop_prs3_busy;
  wire        _slots_2_io_out_uop_ppred_busy;
  wire        _slots_2_io_out_uop_bypassable;
  wire [4:0]  _slots_2_io_out_uop_mem_cmd;
  wire [1:0]  _slots_2_io_out_uop_mem_size;
  wire        _slots_2_io_out_uop_mem_signed;
  wire        _slots_2_io_out_uop_is_fence;
  wire        _slots_2_io_out_uop_is_amo;
  wire        _slots_2_io_out_uop_uses_ldq;
  wire        _slots_2_io_out_uop_uses_stq;
  wire        _slots_2_io_out_uop_ldst_val;
  wire [1:0]  _slots_2_io_out_uop_dst_rtype;
  wire [1:0]  _slots_2_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_2_io_out_uop_lrs2_rtype;
  wire        _slots_2_io_out_uop_fp_val;
  wire [6:0]  _slots_2_io_uop_uopc;
  wire        _slots_2_io_uop_is_rvc;
  wire [9:0]  _slots_2_io_uop_fu_code;
  wire        _slots_2_io_uop_iw_p1_poisoned;
  wire        _slots_2_io_uop_iw_p2_poisoned;
  wire        _slots_2_io_uop_is_br;
  wire        _slots_2_io_uop_is_jalr;
  wire        _slots_2_io_uop_is_jal;
  wire        _slots_2_io_uop_is_sfb;
  wire [19:0] _slots_2_io_uop_br_mask;
  wire [4:0]  _slots_2_io_uop_br_tag;
  wire [5:0]  _slots_2_io_uop_ftq_idx;
  wire        _slots_2_io_uop_edge_inst;
  wire [5:0]  _slots_2_io_uop_pc_lob;
  wire        _slots_2_io_uop_taken;
  wire [19:0] _slots_2_io_uop_imm_packed;
  wire [6:0]  _slots_2_io_uop_rob_idx;
  wire [4:0]  _slots_2_io_uop_ldq_idx;
  wire [4:0]  _slots_2_io_uop_stq_idx;
  wire [6:0]  _slots_2_io_uop_pdst;
  wire [6:0]  _slots_2_io_uop_prs1;
  wire [6:0]  _slots_2_io_uop_prs2;
  wire        _slots_2_io_uop_bypassable;
  wire [4:0]  _slots_2_io_uop_mem_cmd;
  wire        _slots_2_io_uop_is_amo;
  wire        _slots_2_io_uop_uses_stq;
  wire        _slots_2_io_uop_ldst_val;
  wire [1:0]  _slots_2_io_uop_dst_rtype;
  wire [1:0]  _slots_2_io_uop_lrs1_rtype;
  wire [1:0]  _slots_2_io_uop_lrs2_rtype;
  wire        _slots_2_io_uop_fp_val;
  wire        _slots_1_io_valid;
  wire        _slots_1_io_will_be_valid;
  wire        _slots_1_io_request;
  wire [6:0]  _slots_1_io_out_uop_uopc;
  wire        _slots_1_io_out_uop_is_rvc;
  wire [9:0]  _slots_1_io_out_uop_fu_code;
  wire [1:0]  _slots_1_io_out_uop_iw_state;
  wire        _slots_1_io_out_uop_iw_p1_poisoned;
  wire        _slots_1_io_out_uop_iw_p2_poisoned;
  wire        _slots_1_io_out_uop_is_br;
  wire        _slots_1_io_out_uop_is_jalr;
  wire        _slots_1_io_out_uop_is_jal;
  wire        _slots_1_io_out_uop_is_sfb;
  wire [19:0] _slots_1_io_out_uop_br_mask;
  wire [4:0]  _slots_1_io_out_uop_br_tag;
  wire [5:0]  _slots_1_io_out_uop_ftq_idx;
  wire        _slots_1_io_out_uop_edge_inst;
  wire [5:0]  _slots_1_io_out_uop_pc_lob;
  wire        _slots_1_io_out_uop_taken;
  wire [19:0] _slots_1_io_out_uop_imm_packed;
  wire [6:0]  _slots_1_io_out_uop_rob_idx;
  wire [4:0]  _slots_1_io_out_uop_ldq_idx;
  wire [4:0]  _slots_1_io_out_uop_stq_idx;
  wire [6:0]  _slots_1_io_out_uop_pdst;
  wire [6:0]  _slots_1_io_out_uop_prs1;
  wire [6:0]  _slots_1_io_out_uop_prs2;
  wire [6:0]  _slots_1_io_out_uop_prs3;
  wire        _slots_1_io_out_uop_prs1_busy;
  wire        _slots_1_io_out_uop_prs2_busy;
  wire        _slots_1_io_out_uop_prs3_busy;
  wire        _slots_1_io_out_uop_ppred_busy;
  wire        _slots_1_io_out_uop_bypassable;
  wire [4:0]  _slots_1_io_out_uop_mem_cmd;
  wire [1:0]  _slots_1_io_out_uop_mem_size;
  wire        _slots_1_io_out_uop_mem_signed;
  wire        _slots_1_io_out_uop_is_fence;
  wire        _slots_1_io_out_uop_is_amo;
  wire        _slots_1_io_out_uop_uses_ldq;
  wire        _slots_1_io_out_uop_uses_stq;
  wire        _slots_1_io_out_uop_ldst_val;
  wire [1:0]  _slots_1_io_out_uop_dst_rtype;
  wire [1:0]  _slots_1_io_out_uop_lrs1_rtype;
  wire [1:0]  _slots_1_io_out_uop_lrs2_rtype;
  wire        _slots_1_io_out_uop_fp_val;
  wire [6:0]  _slots_1_io_uop_uopc;
  wire        _slots_1_io_uop_is_rvc;
  wire [9:0]  _slots_1_io_uop_fu_code;
  wire        _slots_1_io_uop_iw_p1_poisoned;
  wire        _slots_1_io_uop_iw_p2_poisoned;
  wire        _slots_1_io_uop_is_br;
  wire        _slots_1_io_uop_is_jalr;
  wire        _slots_1_io_uop_is_jal;
  wire        _slots_1_io_uop_is_sfb;
  wire [19:0] _slots_1_io_uop_br_mask;
  wire [4:0]  _slots_1_io_uop_br_tag;
  wire [5:0]  _slots_1_io_uop_ftq_idx;
  wire        _slots_1_io_uop_edge_inst;
  wire [5:0]  _slots_1_io_uop_pc_lob;
  wire        _slots_1_io_uop_taken;
  wire [19:0] _slots_1_io_uop_imm_packed;
  wire [6:0]  _slots_1_io_uop_rob_idx;
  wire [4:0]  _slots_1_io_uop_ldq_idx;
  wire [4:0]  _slots_1_io_uop_stq_idx;
  wire [6:0]  _slots_1_io_uop_pdst;
  wire [6:0]  _slots_1_io_uop_prs1;
  wire [6:0]  _slots_1_io_uop_prs2;
  wire        _slots_1_io_uop_bypassable;
  wire [4:0]  _slots_1_io_uop_mem_cmd;
  wire        _slots_1_io_uop_is_amo;
  wire        _slots_1_io_uop_uses_stq;
  wire        _slots_1_io_uop_ldst_val;
  wire [1:0]  _slots_1_io_uop_dst_rtype;
  wire [1:0]  _slots_1_io_uop_lrs1_rtype;
  wire [1:0]  _slots_1_io_uop_lrs2_rtype;
  wire        _slots_1_io_uop_fp_val;
  wire        _slots_0_io_valid;
  wire        _slots_0_io_will_be_valid;
  wire        _slots_0_io_request;
  wire [6:0]  _slots_0_io_uop_uopc;
  wire        _slots_0_io_uop_is_rvc;
  wire [9:0]  _slots_0_io_uop_fu_code;
  wire        _slots_0_io_uop_iw_p1_poisoned;
  wire        _slots_0_io_uop_iw_p2_poisoned;
  wire        _slots_0_io_uop_is_br;
  wire        _slots_0_io_uop_is_jalr;
  wire        _slots_0_io_uop_is_jal;
  wire        _slots_0_io_uop_is_sfb;
  wire [19:0] _slots_0_io_uop_br_mask;
  wire [4:0]  _slots_0_io_uop_br_tag;
  wire [5:0]  _slots_0_io_uop_ftq_idx;
  wire        _slots_0_io_uop_edge_inst;
  wire [5:0]  _slots_0_io_uop_pc_lob;
  wire        _slots_0_io_uop_taken;
  wire [19:0] _slots_0_io_uop_imm_packed;
  wire [6:0]  _slots_0_io_uop_rob_idx;
  wire [4:0]  _slots_0_io_uop_ldq_idx;
  wire [4:0]  _slots_0_io_uop_stq_idx;
  wire [6:0]  _slots_0_io_uop_pdst;
  wire [6:0]  _slots_0_io_uop_prs1;
  wire [6:0]  _slots_0_io_uop_prs2;
  wire        _slots_0_io_uop_bypassable;
  wire [4:0]  _slots_0_io_uop_mem_cmd;
  wire        _slots_0_io_uop_is_amo;
  wire        _slots_0_io_uop_uses_stq;
  wire        _slots_0_io_uop_ldst_val;
  wire [1:0]  _slots_0_io_uop_dst_rtype;
  wire [1:0]  _slots_0_io_uop_lrs1_rtype;
  wire [1:0]  _slots_0_io_uop_lrs2_rtype;
  wire        _slots_0_io_uop_fp_val;
  wire        _GEN = io_dis_uops_0_bits_uopc == 7'h2;
  wire        _GEN_0 = _GEN & ~(|io_dis_uops_0_bits_lrs2_rtype) | io_dis_uops_0_bits_uopc == 7'h43;
  wire [1:0]  _GEN_12648 = _GEN_0 ? 2'h2 : 2'h1;
  wire        _GEN_1 = _GEN_0 | ~(_GEN & (|io_dis_uops_0_bits_lrs2_rtype));
  wire [1:0]  _GEN_12597 = _GEN_1 ? io_dis_uops_0_bits_lrs2_rtype : 2'h2;
  wire        _GEN_12623 = _GEN_1 & io_dis_uops_0_bits_prs2_busy;
  wire        _GEN_2 = io_dis_uops_1_bits_uopc == 7'h2;
  wire        _GEN_3 = _GEN_2 & ~(|io_dis_uops_1_bits_lrs2_rtype) | io_dis_uops_1_bits_uopc == 7'h43;
  wire [1:0]  _GEN_7 = _GEN_3 ? 2'h2 : 2'h1;
  wire        _GEN_4 = _GEN_3 | ~(_GEN_2 & (|io_dis_uops_1_bits_lrs2_rtype));
  wire [1:0]  _GEN_8 = _GEN_4 ? io_dis_uops_1_bits_lrs2_rtype : 2'h2;
  wire        _GEN_9 = _GEN_4 & io_dis_uops_1_bits_prs2_busy;
  wire        _GEN_5 = io_dis_uops_2_bits_uopc == 7'h2;
  wire        _GEN_6 = _GEN_5 & ~(|io_dis_uops_2_bits_lrs2_rtype) | io_dis_uops_2_bits_uopc == 7'h43;
  wire        _GEN_10 = _GEN_6 | ~(_GEN_5 & (|io_dis_uops_2_bits_lrs2_rtype));
  wire [1:0]  _GEN_13 = _GEN_10 ? io_dis_uops_2_bits_lrs2_rtype : 2'h2;
  wire        _GEN_14 = _GEN_10 & io_dis_uops_2_bits_prs2_busy;
  wire        _GEN_11 = io_dis_uops_3_bits_uopc == 7'h2;
  wire        _GEN_12 = _GEN_11 & ~(|io_dis_uops_3_bits_lrs2_rtype) | io_dis_uops_3_bits_uopc == 7'h43;
  wire        _GEN_15 = _GEN_12 | ~(_GEN_11 & (|io_dis_uops_3_bits_lrs2_rtype));
  wire [9:0]  _can_allocate_T_2 = _slots_0_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_16 = {_slots_0_io_uop_fu_code[5], _slots_0_io_uop_fu_code[0]};
  wire [9:0]  _can_allocate_T = _slots_0_io_uop_fu_code & io_fu_types_0;
  wire        _GEN_17 = _slots_0_io_request & (|_can_allocate_T);
  wire        _GEN_18 = _slots_0_io_request & (|_GEN_16) | _GEN_17;
  wire        _GEN_19 = _slots_0_io_request & ~(_slots_0_io_request & (|_can_allocate_T_2) | _GEN_18);
  wire [9:0]  _can_allocate_T_3 = _slots_0_io_uop_fu_code & io_fu_types_3;
  wire        _GEN_13149 = _GEN_19 & (|_can_allocate_T_3);
  wire        _GEN_20 = _slots_0_io_request & ~_GEN_18;
  wire        _GEN_13068 = _GEN_20 & (|_can_allocate_T_2);
  wire        _GEN_21 = _slots_0_io_request & ~_GEN_17;
  wire        _GEN_12987 = _GEN_21 & (|_GEN_16);
  wire        _GEN_12906 = _slots_0_io_request & (|_can_allocate_T);
  wire        issue_slots_0_grant = _GEN_13149 | _GEN_13068 | _GEN_12987 | _GEN_12906;
  wire [9:0]  _can_allocate_T_6 = _slots_1_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_22 = _GEN_20 & (|_can_allocate_T_2);
  wire [1:0]  _GEN_23 = {_slots_1_io_uop_fu_code[5], _slots_1_io_uop_fu_code[0]};
  wire        _GEN_24 = _GEN_21 & (|_GEN_16);
  wire        _GEN_26 = _slots_1_io_request & (|(_slots_1_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_28 = _GEN_26 & ~_GEN_17;
  wire        _GEN_30 = _slots_1_io_request & (|_GEN_23) & ~_GEN_24 | _GEN_28;
  wire        _GEN_32 = _slots_1_io_request & ~(_slots_1_io_request & (|_can_allocate_T_6) & ~_GEN_22 | _GEN_30) & (|(_slots_1_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_34 = _GEN_19 & (|_can_allocate_T_3);
  wire        _GEN_36 = _GEN_32 & ~_GEN_34;
  wire        _GEN_38 = _slots_1_io_request & ~_GEN_30 & (|_can_allocate_T_6);
  wire        _GEN_40 = _GEN_38 & ~_GEN_22;
  wire        _GEN_42 = _slots_1_io_request & ~_GEN_28 & (|_GEN_23);
  wire        _GEN_44 = _GEN_42 & ~_GEN_24;
  wire        _GEN_13229 = _GEN_26 & ~_GEN_17;
  wire        issue_slots_1_grant = _GEN_36 | _GEN_40 | _GEN_44 | _GEN_13229;
  wire [9:0]  _can_allocate_T_14 = _slots_3_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_46 = {_slots_2_io_uop_fu_code[5], _slots_2_io_uop_fu_code[0]};
  wire        _GEN_48 = _GEN_42 | _GEN_24;
  wire        _GEN_50 = _slots_2_io_request & (|(_slots_2_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_52 = _GEN_26 | _GEN_17;
  wire        _GEN_54 = _GEN_50 & ~_GEN_52;
  wire        _GEN_56 = _slots_2_io_request & (|_GEN_46) & ~_GEN_48 | _GEN_54;
  wire [9:0]  _can_allocate_T_10 = _slots_2_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_58 = _slots_2_io_request & ~_GEN_56 & (|_can_allocate_T_10);
  wire        _GEN_60 = _GEN_38 | _GEN_22;
  wire        _GEN_62 = _GEN_58 | _GEN_60;
  wire [1:0]  _GEN_64 = {_slots_3_io_uop_fu_code[5], _slots_3_io_uop_fu_code[0]};
  wire        _GEN_66 = _slots_2_io_request & ~_GEN_54 & (|_GEN_46);
  wire        _GEN_68 = _GEN_66 | _GEN_48;
  wire        _GEN_70 = _slots_3_io_request & (|(_slots_3_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_72 = _GEN_50 | _GEN_52;
  wire        _GEN_74 = _GEN_70 & ~_GEN_72;
  wire        _GEN_76 = _slots_3_io_request & (|_GEN_64) & ~_GEN_68 | _GEN_74;
  wire        _GEN_78 = _slots_3_io_request & ~(_slots_3_io_request & (|_can_allocate_T_14) & ~_GEN_62 | _GEN_76) & (|(_slots_3_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_80 = _slots_2_io_request & ~(_slots_2_io_request & (|_can_allocate_T_10) & ~_GEN_60 | _GEN_56) & (|(_slots_2_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_82 = _GEN_32 | _GEN_34;
  wire        _GEN_84 = _GEN_80 | _GEN_82;
  wire        _GEN_86 = _GEN_78 & ~_GEN_84;
  wire        _GEN_88 = _slots_3_io_request & ~_GEN_76 & (|_can_allocate_T_14);
  wire        _GEN_90 = _GEN_88 & ~_GEN_62;
  wire        _GEN_92 = _slots_3_io_request & ~_GEN_74 & (|_GEN_64);
  wire        _GEN_94 = _GEN_92 & ~_GEN_68;
  wire        _GEN_13877 = _GEN_70 & ~_GEN_72;
  wire        issue_slots_3_grant = _GEN_86 | _GEN_90 | _GEN_94 | _GEN_13877;
  wire [9:0]  _can_allocate_T_18 = _slots_4_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_96 = _GEN_88 | _GEN_62;
  wire [1:0]  _GEN_98 = {_slots_4_io_uop_fu_code[5], _slots_4_io_uop_fu_code[0]};
  wire        _GEN_99 = _GEN_92 | _GEN_68;
  wire        _GEN_100 = _slots_4_io_request & (|(_slots_4_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_101 = _GEN_70 | _GEN_72;
  wire        _GEN_102 = _GEN_100 & ~_GEN_101;
  wire        _GEN_103 = _slots_4_io_request & (|_GEN_98) & ~_GEN_99 | _GEN_102;
  wire        _GEN_104 = _slots_4_io_request & ~(_slots_4_io_request & (|_can_allocate_T_18) & ~_GEN_96 | _GEN_103) & (|(_slots_4_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_105 = _GEN_78 | _GEN_84;
  wire        _GEN_106 = _GEN_104 & ~_GEN_105;
  wire        _GEN_107 = _slots_4_io_request & ~_GEN_103 & (|_can_allocate_T_18);
  wire        _GEN_108 = _GEN_107 & ~_GEN_96;
  wire        _GEN_109 = _slots_4_io_request & ~_GEN_102 & (|_GEN_98);
  wire        _GEN_110 = _GEN_109 & ~_GEN_99;
  wire        _GEN_14201 = _GEN_100 & ~_GEN_101;
  wire        issue_slots_4_grant = _GEN_106 | _GEN_108 | _GEN_110 | _GEN_14201;
  wire        _GEN_111 = _GEN_80 & ~_GEN_82;
  wire        _GEN_112 = _GEN_58 & ~_GEN_60;
  wire        _GEN_113 = _GEN_66 & ~_GEN_48;
  wire        _GEN_13553 = _GEN_50 & ~_GEN_52;
  wire        issue_slots_2_grant = _GEN_111 | _GEN_112 | _GEN_113 | _GEN_13553;
  wire [9:0]  _can_allocate_T_22 = _slots_5_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_114 = _GEN_107 | _GEN_96;
  wire [1:0]  _GEN_115 = {_slots_5_io_uop_fu_code[5], _slots_5_io_uop_fu_code[0]};
  wire        _GEN_116 = _GEN_109 | _GEN_99;
  wire        _GEN_117 = _slots_5_io_request & (|(_slots_5_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_118 = _GEN_100 | _GEN_101;
  wire        _GEN_119 = _GEN_117 & ~_GEN_118;
  wire        _GEN_120 = _slots_5_io_request & (|_GEN_115) & ~_GEN_116 | _GEN_119;
  wire        _GEN_121 = _slots_5_io_request & ~(_slots_5_io_request & (|_can_allocate_T_22) & ~_GEN_114 | _GEN_120) & (|(_slots_5_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_122 = _GEN_104 | _GEN_105;
  wire        _GEN_123 = _GEN_121 & ~_GEN_122;
  wire        _GEN_124 = _slots_5_io_request & ~_GEN_120 & (|_can_allocate_T_22);
  wire        _GEN_125 = _GEN_124 & ~_GEN_114;
  wire        _GEN_126 = _slots_5_io_request & ~_GEN_119 & (|_GEN_115);
  wire        _GEN_127 = _GEN_126 & ~_GEN_116;
  wire        _GEN_14525 = _GEN_117 & ~_GEN_118;
  wire        issue_slots_5_grant = _GEN_123 | _GEN_125 | _GEN_127 | _GEN_14525;
  wire [9:0]  _can_allocate_T_26 = _slots_6_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_128 = _GEN_124 | _GEN_114;
  wire [1:0]  _GEN_129 = {_slots_6_io_uop_fu_code[5], _slots_6_io_uop_fu_code[0]};
  wire        _GEN_130 = _GEN_126 | _GEN_116;
  wire        _GEN_131 = _slots_6_io_request & (|(_slots_6_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_132 = _GEN_117 | _GEN_118;
  wire        _GEN_133 = _GEN_131 & ~_GEN_132;
  wire        _GEN_134 = _slots_6_io_request & (|_GEN_129) & ~_GEN_130 | _GEN_133;
  wire        _GEN_135 = _slots_6_io_request & ~(_slots_6_io_request & (|_can_allocate_T_26) & ~_GEN_128 | _GEN_134) & (|(_slots_6_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_136 = _GEN_121 | _GEN_122;
  wire        _GEN_137 = _GEN_135 & ~_GEN_136;
  wire        _GEN_138 = _slots_6_io_request & ~_GEN_134 & (|_can_allocate_T_26);
  wire        _GEN_139 = _GEN_138 & ~_GEN_128;
  wire        _GEN_140 = _slots_6_io_request & ~_GEN_133 & (|_GEN_129);
  wire        _GEN_141 = _GEN_140 & ~_GEN_130;
  wire        _GEN_14849 = _GEN_131 & ~_GEN_132;
  wire        issue_slots_6_grant = _GEN_137 | _GEN_139 | _GEN_141 | _GEN_14849;
  wire [9:0]  _can_allocate_T_34 = _slots_8_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_142 = {_slots_7_io_uop_fu_code[5], _slots_7_io_uop_fu_code[0]};
  wire        _GEN_143 = _GEN_140 | _GEN_130;
  wire        _GEN_144 = _slots_7_io_request & (|(_slots_7_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_145 = _GEN_131 | _GEN_132;
  wire        _GEN_146 = _GEN_144 & ~_GEN_145;
  wire        _GEN_147 = _slots_7_io_request & (|_GEN_142) & ~_GEN_143 | _GEN_146;
  wire [9:0]  _can_allocate_T_30 = _slots_7_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_148 = _slots_7_io_request & ~_GEN_147 & (|_can_allocate_T_30);
  wire        _GEN_149 = _GEN_138 | _GEN_128;
  wire        _GEN_150 = _GEN_148 | _GEN_149;
  wire [1:0]  _GEN_151 = {_slots_8_io_uop_fu_code[5], _slots_8_io_uop_fu_code[0]};
  wire        _GEN_152 = _slots_7_io_request & ~_GEN_146 & (|_GEN_142);
  wire        _GEN_153 = _GEN_152 | _GEN_143;
  wire        _GEN_154 = _slots_8_io_request & (|(_slots_8_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_155 = _GEN_144 | _GEN_145;
  wire        _GEN_156 = _GEN_154 & ~_GEN_155;
  wire        _GEN_157 = _slots_8_io_request & (|_GEN_151) & ~_GEN_153 | _GEN_156;
  wire        _GEN_158 = _slots_8_io_request & ~(_slots_8_io_request & (|_can_allocate_T_34) & ~_GEN_150 | _GEN_157) & (|(_slots_8_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_159 = _slots_7_io_request & ~(_slots_7_io_request & (|_can_allocate_T_30) & ~_GEN_149 | _GEN_147) & (|(_slots_7_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_160 = _GEN_135 | _GEN_136;
  wire        _GEN_161 = _GEN_159 | _GEN_160;
  wire        _GEN_162 = _GEN_158 & ~_GEN_161;
  wire        _GEN_163 = _slots_8_io_request & ~_GEN_157 & (|_can_allocate_T_34);
  wire        _GEN_164 = _GEN_163 & ~_GEN_150;
  wire        _GEN_165 = _slots_8_io_request & ~_GEN_156 & (|_GEN_151);
  wire        _GEN_166 = _GEN_165 & ~_GEN_153;
  wire        _GEN_15497 = _GEN_154 & ~_GEN_155;
  wire        issue_slots_8_grant = _GEN_162 | _GEN_164 | _GEN_166 | _GEN_15497;
  wire [9:0]  _can_allocate_T_38 = _slots_9_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_167 = _GEN_163 | _GEN_150;
  wire [1:0]  _GEN_168 = {_slots_9_io_uop_fu_code[5], _slots_9_io_uop_fu_code[0]};
  wire        _GEN_169 = _GEN_165 | _GEN_153;
  wire        _GEN_170 = _slots_9_io_request & (|(_slots_9_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_171 = _GEN_154 | _GEN_155;
  wire        _GEN_172 = _GEN_170 & ~_GEN_171;
  wire        _GEN_173 = _slots_9_io_request & (|_GEN_168) & ~_GEN_169 | _GEN_172;
  wire        _GEN_174 = _slots_9_io_request & ~(_slots_9_io_request & (|_can_allocate_T_38) & ~_GEN_167 | _GEN_173) & (|(_slots_9_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_175 = _GEN_158 | _GEN_161;
  wire        _GEN_176 = _GEN_174 & ~_GEN_175;
  wire        _GEN_177 = _slots_9_io_request & ~_GEN_173 & (|_can_allocate_T_38);
  wire        _GEN_178 = _GEN_177 & ~_GEN_167;
  wire        _GEN_179 = _slots_9_io_request & ~_GEN_172 & (|_GEN_168);
  wire        _GEN_180 = _GEN_179 & ~_GEN_169;
  wire        _GEN_15821 = _GEN_170 & ~_GEN_171;
  wire        issue_slots_9_grant = _GEN_176 | _GEN_178 | _GEN_180 | _GEN_15821;
  wire        _GEN_181 = _GEN_159 & ~_GEN_160;
  wire        _GEN_182 = _GEN_148 & ~_GEN_149;
  wire        _GEN_183 = _GEN_152 & ~_GEN_143;
  wire        _GEN_15173 = _GEN_144 & ~_GEN_145;
  wire        issue_slots_7_grant = _GEN_181 | _GEN_182 | _GEN_183 | _GEN_15173;
  wire [9:0]  _can_allocate_T_42 = _slots_10_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_184 = _GEN_177 | _GEN_167;
  wire [1:0]  _GEN_185 = {_slots_10_io_uop_fu_code[5], _slots_10_io_uop_fu_code[0]};
  wire        _GEN_186 = _GEN_179 | _GEN_169;
  wire        _GEN_187 = _slots_10_io_request & (|(_slots_10_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_188 = _GEN_170 | _GEN_171;
  wire        _GEN_189 = _GEN_187 & ~_GEN_188;
  wire        _GEN_190 = _slots_10_io_request & (|_GEN_185) & ~_GEN_186 | _GEN_189;
  wire        _GEN_191 = _slots_10_io_request & ~(_slots_10_io_request & (|_can_allocate_T_42) & ~_GEN_184 | _GEN_190) & (|(_slots_10_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_192 = _GEN_174 | _GEN_175;
  wire        _GEN_193 = _GEN_191 & ~_GEN_192;
  wire        _GEN_194 = _slots_10_io_request & ~_GEN_190 & (|_can_allocate_T_42);
  wire        _GEN_195 = _GEN_194 & ~_GEN_184;
  wire        _GEN_196 = _slots_10_io_request & ~_GEN_189 & (|_GEN_185);
  wire        _GEN_197 = _GEN_196 & ~_GEN_186;
  wire        _GEN_16145 = _GEN_187 & ~_GEN_188;
  wire        issue_slots_10_grant = _GEN_193 | _GEN_195 | _GEN_197 | _GEN_16145;
  wire [9:0]  _can_allocate_T_46 = _slots_11_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_198 = _GEN_194 | _GEN_184;
  wire [1:0]  _GEN_199 = {_slots_11_io_uop_fu_code[5], _slots_11_io_uop_fu_code[0]};
  wire        _GEN_200 = _GEN_196 | _GEN_186;
  wire        _GEN_201 = _slots_11_io_request & (|(_slots_11_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_202 = _GEN_187 | _GEN_188;
  wire        _GEN_203 = _GEN_201 & ~_GEN_202;
  wire        _GEN_204 = _slots_11_io_request & (|_GEN_199) & ~_GEN_200 | _GEN_203;
  wire        _GEN_205 = _slots_11_io_request & ~(_slots_11_io_request & (|_can_allocate_T_46) & ~_GEN_198 | _GEN_204) & (|(_slots_11_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_206 = _GEN_191 | _GEN_192;
  wire        _GEN_207 = _GEN_205 & ~_GEN_206;
  wire        _GEN_208 = _slots_11_io_request & ~_GEN_204 & (|_can_allocate_T_46);
  wire        _GEN_209 = _GEN_208 & ~_GEN_198;
  wire        _GEN_210 = _slots_11_io_request & ~_GEN_203 & (|_GEN_199);
  wire        _GEN_211 = _GEN_210 & ~_GEN_200;
  wire        _GEN_16469 = _GEN_201 & ~_GEN_202;
  wire        issue_slots_11_grant = _GEN_207 | _GEN_209 | _GEN_211 | _GEN_16469;
  wire [9:0]  _can_allocate_T_54 = _slots_13_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_212 = {_slots_12_io_uop_fu_code[5], _slots_12_io_uop_fu_code[0]};
  wire        _GEN_213 = _GEN_210 | _GEN_200;
  wire        _GEN_214 = _slots_12_io_request & (|(_slots_12_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_215 = _GEN_201 | _GEN_202;
  wire        _GEN_216 = _GEN_214 & ~_GEN_215;
  wire        _GEN_217 = _slots_12_io_request & (|_GEN_212) & ~_GEN_213 | _GEN_216;
  wire [9:0]  _can_allocate_T_50 = _slots_12_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_218 = _slots_12_io_request & ~_GEN_217 & (|_can_allocate_T_50);
  wire        _GEN_219 = _GEN_208 | _GEN_198;
  wire        _GEN_220 = _GEN_218 | _GEN_219;
  wire [1:0]  _GEN_221 = {_slots_13_io_uop_fu_code[5], _slots_13_io_uop_fu_code[0]};
  wire        _GEN_222 = _slots_12_io_request & ~_GEN_216 & (|_GEN_212);
  wire        _GEN_223 = _GEN_222 | _GEN_213;
  wire        _GEN_224 = _slots_13_io_request & (|(_slots_13_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_225 = _GEN_214 | _GEN_215;
  wire        _GEN_226 = _GEN_224 & ~_GEN_225;
  wire        _GEN_227 = _slots_13_io_request & (|_GEN_221) & ~_GEN_223 | _GEN_226;
  wire        _GEN_228 = _slots_13_io_request & ~(_slots_13_io_request & (|_can_allocate_T_54) & ~_GEN_220 | _GEN_227) & (|(_slots_13_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_229 = _slots_12_io_request & ~(_slots_12_io_request & (|_can_allocate_T_50) & ~_GEN_219 | _GEN_217) & (|(_slots_12_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_230 = _GEN_205 | _GEN_206;
  wire        _GEN_231 = _GEN_229 | _GEN_230;
  wire        _GEN_232 = _GEN_228 & ~_GEN_231;
  wire        _GEN_233 = _slots_13_io_request & ~_GEN_227 & (|_can_allocate_T_54);
  wire        _GEN_234 = _GEN_233 & ~_GEN_220;
  wire        _GEN_235 = _slots_13_io_request & ~_GEN_226 & (|_GEN_221);
  wire        _GEN_236 = _GEN_235 & ~_GEN_223;
  wire        _GEN_17117 = _GEN_224 & ~_GEN_225;
  wire        issue_slots_13_grant = _GEN_232 | _GEN_234 | _GEN_236 | _GEN_17117;
  wire [9:0]  _can_allocate_T_58 = _slots_14_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_237 = _GEN_233 | _GEN_220;
  wire [1:0]  _GEN_238 = {_slots_14_io_uop_fu_code[5], _slots_14_io_uop_fu_code[0]};
  wire        _GEN_239 = _GEN_235 | _GEN_223;
  wire        _GEN_240 = _slots_14_io_request & (|(_slots_14_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_241 = _GEN_224 | _GEN_225;
  wire        _GEN_242 = _GEN_240 & ~_GEN_241;
  wire        _GEN_243 = _slots_14_io_request & (|_GEN_238) & ~_GEN_239 | _GEN_242;
  wire        _GEN_244 = _slots_14_io_request & ~(_slots_14_io_request & (|_can_allocate_T_58) & ~_GEN_237 | _GEN_243) & (|(_slots_14_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_245 = _GEN_228 | _GEN_231;
  wire        _GEN_246 = _GEN_244 & ~_GEN_245;
  wire        _GEN_247 = _slots_14_io_request & ~_GEN_243 & (|_can_allocate_T_58);
  wire        _GEN_248 = _GEN_247 & ~_GEN_237;
  wire        _GEN_249 = _slots_14_io_request & ~_GEN_242 & (|_GEN_238);
  wire        _GEN_250 = _GEN_249 & ~_GEN_239;
  wire        _GEN_17441 = _GEN_240 & ~_GEN_241;
  wire        issue_slots_14_grant = _GEN_246 | _GEN_248 | _GEN_250 | _GEN_17441;
  wire        _GEN_251 = _GEN_229 & ~_GEN_230;
  wire        _GEN_252 = _GEN_218 & ~_GEN_219;
  wire        _GEN_253 = _GEN_222 & ~_GEN_213;
  wire        _GEN_16793 = _GEN_214 & ~_GEN_215;
  wire        issue_slots_12_grant = _GEN_251 | _GEN_252 | _GEN_253 | _GEN_16793;
  wire [9:0]  _can_allocate_T_62 = _slots_15_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_254 = _GEN_247 | _GEN_237;
  wire [1:0]  _GEN_255 = {_slots_15_io_uop_fu_code[5], _slots_15_io_uop_fu_code[0]};
  wire        _GEN_256 = _GEN_249 | _GEN_239;
  wire        _GEN_257 = _slots_15_io_request & (|(_slots_15_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_258 = _GEN_240 | _GEN_241;
  wire        _GEN_259 = _GEN_257 & ~_GEN_258;
  wire        _GEN_260 = _slots_15_io_request & (|_GEN_255) & ~_GEN_256 | _GEN_259;
  wire        _GEN_261 = _slots_15_io_request & ~(_slots_15_io_request & (|_can_allocate_T_62) & ~_GEN_254 | _GEN_260) & (|(_slots_15_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_262 = _GEN_244 | _GEN_245;
  wire        _GEN_263 = _GEN_261 & ~_GEN_262;
  wire        _GEN_264 = _slots_15_io_request & ~_GEN_260 & (|_can_allocate_T_62);
  wire        _GEN_265 = _GEN_264 & ~_GEN_254;
  wire        _GEN_266 = _slots_15_io_request & ~_GEN_259 & (|_GEN_255);
  wire        _GEN_267 = _GEN_266 & ~_GEN_256;
  wire        _GEN_17765 = _GEN_257 & ~_GEN_258;
  wire        issue_slots_15_grant = _GEN_263 | _GEN_265 | _GEN_267 | _GEN_17765;
  wire [9:0]  _can_allocate_T_66 = _slots_16_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_268 = _GEN_264 | _GEN_254;
  wire [1:0]  _GEN_269 = {_slots_16_io_uop_fu_code[5], _slots_16_io_uop_fu_code[0]};
  wire        _GEN_270 = _GEN_266 | _GEN_256;
  wire        _GEN_271 = _slots_16_io_request & (|(_slots_16_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_272 = _GEN_257 | _GEN_258;
  wire        _GEN_273 = _GEN_271 & ~_GEN_272;
  wire        _GEN_274 = _slots_16_io_request & (|_GEN_269) & ~_GEN_270 | _GEN_273;
  wire        _GEN_275 = _slots_16_io_request & ~(_slots_16_io_request & (|_can_allocate_T_66) & ~_GEN_268 | _GEN_274) & (|(_slots_16_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_276 = _GEN_261 | _GEN_262;
  wire        _GEN_277 = _GEN_275 & ~_GEN_276;
  wire        _GEN_278 = _slots_16_io_request & ~_GEN_274 & (|_can_allocate_T_66);
  wire        _GEN_279 = _GEN_278 & ~_GEN_268;
  wire        _GEN_280 = _slots_16_io_request & ~_GEN_273 & (|_GEN_269);
  wire        _GEN_281 = _GEN_280 & ~_GEN_270;
  wire        _GEN_18089 = _GEN_271 & ~_GEN_272;
  wire        issue_slots_16_grant = _GEN_277 | _GEN_279 | _GEN_281 | _GEN_18089;
  wire [9:0]  _can_allocate_T_74 = _slots_18_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_282 = {_slots_17_io_uop_fu_code[5], _slots_17_io_uop_fu_code[0]};
  wire        _GEN_283 = _GEN_280 | _GEN_270;
  wire        _GEN_284 = _slots_17_io_request & (|(_slots_17_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_285 = _GEN_271 | _GEN_272;
  wire        _GEN_286 = _GEN_284 & ~_GEN_285;
  wire        _GEN_287 = _slots_17_io_request & (|_GEN_282) & ~_GEN_283 | _GEN_286;
  wire [9:0]  _can_allocate_T_70 = _slots_17_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_288 = _slots_17_io_request & ~_GEN_287 & (|_can_allocate_T_70);
  wire        _GEN_289 = _GEN_278 | _GEN_268;
  wire        _GEN_290 = _GEN_288 | _GEN_289;
  wire [1:0]  _GEN_291 = {_slots_18_io_uop_fu_code[5], _slots_18_io_uop_fu_code[0]};
  wire        _GEN_292 = _slots_17_io_request & ~_GEN_286 & (|_GEN_282);
  wire        _GEN_293 = _GEN_292 | _GEN_283;
  wire        _GEN_294 = _slots_18_io_request & (|(_slots_18_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_295 = _GEN_284 | _GEN_285;
  wire        _GEN_296 = _GEN_294 & ~_GEN_295;
  wire        _GEN_297 = _slots_18_io_request & (|_GEN_291) & ~_GEN_293 | _GEN_296;
  wire        _GEN_298 = _slots_18_io_request & ~(_slots_18_io_request & (|_can_allocate_T_74) & ~_GEN_290 | _GEN_297) & (|(_slots_18_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_299 = _slots_17_io_request & ~(_slots_17_io_request & (|_can_allocate_T_70) & ~_GEN_289 | _GEN_287) & (|(_slots_17_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_300 = _GEN_275 | _GEN_276;
  wire        _GEN_301 = _GEN_299 | _GEN_300;
  wire        _GEN_302 = _GEN_298 & ~_GEN_301;
  wire        _GEN_303 = _slots_18_io_request & ~_GEN_297 & (|_can_allocate_T_74);
  wire        _GEN_304 = _GEN_303 & ~_GEN_290;
  wire        _GEN_305 = _slots_18_io_request & ~_GEN_296 & (|_GEN_291);
  wire        _GEN_306 = _GEN_305 & ~_GEN_293;
  wire        _GEN_18737 = _GEN_294 & ~_GEN_295;
  wire        issue_slots_18_grant = _GEN_302 | _GEN_304 | _GEN_306 | _GEN_18737;
  wire [9:0]  _can_allocate_T_78 = _slots_19_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_307 = _GEN_303 | _GEN_290;
  wire [1:0]  _GEN_308 = {_slots_19_io_uop_fu_code[5], _slots_19_io_uop_fu_code[0]};
  wire        _GEN_309 = _GEN_305 | _GEN_293;
  wire        _GEN_310 = _slots_19_io_request & (|(_slots_19_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_311 = _GEN_294 | _GEN_295;
  wire        _GEN_312 = _GEN_310 & ~_GEN_311;
  wire        _GEN_313 = _slots_19_io_request & (|_GEN_308) & ~_GEN_309 | _GEN_312;
  wire        _GEN_314 = _slots_19_io_request & ~(_slots_19_io_request & (|_can_allocate_T_78) & ~_GEN_307 | _GEN_313) & (|(_slots_19_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_315 = _GEN_298 | _GEN_301;
  wire        _GEN_316 = _GEN_314 & ~_GEN_315;
  wire        _GEN_317 = _slots_19_io_request & ~_GEN_313 & (|_can_allocate_T_78);
  wire        _GEN_318 = _GEN_317 & ~_GEN_307;
  wire        _GEN_319 = _slots_19_io_request & ~_GEN_312 & (|_GEN_308);
  wire        _GEN_320 = _GEN_319 & ~_GEN_309;
  wire        _GEN_19061 = _GEN_310 & ~_GEN_311;
  wire        issue_slots_19_grant = _GEN_316 | _GEN_318 | _GEN_320 | _GEN_19061;
  wire        _GEN_321 = _GEN_299 & ~_GEN_300;
  wire        _GEN_322 = _GEN_288 & ~_GEN_289;
  wire        _GEN_323 = _GEN_292 & ~_GEN_283;
  wire        _GEN_18413 = _GEN_284 & ~_GEN_285;
  wire        issue_slots_17_grant = _GEN_321 | _GEN_322 | _GEN_323 | _GEN_18413;
  wire [9:0]  _can_allocate_T_82 = _slots_20_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_324 = _GEN_317 | _GEN_307;
  wire [1:0]  _GEN_325 = {_slots_20_io_uop_fu_code[5], _slots_20_io_uop_fu_code[0]};
  wire        _GEN_326 = _GEN_319 | _GEN_309;
  wire        _GEN_327 = _slots_20_io_request & (|(_slots_20_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_328 = _GEN_310 | _GEN_311;
  wire        _GEN_329 = _GEN_327 & ~_GEN_328;
  wire        _GEN_330 = _slots_20_io_request & (|_GEN_325) & ~_GEN_326 | _GEN_329;
  wire        _GEN_331 = _slots_20_io_request & ~(_slots_20_io_request & (|_can_allocate_T_82) & ~_GEN_324 | _GEN_330) & (|(_slots_20_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_332 = _GEN_314 | _GEN_315;
  wire        _GEN_333 = _GEN_331 & ~_GEN_332;
  wire        _GEN_334 = _slots_20_io_request & ~_GEN_330 & (|_can_allocate_T_82);
  wire        _GEN_335 = _GEN_334 & ~_GEN_324;
  wire        _GEN_336 = _slots_20_io_request & ~_GEN_329 & (|_GEN_325);
  wire        _GEN_337 = _GEN_336 & ~_GEN_326;
  wire        _GEN_19385 = _GEN_327 & ~_GEN_328;
  wire        issue_slots_20_grant = _GEN_333 | _GEN_335 | _GEN_337 | _GEN_19385;
  wire [9:0]  _can_allocate_T_86 = _slots_21_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_338 = _GEN_334 | _GEN_324;
  wire [1:0]  _GEN_339 = {_slots_21_io_uop_fu_code[5], _slots_21_io_uop_fu_code[0]};
  wire        _GEN_340 = _GEN_336 | _GEN_326;
  wire        _GEN_341 = _slots_21_io_request & (|(_slots_21_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_342 = _GEN_327 | _GEN_328;
  wire        _GEN_343 = _GEN_341 & ~_GEN_342;
  wire        _GEN_344 = _slots_21_io_request & (|_GEN_339) & ~_GEN_340 | _GEN_343;
  wire        _GEN_345 = _slots_21_io_request & ~(_slots_21_io_request & (|_can_allocate_T_86) & ~_GEN_338 | _GEN_344) & (|(_slots_21_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_346 = _GEN_331 | _GEN_332;
  wire        _GEN_347 = _GEN_345 & ~_GEN_346;
  wire        _GEN_348 = _slots_21_io_request & ~_GEN_344 & (|_can_allocate_T_86);
  wire        _GEN_349 = _GEN_348 & ~_GEN_338;
  wire        _GEN_350 = _slots_21_io_request & ~_GEN_343 & (|_GEN_339);
  wire        _GEN_351 = _GEN_350 & ~_GEN_340;
  wire        _GEN_19709 = _GEN_341 & ~_GEN_342;
  wire        issue_slots_21_grant = _GEN_347 | _GEN_349 | _GEN_351 | _GEN_19709;
  wire [9:0]  _can_allocate_T_94 = _slots_23_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_352 = {_slots_22_io_uop_fu_code[5], _slots_22_io_uop_fu_code[0]};
  wire        _GEN_353 = _GEN_350 | _GEN_340;
  wire        _GEN_354 = _slots_22_io_request & (|(_slots_22_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_355 = _GEN_341 | _GEN_342;
  wire        _GEN_356 = _GEN_354 & ~_GEN_355;
  wire        _GEN_357 = _slots_22_io_request & (|_GEN_352) & ~_GEN_353 | _GEN_356;
  wire [9:0]  _can_allocate_T_90 = _slots_22_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_358 = _slots_22_io_request & ~_GEN_357 & (|_can_allocate_T_90);
  wire        _GEN_359 = _GEN_348 | _GEN_338;
  wire        _GEN_360 = _GEN_358 | _GEN_359;
  wire [1:0]  _GEN_361 = {_slots_23_io_uop_fu_code[5], _slots_23_io_uop_fu_code[0]};
  wire        _GEN_362 = _slots_22_io_request & ~_GEN_356 & (|_GEN_352);
  wire        _GEN_363 = _GEN_362 | _GEN_353;
  wire        _GEN_364 = _slots_23_io_request & (|(_slots_23_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_365 = _GEN_354 | _GEN_355;
  wire        _GEN_366 = _GEN_364 & ~_GEN_365;
  wire        _GEN_367 = _slots_23_io_request & (|_GEN_361) & ~_GEN_363 | _GEN_366;
  wire        _GEN_368 = _slots_23_io_request & ~(_slots_23_io_request & (|_can_allocate_T_94) & ~_GEN_360 | _GEN_367) & (|(_slots_23_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_369 = _slots_22_io_request & ~(_slots_22_io_request & (|_can_allocate_T_90) & ~_GEN_359 | _GEN_357) & (|(_slots_22_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_370 = _GEN_345 | _GEN_346;
  wire        _GEN_371 = _GEN_369 | _GEN_370;
  wire        _GEN_372 = _GEN_368 & ~_GEN_371;
  wire        _GEN_373 = _slots_23_io_request & ~_GEN_367 & (|_can_allocate_T_94);
  wire        _GEN_374 = _GEN_373 & ~_GEN_360;
  wire        _GEN_375 = _slots_23_io_request & ~_GEN_366 & (|_GEN_361);
  wire        _GEN_376 = _GEN_375 & ~_GEN_363;
  wire        _GEN_20357 = _GEN_364 & ~_GEN_365;
  wire        issue_slots_23_grant = _GEN_372 | _GEN_374 | _GEN_376 | _GEN_20357;
  wire [9:0]  _can_allocate_T_98 = _slots_24_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_377 = _GEN_373 | _GEN_360;
  wire [1:0]  _GEN_378 = {_slots_24_io_uop_fu_code[5], _slots_24_io_uop_fu_code[0]};
  wire        _GEN_379 = _GEN_375 | _GEN_363;
  wire        _GEN_380 = _slots_24_io_request & (|(_slots_24_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_381 = _GEN_364 | _GEN_365;
  wire        _GEN_382 = _GEN_380 & ~_GEN_381;
  wire        _GEN_383 = _slots_24_io_request & (|_GEN_378) & ~_GEN_379 | _GEN_382;
  wire        _GEN_384 = _slots_24_io_request & ~(_slots_24_io_request & (|_can_allocate_T_98) & ~_GEN_377 | _GEN_383) & (|(_slots_24_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_385 = _GEN_368 | _GEN_371;
  wire        _GEN_386 = _GEN_384 & ~_GEN_385;
  wire        _GEN_387 = _slots_24_io_request & ~_GEN_383 & (|_can_allocate_T_98);
  wire        _GEN_388 = _GEN_387 & ~_GEN_377;
  wire        _GEN_389 = _slots_24_io_request & ~_GEN_382 & (|_GEN_378);
  wire        _GEN_390 = _GEN_389 & ~_GEN_379;
  wire        _GEN_20681 = _GEN_380 & ~_GEN_381;
  wire        issue_slots_24_grant = _GEN_386 | _GEN_388 | _GEN_390 | _GEN_20681;
  wire        _GEN_391 = _GEN_369 & ~_GEN_370;
  wire        _GEN_392 = _GEN_358 & ~_GEN_359;
  wire        _GEN_393 = _GEN_362 & ~_GEN_353;
  wire        _GEN_20033 = _GEN_354 & ~_GEN_355;
  wire        issue_slots_22_grant = _GEN_391 | _GEN_392 | _GEN_393 | _GEN_20033;
  wire [9:0]  _can_allocate_T_102 = _slots_25_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_394 = _GEN_387 | _GEN_377;
  wire [1:0]  _GEN_395 = {_slots_25_io_uop_fu_code[5], _slots_25_io_uop_fu_code[0]};
  wire        _GEN_396 = _GEN_389 | _GEN_379;
  wire        _GEN_397 = _slots_25_io_request & (|(_slots_25_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_398 = _GEN_380 | _GEN_381;
  wire        _GEN_399 = _GEN_397 & ~_GEN_398;
  wire        _GEN_400 = _slots_25_io_request & (|_GEN_395) & ~_GEN_396 | _GEN_399;
  wire        _GEN_401 = _slots_25_io_request & ~(_slots_25_io_request & (|_can_allocate_T_102) & ~_GEN_394 | _GEN_400) & (|(_slots_25_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_402 = _GEN_384 | _GEN_385;
  wire        _GEN_403 = _GEN_401 & ~_GEN_402;
  wire        _GEN_404 = _slots_25_io_request & ~_GEN_400 & (|_can_allocate_T_102);
  wire        _GEN_405 = _GEN_404 & ~_GEN_394;
  wire        _GEN_406 = _slots_25_io_request & ~_GEN_399 & (|_GEN_395);
  wire        _GEN_407 = _GEN_406 & ~_GEN_396;
  wire        _GEN_21005 = _GEN_397 & ~_GEN_398;
  wire        issue_slots_25_grant = _GEN_403 | _GEN_405 | _GEN_407 | _GEN_21005;
  wire [9:0]  _can_allocate_T_106 = _slots_26_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_408 = _GEN_404 | _GEN_394;
  wire [1:0]  _GEN_409 = {_slots_26_io_uop_fu_code[5], _slots_26_io_uop_fu_code[0]};
  wire        _GEN_410 = _GEN_406 | _GEN_396;
  wire        _GEN_411 = _slots_26_io_request & (|(_slots_26_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_412 = _GEN_397 | _GEN_398;
  wire        _GEN_413 = _GEN_411 & ~_GEN_412;
  wire        _GEN_414 = _slots_26_io_request & (|_GEN_409) & ~_GEN_410 | _GEN_413;
  wire        _GEN_415 = _slots_26_io_request & ~(_slots_26_io_request & (|_can_allocate_T_106) & ~_GEN_408 | _GEN_414) & (|(_slots_26_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_416 = _GEN_401 | _GEN_402;
  wire        _GEN_417 = _GEN_415 & ~_GEN_416;
  wire        _GEN_418 = _slots_26_io_request & ~_GEN_414 & (|_can_allocate_T_106);
  wire        _GEN_419 = _GEN_418 & ~_GEN_408;
  wire        _GEN_420 = _slots_26_io_request & ~_GEN_413 & (|_GEN_409);
  wire        _GEN_421 = _GEN_420 & ~_GEN_410;
  wire        _GEN_21329 = _GEN_411 & ~_GEN_412;
  wire        issue_slots_26_grant = _GEN_417 | _GEN_419 | _GEN_421 | _GEN_21329;
  wire [9:0]  _can_allocate_T_114 = _slots_28_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_422 = {_slots_27_io_uop_fu_code[5], _slots_27_io_uop_fu_code[0]};
  wire        _GEN_423 = _GEN_420 | _GEN_410;
  wire        _GEN_424 = _slots_27_io_request & (|(_slots_27_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_425 = _GEN_411 | _GEN_412;
  wire        _GEN_426 = _GEN_424 & ~_GEN_425;
  wire        _GEN_427 = _slots_27_io_request & (|_GEN_422) & ~_GEN_423 | _GEN_426;
  wire [9:0]  _can_allocate_T_110 = _slots_27_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_428 = _slots_27_io_request & ~_GEN_427 & (|_can_allocate_T_110);
  wire        _GEN_429 = _GEN_418 | _GEN_408;
  wire        _GEN_430 = _GEN_428 | _GEN_429;
  wire [1:0]  _GEN_431 = {_slots_28_io_uop_fu_code[5], _slots_28_io_uop_fu_code[0]};
  wire        _GEN_432 = _slots_27_io_request & ~_GEN_426 & (|_GEN_422);
  wire        _GEN_433 = _GEN_432 | _GEN_423;
  wire        _GEN_434 = _slots_28_io_request & (|(_slots_28_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_435 = _GEN_424 | _GEN_425;
  wire        _GEN_436 = _GEN_434 & ~_GEN_435;
  wire        _GEN_437 = _slots_28_io_request & (|_GEN_431) & ~_GEN_433 | _GEN_436;
  wire        _GEN_438 = _slots_28_io_request & ~(_slots_28_io_request & (|_can_allocate_T_114) & ~_GEN_430 | _GEN_437) & (|(_slots_28_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_439 = _slots_27_io_request & ~(_slots_27_io_request & (|_can_allocate_T_110) & ~_GEN_429 | _GEN_427) & (|(_slots_27_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_440 = _GEN_415 | _GEN_416;
  wire        _GEN_441 = _GEN_439 | _GEN_440;
  wire        _GEN_442 = _GEN_438 & ~_GEN_441;
  wire        _GEN_443 = _slots_28_io_request & ~_GEN_437 & (|_can_allocate_T_114);
  wire        _GEN_444 = _GEN_443 & ~_GEN_430;
  wire        _GEN_445 = _slots_28_io_request & ~_GEN_436 & (|_GEN_431);
  wire        _GEN_446 = _GEN_445 & ~_GEN_433;
  wire        _GEN_21977 = _GEN_434 & ~_GEN_435;
  wire        issue_slots_28_grant = _GEN_442 | _GEN_444 | _GEN_446 | _GEN_21977;
  wire [9:0]  _can_allocate_T_118 = _slots_29_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_447 = _GEN_443 | _GEN_430;
  wire [1:0]  _GEN_448 = {_slots_29_io_uop_fu_code[5], _slots_29_io_uop_fu_code[0]};
  wire        _GEN_449 = _GEN_445 | _GEN_433;
  wire        _GEN_450 = _slots_29_io_request & (|(_slots_29_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_451 = _GEN_434 | _GEN_435;
  wire        _GEN_452 = _GEN_450 & ~_GEN_451;
  wire        _GEN_453 = _slots_29_io_request & (|_GEN_448) & ~_GEN_449 | _GEN_452;
  wire        _GEN_454 = _slots_29_io_request & ~(_slots_29_io_request & (|_can_allocate_T_118) & ~_GEN_447 | _GEN_453) & (|(_slots_29_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_455 = _GEN_438 | _GEN_441;
  wire        _GEN_456 = _GEN_454 & ~_GEN_455;
  wire        _GEN_457 = _slots_29_io_request & ~_GEN_453 & (|_can_allocate_T_118);
  wire        _GEN_458 = _GEN_457 & ~_GEN_447;
  wire        _GEN_459 = _slots_29_io_request & ~_GEN_452 & (|_GEN_448);
  wire        _GEN_460 = _GEN_459 & ~_GEN_449;
  wire        _GEN_22301 = _GEN_450 & ~_GEN_451;
  wire        issue_slots_29_grant = _GEN_456 | _GEN_458 | _GEN_460 | _GEN_22301;
  wire        _GEN_461 = _GEN_439 & ~_GEN_440;
  wire        _GEN_462 = _GEN_428 & ~_GEN_429;
  wire        _GEN_463 = _GEN_432 & ~_GEN_423;
  wire        _GEN_21653 = _GEN_424 & ~_GEN_425;
  wire        issue_slots_27_grant = _GEN_461 | _GEN_462 | _GEN_463 | _GEN_21653;
  wire [9:0]  _can_allocate_T_122 = _slots_30_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_464 = _GEN_457 | _GEN_447;
  wire [1:0]  _GEN_465 = {_slots_30_io_uop_fu_code[5], _slots_30_io_uop_fu_code[0]};
  wire        _GEN_466 = _GEN_459 | _GEN_449;
  wire        _GEN_467 = _slots_30_io_request & (|(_slots_30_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_468 = _GEN_450 | _GEN_451;
  wire        _GEN_469 = _GEN_467 & ~_GEN_468;
  wire        _GEN_470 = _slots_30_io_request & (|_GEN_465) & ~_GEN_466 | _GEN_469;
  wire        _GEN_471 = _slots_30_io_request & ~(_slots_30_io_request & (|_can_allocate_T_122) & ~_GEN_464 | _GEN_470) & (|(_slots_30_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_472 = _GEN_454 | _GEN_455;
  wire        _GEN_473 = _GEN_471 & ~_GEN_472;
  wire        _GEN_474 = _slots_30_io_request & ~_GEN_470 & (|_can_allocate_T_122);
  wire        _GEN_475 = _GEN_474 & ~_GEN_464;
  wire        _GEN_476 = _slots_30_io_request & ~_GEN_469 & (|_GEN_465);
  wire        _GEN_477 = _GEN_476 & ~_GEN_466;
  wire        _GEN_22625 = _GEN_467 & ~_GEN_468;
  wire        issue_slots_30_grant = _GEN_473 | _GEN_475 | _GEN_477 | _GEN_22625;
  wire [9:0]  _can_allocate_T_126 = _slots_31_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_478 = _GEN_474 | _GEN_464;
  wire [1:0]  _GEN_479 = {_slots_31_io_uop_fu_code[5], _slots_31_io_uop_fu_code[0]};
  wire        _GEN_480 = _GEN_476 | _GEN_466;
  wire        _GEN_481 = _slots_31_io_request & (|(_slots_31_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_482 = _GEN_467 | _GEN_468;
  wire        _GEN_483 = _GEN_481 & ~_GEN_482;
  wire        _GEN_484 = _slots_31_io_request & (|_GEN_479) & ~_GEN_480 | _GEN_483;
  wire        _GEN_485 = _slots_31_io_request & ~(_slots_31_io_request & (|_can_allocate_T_126) & ~_GEN_478 | _GEN_484) & (|(_slots_31_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_486 = _GEN_471 | _GEN_472;
  wire        _GEN_487 = _GEN_485 & ~_GEN_486;
  wire        _GEN_488 = _slots_31_io_request & ~_GEN_484 & (|_can_allocate_T_126);
  wire        _GEN_489 = _GEN_488 & ~_GEN_478;
  wire        _GEN_490 = _slots_31_io_request & ~_GEN_483 & (|_GEN_479);
  wire        _GEN_491 = _GEN_490 & ~_GEN_480;
  wire        _GEN_22949 = _GEN_481 & ~_GEN_482;
  wire        issue_slots_31_grant = _GEN_487 | _GEN_489 | _GEN_491 | _GEN_22949;
  wire [9:0]  _can_allocate_T_134 = _slots_33_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_492 = {_slots_32_io_uop_fu_code[5], _slots_32_io_uop_fu_code[0]};
  wire        _GEN_493 = _GEN_490 | _GEN_480;
  wire        _GEN_494 = _slots_32_io_request & (|(_slots_32_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_495 = _GEN_481 | _GEN_482;
  wire        _GEN_496 = _GEN_494 & ~_GEN_495;
  wire        _GEN_497 = _slots_32_io_request & (|_GEN_492) & ~_GEN_493 | _GEN_496;
  wire [9:0]  _can_allocate_T_130 = _slots_32_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_498 = _slots_32_io_request & ~_GEN_497 & (|_can_allocate_T_130);
  wire        _GEN_499 = _GEN_488 | _GEN_478;
  wire        _GEN_500 = _GEN_498 | _GEN_499;
  wire [1:0]  _GEN_501 = {_slots_33_io_uop_fu_code[5], _slots_33_io_uop_fu_code[0]};
  wire        _GEN_502 = _slots_32_io_request & ~_GEN_496 & (|_GEN_492);
  wire        _GEN_503 = _GEN_502 | _GEN_493;
  wire        _GEN_504 = _slots_33_io_request & (|(_slots_33_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_505 = _GEN_494 | _GEN_495;
  wire        _GEN_506 = _GEN_504 & ~_GEN_505;
  wire        _GEN_507 = _slots_33_io_request & (|_GEN_501) & ~_GEN_503 | _GEN_506;
  wire        _GEN_508 = _slots_33_io_request & ~(_slots_33_io_request & (|_can_allocate_T_134) & ~_GEN_500 | _GEN_507) & (|(_slots_33_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_509 = _slots_32_io_request & ~(_slots_32_io_request & (|_can_allocate_T_130) & ~_GEN_499 | _GEN_497) & (|(_slots_32_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_510 = _GEN_485 | _GEN_486;
  wire        _GEN_511 = _GEN_509 | _GEN_510;
  wire        _GEN_512 = _GEN_508 & ~_GEN_511;
  wire        _GEN_513 = _slots_33_io_request & ~_GEN_507 & (|_can_allocate_T_134);
  wire        _GEN_514 = _GEN_513 & ~_GEN_500;
  wire        _GEN_515 = _slots_33_io_request & ~_GEN_506 & (|_GEN_501);
  wire        _GEN_516 = _GEN_515 & ~_GEN_503;
  wire        _GEN_23597 = _GEN_504 & ~_GEN_505;
  wire        issue_slots_33_grant = _GEN_512 | _GEN_514 | _GEN_516 | _GEN_23597;
  wire [9:0]  _can_allocate_T_138 = _slots_34_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_517 = _GEN_513 | _GEN_500;
  wire [1:0]  _GEN_518 = {_slots_34_io_uop_fu_code[5], _slots_34_io_uop_fu_code[0]};
  wire        _GEN_519 = _GEN_515 | _GEN_503;
  wire        _GEN_520 = _slots_34_io_request & (|(_slots_34_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_521 = _GEN_504 | _GEN_505;
  wire        _GEN_522 = _GEN_520 & ~_GEN_521;
  wire        _GEN_523 = _slots_34_io_request & (|_GEN_518) & ~_GEN_519 | _GEN_522;
  wire        _GEN_524 = _slots_34_io_request & ~(_slots_34_io_request & (|_can_allocate_T_138) & ~_GEN_517 | _GEN_523) & (|(_slots_34_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_525 = _GEN_508 | _GEN_511;
  wire        _GEN_526 = _GEN_524 & ~_GEN_525;
  wire        _GEN_527 = _slots_34_io_request & ~_GEN_523 & (|_can_allocate_T_138);
  wire        _GEN_528 = _GEN_527 & ~_GEN_517;
  wire        _GEN_529 = _slots_34_io_request & ~_GEN_522 & (|_GEN_518);
  wire        _GEN_530 = _GEN_529 & ~_GEN_519;
  wire        _GEN_23921 = _GEN_520 & ~_GEN_521;
  wire        issue_slots_34_grant = _GEN_526 | _GEN_528 | _GEN_530 | _GEN_23921;
  wire        _GEN_531 = _GEN_509 & ~_GEN_510;
  wire        _GEN_532 = _GEN_498 & ~_GEN_499;
  wire        _GEN_533 = _GEN_502 & ~_GEN_493;
  wire        _GEN_23273 = _GEN_494 & ~_GEN_495;
  wire        issue_slots_32_grant = _GEN_531 | _GEN_532 | _GEN_533 | _GEN_23273;
  wire [9:0]  _can_allocate_T_142 = _slots_35_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_534 = _GEN_527 | _GEN_517;
  wire [1:0]  _GEN_535 = {_slots_35_io_uop_fu_code[5], _slots_35_io_uop_fu_code[0]};
  wire        _GEN_536 = _GEN_529 | _GEN_519;
  wire        _GEN_537 = _slots_35_io_request & (|(_slots_35_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_538 = _GEN_520 | _GEN_521;
  wire        _GEN_539 = _GEN_537 & ~_GEN_538;
  wire        _GEN_540 = _slots_35_io_request & (|_GEN_535) & ~_GEN_536 | _GEN_539;
  wire        _GEN_541 = _slots_35_io_request & ~(_slots_35_io_request & (|_can_allocate_T_142) & ~_GEN_534 | _GEN_540) & (|(_slots_35_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_542 = _GEN_524 | _GEN_525;
  wire        _GEN_543 = _GEN_541 & ~_GEN_542;
  wire        _GEN_544 = _slots_35_io_request & ~_GEN_540 & (|_can_allocate_T_142);
  wire        _GEN_545 = _GEN_544 & ~_GEN_534;
  wire        _GEN_546 = _slots_35_io_request & ~_GEN_539 & (|_GEN_535);
  wire        _GEN_547 = _GEN_546 & ~_GEN_536;
  wire        _GEN_24245 = _GEN_537 & ~_GEN_538;
  wire        issue_slots_35_grant = _GEN_543 | _GEN_545 | _GEN_547 | _GEN_24245;
  wire [9:0]  _can_allocate_T_146 = _slots_36_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_548 = _GEN_544 | _GEN_534;
  wire [1:0]  _GEN_549 = {_slots_36_io_uop_fu_code[5], _slots_36_io_uop_fu_code[0]};
  wire        _GEN_550 = _GEN_546 | _GEN_536;
  wire        _GEN_551 = _slots_36_io_request & (|(_slots_36_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_552 = _GEN_537 | _GEN_538;
  wire        _GEN_553 = _GEN_551 & ~_GEN_552;
  wire        _GEN_554 = _slots_36_io_request & (|_GEN_549) & ~_GEN_550 | _GEN_553;
  wire        _GEN_555 = _slots_36_io_request & ~(_slots_36_io_request & (|_can_allocate_T_146) & ~_GEN_548 | _GEN_554) & (|(_slots_36_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_556 = _GEN_541 | _GEN_542;
  wire        _GEN_557 = _GEN_555 & ~_GEN_556;
  wire        _GEN_558 = _slots_36_io_request & ~_GEN_554 & (|_can_allocate_T_146);
  wire        _GEN_559 = _GEN_558 & ~_GEN_548;
  wire        _GEN_560 = _slots_36_io_request & ~_GEN_553 & (|_GEN_549);
  wire        _GEN_561 = _GEN_560 & ~_GEN_550;
  wire        _GEN_24569 = _GEN_551 & ~_GEN_552;
  wire        issue_slots_36_grant = _GEN_557 | _GEN_559 | _GEN_561 | _GEN_24569;
  wire [9:0]  _can_allocate_T_154 = _slots_38_io_uop_fu_code & io_fu_types_2;
  wire [1:0]  _GEN_562 = {_slots_37_io_uop_fu_code[5], _slots_37_io_uop_fu_code[0]};
  wire        _GEN_563 = _GEN_560 | _GEN_550;
  wire        _GEN_564 = _slots_37_io_request & (|(_slots_37_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_565 = _GEN_551 | _GEN_552;
  wire        _GEN_566 = _GEN_564 & ~_GEN_565;
  wire        _GEN_567 = _slots_37_io_request & (|_GEN_562) & ~_GEN_563 | _GEN_566;
  wire [9:0]  _can_allocate_T_150 = _slots_37_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_568 = _slots_37_io_request & ~_GEN_567 & (|_can_allocate_T_150);
  wire        _GEN_569 = _GEN_558 | _GEN_548;
  wire        _GEN_570 = _GEN_568 | _GEN_569;
  wire [1:0]  _GEN_571 = {_slots_38_io_uop_fu_code[5], _slots_38_io_uop_fu_code[0]};
  wire        _GEN_572 = _slots_37_io_request & ~_GEN_566 & (|_GEN_562);
  wire        _GEN_573 = _GEN_572 | _GEN_563;
  wire        _GEN_574 = _slots_38_io_request & (|(_slots_38_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_575 = _GEN_564 | _GEN_565;
  wire        _GEN_576 = _GEN_574 & ~_GEN_575;
  wire        _GEN_577 = _slots_38_io_request & (|_GEN_571) & ~_GEN_573 | _GEN_576;
  wire        _GEN_578 = _slots_38_io_request & ~(_slots_38_io_request & (|_can_allocate_T_154) & ~_GEN_570 | _GEN_577) & (|(_slots_38_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_579 = _slots_37_io_request & ~(_slots_37_io_request & (|_can_allocate_T_150) & ~_GEN_569 | _GEN_567) & (|(_slots_37_io_uop_fu_code & io_fu_types_3));
  wire        _GEN_580 = _GEN_555 | _GEN_556;
  wire        _GEN_581 = _GEN_579 | _GEN_580;
  wire        _GEN_582 = _GEN_578 & ~_GEN_581;
  wire        _GEN_583 = _slots_38_io_request & ~_GEN_577 & (|_can_allocate_T_154);
  wire        _GEN_584 = _GEN_583 & ~_GEN_570;
  wire        _GEN_585 = _slots_38_io_request & ~_GEN_576 & (|_GEN_571);
  wire        _GEN_586 = _GEN_585 & ~_GEN_573;
  wire        _GEN_25217 = _GEN_574 & ~_GEN_575;
  wire        issue_slots_38_grant = _GEN_582 | _GEN_584 | _GEN_586 | _GEN_25217;
  wire [9:0]  _can_allocate_T_158 = _slots_39_io_uop_fu_code & io_fu_types_2;
  wire        _GEN_587 = _GEN_583 | _GEN_570;
  wire [1:0]  _GEN_588 = {_slots_39_io_uop_fu_code[5], _slots_39_io_uop_fu_code[0]};
  wire        _GEN_589 = _GEN_585 | _GEN_573;
  wire        _GEN_590 = _slots_39_io_request & (|(_slots_39_io_uop_fu_code & io_fu_types_0));
  wire        _GEN_591 = _GEN_574 | _GEN_575;
  wire        _GEN_592 = _GEN_590 & ~_GEN_591;
  wire        _GEN_593 = _slots_39_io_request & (|_GEN_588) & ~_GEN_589 | _GEN_592;
  wire        _GEN_594 = _slots_39_io_request & ~(_slots_39_io_request & (|_can_allocate_T_158) & ~_GEN_587 | _GEN_593) & (|(_slots_39_io_uop_fu_code & io_fu_types_3)) & ~(_GEN_578 | _GEN_581);
  wire        _GEN_595 = _slots_39_io_request & ~_GEN_593 & (|_can_allocate_T_158) & ~_GEN_587;
  wire        _GEN_596 = _slots_39_io_request & ~_GEN_592 & (|_GEN_588) & ~_GEN_589;
  wire        _GEN_25541 = _GEN_590 & ~_GEN_591;
  wire        issue_slots_39_grant = _GEN_594 | _GEN_595 | _GEN_596 | _GEN_25541;
  wire        _GEN_597 = _GEN_579 & ~_GEN_580;
  wire        _GEN_598 = _GEN_568 & ~_GEN_569;
  wire        _GEN_599 = _GEN_572 & ~_GEN_563;
  wire        _GEN_24893 = _GEN_564 & ~_GEN_565;
  wire        issue_slots_37_grant = _GEN_597 | _GEN_598 | _GEN_599 | _GEN_24893;
  wire [3:0]  _GEN_23_0 = _slots_0_io_valid & ~_slots_1_io_valid ? 4'h1 : _slots_1_io_valid ? {3'h0, ~_slots_0_io_valid} : {2'h0, ~_slots_0_io_valid, 1'h0};
  assign _GEN_23_1to0 = _GEN_23_0[1:0];
  assign _GEN_25 = _GEN_23_1to0 == 2'h0 & ~_slots_2_io_valid ? 4'h1 : _GEN_23_0[3] | _slots_2_io_valid ? _GEN_23_0 : {_GEN_23_0[2:0], 1'h0};
  assign _GEN_27 = _GEN_25 == 4'h0 & ~_slots_3_io_valid ? 4'h1 : _GEN_25[3] | _slots_3_io_valid ? _GEN_25 : {_GEN_25[2:0], 1'h0};
  assign _GEN_29 = _GEN_27 == 4'h0 & ~_slots_4_io_valid ? 4'h1 : _GEN_27[3] | _slots_4_io_valid ? _GEN_27 : {_GEN_27[2:0], 1'h0};
  assign _GEN_31 = _GEN_29 == 4'h0 & ~_slots_5_io_valid ? 4'h1 : _GEN_29[3] | _slots_5_io_valid ? _GEN_29 : {_GEN_29[2:0], 1'h0};
  assign _GEN_33 = _GEN_31 == 4'h0 & ~_slots_6_io_valid ? 4'h1 : _GEN_31[3] | _slots_6_io_valid ? _GEN_31 : {_GEN_31[2:0], 1'h0};
  assign _GEN_35 = _GEN_33 == 4'h0 & ~_slots_7_io_valid ? 4'h1 : _GEN_33[3] | _slots_7_io_valid ? _GEN_33 : {_GEN_33[2:0], 1'h0};
  assign _GEN_37 = _GEN_35 == 4'h0 & ~_slots_8_io_valid ? 4'h1 : _GEN_35[3] | _slots_8_io_valid ? _GEN_35 : {_GEN_35[2:0], 1'h0};
  assign _GEN_39 = _GEN_37 == 4'h0 & ~_slots_9_io_valid ? 4'h1 : _GEN_37[3] | _slots_9_io_valid ? _GEN_37 : {_GEN_37[2:0], 1'h0};
  assign _GEN_41 = _GEN_39 == 4'h0 & ~_slots_10_io_valid ? 4'h1 : _GEN_39[3] | _slots_10_io_valid ? _GEN_39 : {_GEN_39[2:0], 1'h0};
  assign _GEN_43 = _GEN_41 == 4'h0 & ~_slots_11_io_valid ? 4'h1 : _GEN_41[3] | _slots_11_io_valid ? _GEN_41 : {_GEN_41[2:0], 1'h0};
  assign _GEN_45 = _GEN_43 == 4'h0 & ~_slots_12_io_valid ? 4'h1 : _GEN_43[3] | _slots_12_io_valid ? _GEN_43 : {_GEN_43[2:0], 1'h0};
  assign _GEN_47 = _GEN_45 == 4'h0 & ~_slots_13_io_valid ? 4'h1 : _GEN_45[3] | _slots_13_io_valid ? _GEN_45 : {_GEN_45[2:0], 1'h0};
  assign _GEN_49 = _GEN_47 == 4'h0 & ~_slots_14_io_valid ? 4'h1 : _GEN_47[3] | _slots_14_io_valid ? _GEN_47 : {_GEN_47[2:0], 1'h0};
  assign _GEN_51 = _GEN_49 == 4'h0 & ~_slots_15_io_valid ? 4'h1 : _GEN_49[3] | _slots_15_io_valid ? _GEN_49 : {_GEN_49[2:0], 1'h0};
  assign _GEN_53 = _GEN_51 == 4'h0 & ~_slots_16_io_valid ? 4'h1 : _GEN_51[3] | _slots_16_io_valid ? _GEN_51 : {_GEN_51[2:0], 1'h0};
  assign _GEN_55 = _GEN_53 == 4'h0 & ~_slots_17_io_valid ? 4'h1 : _GEN_53[3] | _slots_17_io_valid ? _GEN_53 : {_GEN_53[2:0], 1'h0};
  assign _GEN_57 = _GEN_55 == 4'h0 & ~_slots_18_io_valid ? 4'h1 : _GEN_55[3] | _slots_18_io_valid ? _GEN_55 : {_GEN_55[2:0], 1'h0};
  assign _GEN_59 = _GEN_57 == 4'h0 & ~_slots_19_io_valid ? 4'h1 : _GEN_57[3] | _slots_19_io_valid ? _GEN_57 : {_GEN_57[2:0], 1'h0};
  assign _GEN_61 = _GEN_59 == 4'h0 & ~_slots_20_io_valid ? 4'h1 : _GEN_59[3] | _slots_20_io_valid ? _GEN_59 : {_GEN_59[2:0], 1'h0};
  assign _GEN_63 = _GEN_61 == 4'h0 & ~_slots_21_io_valid ? 4'h1 : _GEN_61[3] | _slots_21_io_valid ? _GEN_61 : {_GEN_61[2:0], 1'h0};
  assign _GEN_65 = _GEN_63 == 4'h0 & ~_slots_22_io_valid ? 4'h1 : _GEN_63[3] | _slots_22_io_valid ? _GEN_63 : {_GEN_63[2:0], 1'h0};
  assign _GEN_67 = _GEN_65 == 4'h0 & ~_slots_23_io_valid ? 4'h1 : _GEN_65[3] | _slots_23_io_valid ? _GEN_65 : {_GEN_65[2:0], 1'h0};
  assign _GEN_69 = _GEN_67 == 4'h0 & ~_slots_24_io_valid ? 4'h1 : _GEN_67[3] | _slots_24_io_valid ? _GEN_67 : {_GEN_67[2:0], 1'h0};
  assign _GEN_71 = _GEN_69 == 4'h0 & ~_slots_25_io_valid ? 4'h1 : _GEN_69[3] | _slots_25_io_valid ? _GEN_69 : {_GEN_69[2:0], 1'h0};
  assign _GEN_73 = _GEN_71 == 4'h0 & ~_slots_26_io_valid ? 4'h1 : _GEN_71[3] | _slots_26_io_valid ? _GEN_71 : {_GEN_71[2:0], 1'h0};
  assign _GEN_75 = _GEN_73 == 4'h0 & ~_slots_27_io_valid ? 4'h1 : _GEN_73[3] | _slots_27_io_valid ? _GEN_73 : {_GEN_73[2:0], 1'h0};
  assign _GEN_77 = _GEN_75 == 4'h0 & ~_slots_28_io_valid ? 4'h1 : _GEN_75[3] | _slots_28_io_valid ? _GEN_75 : {_GEN_75[2:0], 1'h0};
  assign _GEN_79 = _GEN_77 == 4'h0 & ~_slots_29_io_valid ? 4'h1 : _GEN_77[3] | _slots_29_io_valid ? _GEN_77 : {_GEN_77[2:0], 1'h0};
  assign _GEN_81 = _GEN_79 == 4'h0 & ~_slots_30_io_valid ? 4'h1 : _GEN_79[3] | _slots_30_io_valid ? _GEN_79 : {_GEN_79[2:0], 1'h0};
  assign _GEN_83 = _GEN_81 == 4'h0 & ~_slots_31_io_valid ? 4'h1 : _GEN_81[3] | _slots_31_io_valid ? _GEN_81 : {_GEN_81[2:0], 1'h0};
  assign _GEN_85 = _GEN_83 == 4'h0 & ~_slots_32_io_valid ? 4'h1 : _GEN_83[3] | _slots_32_io_valid ? _GEN_83 : {_GEN_83[2:0], 1'h0};
  assign _GEN_87 = _GEN_85 == 4'h0 & ~_slots_33_io_valid ? 4'h1 : _GEN_85[3] | _slots_33_io_valid ? _GEN_85 : {_GEN_85[2:0], 1'h0};
  assign _GEN_89 = _GEN_87 == 4'h0 & ~_slots_34_io_valid ? 4'h1 : _GEN_87[3] | _slots_34_io_valid ? _GEN_87 : {_GEN_87[2:0], 1'h0};
  assign _GEN_91 = _GEN_89 == 4'h0 & ~_slots_35_io_valid ? 4'h1 : _GEN_89[3] | _slots_35_io_valid ? _GEN_89 : {_GEN_89[2:0], 1'h0};
  assign _GEN_93 = _GEN_91 == 4'h0 & ~_slots_36_io_valid ? 4'h1 : _GEN_91[3] | _slots_36_io_valid ? _GEN_91 : {_GEN_91[2:0], 1'h0};
  assign _GEN_95 = _GEN_93 == 4'h0 & ~_slots_37_io_valid ? 4'h1 : _GEN_93[3] | _slots_37_io_valid ? _GEN_93 : {_GEN_93[2:0], 1'h0};
  assign _GEN_97 = _GEN_95 == 4'h0 & ~_slots_38_io_valid ? 4'h1 : _GEN_95[3] | _slots_38_io_valid ? _GEN_95 : {_GEN_95[2:0], 1'h0};
  wire [3:0]  _GEN_99_0 = _GEN_97 == 4'h0 & ~_slots_39_io_valid ? 4'h1 : _GEN_97[3] | _slots_39_io_valid ? _GEN_97 : {_GEN_97[2:0], 1'h0};
  wire [3:0]  _GEN_101_0 = _GEN_99_0 == 4'h0 & ~io_dis_uops_0_valid ? 4'h1 : _GEN_99_0[3] | io_dis_uops_0_valid ? _GEN_99_0 : {_GEN_99_0[2:0], 1'h0};
  wire [3:0]  _GEN_103_0 = _GEN_101_0 == 4'h0 & ~io_dis_uops_1_valid ? 4'h1 : _GEN_101_0[3] | io_dis_uops_1_valid ? _GEN_101_0 : {_GEN_101_0[2:0], 1'h0};
  wire        will_be_valid_40 = io_dis_uops_0_valid & ~io_dis_uops_0_bits_exception & ~io_dis_uops_0_bits_is_fence & ~io_dis_uops_0_bits_is_fencei;
  wire        will_be_valid_41 = io_dis_uops_1_valid & ~io_dis_uops_1_bits_exception & ~io_dis_uops_1_bits_is_fence & ~io_dis_uops_1_bits_is_fencei;
  wire        will_be_valid_42 = io_dis_uops_2_valid & ~io_dis_uops_2_bits_exception & ~io_dis_uops_2_bits_is_fence & ~io_dis_uops_2_bits_is_fencei;
  wire        _GEN_600 = _GEN_23_1to0 == 2'h2;
  wire        _GEN_601 = _GEN_25 == 4'h4;
  wire        _GEN_602 = _GEN_27 == 4'h8;
  wire        issue_slots_0_in_uop_valid = _GEN_602 ? _slots_4_io_will_be_valid : _GEN_601 ? _slots_3_io_will_be_valid : _GEN_600 ? _slots_2_io_will_be_valid : ~_slots_0_io_valid & _slots_1_io_will_be_valid;
  wire        _GEN_603 = _GEN_25 == 4'h2;
  wire        _GEN_604 = _GEN_27 == 4'h4;
  wire        _GEN_605 = _GEN_29 == 4'h8;
  wire        issue_slots_1_in_uop_valid = _GEN_605 ? _slots_5_io_will_be_valid : _GEN_604 ? _slots_4_io_will_be_valid : _GEN_603 ? _slots_3_io_will_be_valid : _GEN_23_1to0 == 2'h1 & _slots_2_io_will_be_valid;
  wire        _GEN_606 = _GEN_27 == 4'h2;
  wire        _GEN_607 = _GEN_29 == 4'h4;
  wire        _GEN_608 = _GEN_31 == 4'h8;
  wire        issue_slots_2_in_uop_valid = _GEN_608 ? _slots_6_io_will_be_valid : _GEN_607 ? _slots_5_io_will_be_valid : _GEN_606 ? _slots_4_io_will_be_valid : _GEN_25 == 4'h1 & _slots_3_io_will_be_valid;
  wire        _GEN_609 = _GEN_29 == 4'h2;
  wire        _GEN_610 = _GEN_31 == 4'h4;
  wire        _GEN_611 = _GEN_33 == 4'h8;
  wire        issue_slots_3_in_uop_valid = _GEN_611 ? _slots_7_io_will_be_valid : _GEN_610 ? _slots_6_io_will_be_valid : _GEN_609 ? _slots_5_io_will_be_valid : _GEN_27 == 4'h1 & _slots_4_io_will_be_valid;
  wire        _GEN_612 = _GEN_31 == 4'h2;
  wire        _GEN_613 = _GEN_33 == 4'h4;
  wire        _GEN_614 = _GEN_35 == 4'h8;
  wire        issue_slots_4_in_uop_valid = _GEN_614 ? _slots_8_io_will_be_valid : _GEN_613 ? _slots_7_io_will_be_valid : _GEN_612 ? _slots_6_io_will_be_valid : _GEN_29 == 4'h1 & _slots_5_io_will_be_valid;
  wire        _GEN_615 = _GEN_33 == 4'h2;
  wire        _GEN_616 = _GEN_35 == 4'h4;
  wire        _GEN_617 = _GEN_37 == 4'h8;
  wire        issue_slots_5_in_uop_valid = _GEN_617 ? _slots_9_io_will_be_valid : _GEN_616 ? _slots_8_io_will_be_valid : _GEN_615 ? _slots_7_io_will_be_valid : _GEN_31 == 4'h1 & _slots_6_io_will_be_valid;
  wire        _GEN_618 = _GEN_35 == 4'h2;
  wire        _GEN_619 = _GEN_37 == 4'h4;
  wire        _GEN_620 = _GEN_39 == 4'h8;
  wire        issue_slots_6_in_uop_valid = _GEN_620 ? _slots_10_io_will_be_valid : _GEN_619 ? _slots_9_io_will_be_valid : _GEN_618 ? _slots_8_io_will_be_valid : _GEN_33 == 4'h1 & _slots_7_io_will_be_valid;
  wire        _GEN_621 = _GEN_37 == 4'h2;
  wire        _GEN_622 = _GEN_39 == 4'h4;
  wire        _GEN_623 = _GEN_41 == 4'h8;
  wire        issue_slots_7_in_uop_valid = _GEN_623 ? _slots_11_io_will_be_valid : _GEN_622 ? _slots_10_io_will_be_valid : _GEN_621 ? _slots_9_io_will_be_valid : _GEN_35 == 4'h1 & _slots_8_io_will_be_valid;
  wire        _GEN_624 = _GEN_39 == 4'h2;
  wire        _GEN_625 = _GEN_41 == 4'h4;
  wire        _GEN_626 = _GEN_43 == 4'h8;
  wire        issue_slots_8_in_uop_valid = _GEN_626 ? _slots_12_io_will_be_valid : _GEN_625 ? _slots_11_io_will_be_valid : _GEN_624 ? _slots_10_io_will_be_valid : _GEN_37 == 4'h1 & _slots_9_io_will_be_valid;
  wire        _GEN_627 = _GEN_41 == 4'h2;
  wire        _GEN_628 = _GEN_43 == 4'h4;
  wire        _GEN_629 = _GEN_45 == 4'h8;
  wire        issue_slots_9_in_uop_valid = _GEN_629 ? _slots_13_io_will_be_valid : _GEN_628 ? _slots_12_io_will_be_valid : _GEN_627 ? _slots_11_io_will_be_valid : _GEN_39 == 4'h1 & _slots_10_io_will_be_valid;
  wire        _GEN_630 = _GEN_43 == 4'h2;
  wire        _GEN_631 = _GEN_45 == 4'h4;
  wire        _GEN_632 = _GEN_47 == 4'h8;
  wire        issue_slots_10_in_uop_valid = _GEN_632 ? _slots_14_io_will_be_valid : _GEN_631 ? _slots_13_io_will_be_valid : _GEN_630 ? _slots_12_io_will_be_valid : _GEN_41 == 4'h1 & _slots_11_io_will_be_valid;
  wire        _GEN_633 = _GEN_45 == 4'h2;
  wire        _GEN_634 = _GEN_47 == 4'h4;
  wire        _GEN_635 = _GEN_49 == 4'h8;
  wire        issue_slots_11_in_uop_valid = _GEN_635 ? _slots_15_io_will_be_valid : _GEN_634 ? _slots_14_io_will_be_valid : _GEN_633 ? _slots_13_io_will_be_valid : _GEN_43 == 4'h1 & _slots_12_io_will_be_valid;
  wire        _GEN_636 = _GEN_47 == 4'h2;
  wire        _GEN_637 = _GEN_49 == 4'h4;
  wire        _GEN_638 = _GEN_51 == 4'h8;
  wire        issue_slots_12_in_uop_valid = _GEN_638 ? _slots_16_io_will_be_valid : _GEN_637 ? _slots_15_io_will_be_valid : _GEN_636 ? _slots_14_io_will_be_valid : _GEN_45 == 4'h1 & _slots_13_io_will_be_valid;
  wire        _GEN_639 = _GEN_49 == 4'h2;
  wire        _GEN_640 = _GEN_51 == 4'h4;
  wire        _GEN_641 = _GEN_53 == 4'h8;
  wire        issue_slots_13_in_uop_valid = _GEN_641 ? _slots_17_io_will_be_valid : _GEN_640 ? _slots_16_io_will_be_valid : _GEN_639 ? _slots_15_io_will_be_valid : _GEN_47 == 4'h1 & _slots_14_io_will_be_valid;
  wire        _GEN_642 = _GEN_51 == 4'h2;
  wire        _GEN_643 = _GEN_53 == 4'h4;
  wire        _GEN_644 = _GEN_55 == 4'h8;
  wire        issue_slots_14_in_uop_valid = _GEN_644 ? _slots_18_io_will_be_valid : _GEN_643 ? _slots_17_io_will_be_valid : _GEN_642 ? _slots_16_io_will_be_valid : _GEN_49 == 4'h1 & _slots_15_io_will_be_valid;
  wire        _GEN_645 = _GEN_53 == 4'h2;
  wire        _GEN_646 = _GEN_55 == 4'h4;
  wire        _GEN_647 = _GEN_57 == 4'h8;
  wire        issue_slots_15_in_uop_valid = _GEN_647 ? _slots_19_io_will_be_valid : _GEN_646 ? _slots_18_io_will_be_valid : _GEN_645 ? _slots_17_io_will_be_valid : _GEN_51 == 4'h1 & _slots_16_io_will_be_valid;
  wire        _GEN_648 = _GEN_55 == 4'h2;
  wire        _GEN_649 = _GEN_57 == 4'h4;
  wire        _GEN_650 = _GEN_59 == 4'h8;
  wire        issue_slots_16_in_uop_valid = _GEN_650 ? _slots_20_io_will_be_valid : _GEN_649 ? _slots_19_io_will_be_valid : _GEN_648 ? _slots_18_io_will_be_valid : _GEN_53 == 4'h1 & _slots_17_io_will_be_valid;
  wire        _GEN_651 = _GEN_57 == 4'h2;
  wire        _GEN_652 = _GEN_59 == 4'h4;
  wire        _GEN_653 = _GEN_61 == 4'h8;
  wire        issue_slots_17_in_uop_valid = _GEN_653 ? _slots_21_io_will_be_valid : _GEN_652 ? _slots_20_io_will_be_valid : _GEN_651 ? _slots_19_io_will_be_valid : _GEN_55 == 4'h1 & _slots_18_io_will_be_valid;
  wire        _GEN_654 = _GEN_59 == 4'h2;
  wire        _GEN_655 = _GEN_61 == 4'h4;
  wire        _GEN_656 = _GEN_63 == 4'h8;
  wire        issue_slots_18_in_uop_valid = _GEN_656 ? _slots_22_io_will_be_valid : _GEN_655 ? _slots_21_io_will_be_valid : _GEN_654 ? _slots_20_io_will_be_valid : _GEN_57 == 4'h1 & _slots_19_io_will_be_valid;
  wire        _GEN_657 = _GEN_61 == 4'h2;
  wire        _GEN_658 = _GEN_63 == 4'h4;
  wire        _GEN_659 = _GEN_65 == 4'h8;
  wire        issue_slots_19_in_uop_valid = _GEN_659 ? _slots_23_io_will_be_valid : _GEN_658 ? _slots_22_io_will_be_valid : _GEN_657 ? _slots_21_io_will_be_valid : _GEN_59 == 4'h1 & _slots_20_io_will_be_valid;
  wire        _GEN_660 = _GEN_63 == 4'h2;
  wire        _GEN_661 = _GEN_65 == 4'h4;
  wire        _GEN_662 = _GEN_67 == 4'h8;
  wire        issue_slots_20_in_uop_valid = _GEN_662 ? _slots_24_io_will_be_valid : _GEN_661 ? _slots_23_io_will_be_valid : _GEN_660 ? _slots_22_io_will_be_valid : _GEN_61 == 4'h1 & _slots_21_io_will_be_valid;
  wire        _GEN_663 = _GEN_65 == 4'h2;
  wire        _GEN_664 = _GEN_67 == 4'h4;
  wire        _GEN_665 = _GEN_69 == 4'h8;
  wire        issue_slots_21_in_uop_valid = _GEN_665 ? _slots_25_io_will_be_valid : _GEN_664 ? _slots_24_io_will_be_valid : _GEN_663 ? _slots_23_io_will_be_valid : _GEN_63 == 4'h1 & _slots_22_io_will_be_valid;
  wire        _GEN_666 = _GEN_67 == 4'h2;
  wire        _GEN_667 = _GEN_69 == 4'h4;
  wire        _GEN_668 = _GEN_71 == 4'h8;
  wire        issue_slots_22_in_uop_valid = _GEN_668 ? _slots_26_io_will_be_valid : _GEN_667 ? _slots_25_io_will_be_valid : _GEN_666 ? _slots_24_io_will_be_valid : _GEN_65 == 4'h1 & _slots_23_io_will_be_valid;
  wire        _GEN_669 = _GEN_69 == 4'h2;
  wire        _GEN_670 = _GEN_71 == 4'h4;
  wire        _GEN_671 = _GEN_73 == 4'h8;
  wire        issue_slots_23_in_uop_valid = _GEN_671 ? _slots_27_io_will_be_valid : _GEN_670 ? _slots_26_io_will_be_valid : _GEN_669 ? _slots_25_io_will_be_valid : _GEN_67 == 4'h1 & _slots_24_io_will_be_valid;
  wire        _GEN_672 = _GEN_71 == 4'h2;
  wire        _GEN_673 = _GEN_73 == 4'h4;
  wire        _GEN_674 = _GEN_75 == 4'h8;
  wire        issue_slots_24_in_uop_valid = _GEN_674 ? _slots_28_io_will_be_valid : _GEN_673 ? _slots_27_io_will_be_valid : _GEN_672 ? _slots_26_io_will_be_valid : _GEN_69 == 4'h1 & _slots_25_io_will_be_valid;
  wire        _GEN_675 = _GEN_73 == 4'h2;
  wire        _GEN_676 = _GEN_75 == 4'h4;
  wire        _GEN_677 = _GEN_77 == 4'h8;
  wire        issue_slots_25_in_uop_valid = _GEN_677 ? _slots_29_io_will_be_valid : _GEN_676 ? _slots_28_io_will_be_valid : _GEN_675 ? _slots_27_io_will_be_valid : _GEN_71 == 4'h1 & _slots_26_io_will_be_valid;
  wire        _GEN_678 = _GEN_75 == 4'h2;
  wire        _GEN_679 = _GEN_77 == 4'h4;
  wire        _GEN_680 = _GEN_79 == 4'h8;
  wire        issue_slots_26_in_uop_valid = _GEN_680 ? _slots_30_io_will_be_valid : _GEN_679 ? _slots_29_io_will_be_valid : _GEN_678 ? _slots_28_io_will_be_valid : _GEN_73 == 4'h1 & _slots_27_io_will_be_valid;
  wire        _GEN_681 = _GEN_77 == 4'h2;
  wire        _GEN_682 = _GEN_79 == 4'h4;
  wire        _GEN_683 = _GEN_81 == 4'h8;
  wire        issue_slots_27_in_uop_valid = _GEN_683 ? _slots_31_io_will_be_valid : _GEN_682 ? _slots_30_io_will_be_valid : _GEN_681 ? _slots_29_io_will_be_valid : _GEN_75 == 4'h1 & _slots_28_io_will_be_valid;
  wire        _GEN_684 = _GEN_79 == 4'h2;
  wire        _GEN_685 = _GEN_81 == 4'h4;
  wire        _GEN_686 = _GEN_83 == 4'h8;
  wire        issue_slots_28_in_uop_valid = _GEN_686 ? _slots_32_io_will_be_valid : _GEN_685 ? _slots_31_io_will_be_valid : _GEN_684 ? _slots_30_io_will_be_valid : _GEN_77 == 4'h1 & _slots_29_io_will_be_valid;
  wire        _GEN_687 = _GEN_81 == 4'h2;
  wire        _GEN_688 = _GEN_83 == 4'h4;
  wire        _GEN_689 = _GEN_85 == 4'h8;
  wire        issue_slots_29_in_uop_valid = _GEN_689 ? _slots_33_io_will_be_valid : _GEN_688 ? _slots_32_io_will_be_valid : _GEN_687 ? _slots_31_io_will_be_valid : _GEN_79 == 4'h1 & _slots_30_io_will_be_valid;
  wire        _GEN_690 = _GEN_83 == 4'h2;
  wire        _GEN_691 = _GEN_85 == 4'h4;
  wire        _GEN_692 = _GEN_87 == 4'h8;
  wire        issue_slots_30_in_uop_valid = _GEN_692 ? _slots_34_io_will_be_valid : _GEN_691 ? _slots_33_io_will_be_valid : _GEN_690 ? _slots_32_io_will_be_valid : _GEN_81 == 4'h1 & _slots_31_io_will_be_valid;
  wire        _GEN_693 = _GEN_85 == 4'h2;
  wire        _GEN_694 = _GEN_87 == 4'h4;
  wire        _GEN_695 = _GEN_89 == 4'h8;
  wire        issue_slots_31_in_uop_valid = _GEN_695 ? _slots_35_io_will_be_valid : _GEN_694 ? _slots_34_io_will_be_valid : _GEN_693 ? _slots_33_io_will_be_valid : _GEN_83 == 4'h1 & _slots_32_io_will_be_valid;
  wire        _GEN_696 = _GEN_87 == 4'h2;
  wire        _GEN_697 = _GEN_89 == 4'h4;
  wire        _GEN_698 = _GEN_91 == 4'h8;
  wire        issue_slots_32_in_uop_valid = _GEN_698 ? _slots_36_io_will_be_valid : _GEN_697 ? _slots_35_io_will_be_valid : _GEN_696 ? _slots_34_io_will_be_valid : _GEN_85 == 4'h1 & _slots_33_io_will_be_valid;
  wire        _GEN_699 = _GEN_89 == 4'h2;
  wire        _GEN_700 = _GEN_91 == 4'h4;
  wire        _GEN_701 = _GEN_93 == 4'h8;
  wire        issue_slots_33_in_uop_valid = _GEN_701 ? _slots_37_io_will_be_valid : _GEN_700 ? _slots_36_io_will_be_valid : _GEN_699 ? _slots_35_io_will_be_valid : _GEN_87 == 4'h1 & _slots_34_io_will_be_valid;
  wire        _GEN_702 = _GEN_91 == 4'h2;
  wire        _GEN_703 = _GEN_93 == 4'h4;
  wire        _GEN_704 = _GEN_95 == 4'h8;
  wire        issue_slots_34_in_uop_valid = _GEN_704 ? _slots_38_io_will_be_valid : _GEN_703 ? _slots_37_io_will_be_valid : _GEN_702 ? _slots_36_io_will_be_valid : _GEN_89 == 4'h1 & _slots_35_io_will_be_valid;
  wire        _GEN_705 = _GEN_93 == 4'h2;
  wire        _GEN_706 = _GEN_95 == 4'h4;
  wire        _GEN_707 = _GEN_97 == 4'h8;
  wire        issue_slots_35_in_uop_valid = _GEN_707 ? _slots_39_io_will_be_valid : _GEN_706 ? _slots_38_io_will_be_valid : _GEN_705 ? _slots_37_io_will_be_valid : _GEN_91 == 4'h1 & _slots_36_io_will_be_valid;
  wire        _GEN_708 = _GEN_95 == 4'h2;
  wire        _GEN_709 = _GEN_97 == 4'h4;
  wire        _GEN_710 = _GEN_99_0 == 4'h8;
  wire        issue_slots_36_in_uop_valid = _GEN_710 ? will_be_valid_40 : _GEN_709 ? _slots_39_io_will_be_valid : _GEN_708 ? _slots_38_io_will_be_valid : _GEN_93 == 4'h1 & _slots_37_io_will_be_valid;
  wire        _GEN_711 = _GEN_97 == 4'h2;
  wire        _GEN_712 = _GEN_99_0 == 4'h4;
  wire        _GEN_713 = _GEN_101_0 == 4'h8;
  wire        issue_slots_37_in_uop_valid = _GEN_713 ? will_be_valid_41 : _GEN_712 ? will_be_valid_40 : _GEN_711 ? _slots_39_io_will_be_valid : _GEN_95 == 4'h1 & _slots_38_io_will_be_valid;
  wire        _GEN_714 = _GEN_713 | _GEN_712;
  wire        _GEN_715 = _GEN_99_0 == 4'h2;
  wire        _GEN_716 = _GEN_101_0 == 4'h4;
  wire        _GEN_717 = _GEN_103_0 == 4'h8;
  wire        issue_slots_38_in_uop_valid = _GEN_717 ? will_be_valid_42 : _GEN_716 ? will_be_valid_41 : _GEN_715 ? will_be_valid_40 : _GEN_97 == 4'h1 & _slots_39_io_will_be_valid;
  wire        _GEN_718 = _GEN_717 | _GEN_716 | _GEN_715;
  wire        _GEN_719 = _GEN_101_0 == 4'h2;
  wire        _GEN_720 = _GEN_103_0 == 4'h4;
  wire        _GEN_721 = (_GEN_103_0 == 4'h0 & ~io_dis_uops_2_valid ? 4'h1 : _GEN_103_0[3] | io_dis_uops_2_valid ? _GEN_103_0 : {_GEN_103_0[2:0], 1'h0}) == 4'h8;
  wire        issue_slots_39_in_uop_valid = _GEN_721 ? io_dis_uops_3_valid & ~io_dis_uops_3_bits_exception & ~io_dis_uops_3_bits_is_fence & ~io_dis_uops_3_bits_is_fencei : _GEN_720 ? will_be_valid_42 : _GEN_719 ? will_be_valid_41 : _GEN_99_0 == 4'h1 & will_be_valid_40;
  reg         io_dis_uops_0_ready_REG;
  reg         io_dis_uops_1_ready_REG;
  reg         io_dis_uops_2_ready_REG;
  reg         io_dis_uops_3_ready_REG;
  wire [5:0]  num_available =
    {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, ~_slots_0_io_will_be_valid & ~issue_slots_0_in_uop_valid} + {1'h0, (~_slots_1_io_will_be_valid | ~_slots_0_io_valid) & ~issue_slots_1_in_uop_valid}} + {1'h0, {1'h0, (~_slots_2_io_will_be_valid | (|_GEN_23_1to0)) & ~issue_slots_2_in_uop_valid} + {1'h0, (~_slots_3_io_will_be_valid | (|_GEN_25)) & ~issue_slots_3_in_uop_valid} + {1'h0, (~_slots_4_io_will_be_valid | (|_GEN_27)) & ~issue_slots_4_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_5_io_will_be_valid | (|_GEN_29)) & ~issue_slots_5_in_uop_valid} + {1'h0, (~_slots_6_io_will_be_valid | (|_GEN_31)) & ~issue_slots_6_in_uop_valid}} + {1'h0, {1'h0, (~_slots_7_io_will_be_valid | (|_GEN_33)) & ~issue_slots_7_in_uop_valid} + {1'h0, (~_slots_8_io_will_be_valid | (|_GEN_35)) & ~issue_slots_8_in_uop_valid} + {1'h0, (~_slots_9_io_will_be_valid | (|_GEN_37)) & ~issue_slots_9_in_uop_valid}}}} + {1'h0, {1'h0, {1'h0, {1'h0, (~_slots_10_io_will_be_valid | (|_GEN_39)) & ~issue_slots_10_in_uop_valid} + {1'h0, (~_slots_11_io_will_be_valid | (|_GEN_41)) & ~issue_slots_11_in_uop_valid}} + {1'h0, {1'h0, (~_slots_12_io_will_be_valid | (|_GEN_43)) & ~issue_slots_12_in_uop_valid} + {1'h0, (~_slots_13_io_will_be_valid | (|_GEN_45)) & ~issue_slots_13_in_uop_valid} + {1'h0, (~_slots_14_io_will_be_valid | (|_GEN_47)) & ~issue_slots_14_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_15_io_will_be_valid | (|_GEN_49)) & ~issue_slots_15_in_uop_valid} + {1'h0, (~_slots_16_io_will_be_valid | (|_GEN_51)) & ~issue_slots_16_in_uop_valid}} + {1'h0, {1'h0, (~_slots_17_io_will_be_valid | (|_GEN_53)) & ~issue_slots_17_in_uop_valid} + {1'h0, (~_slots_18_io_will_be_valid | (|_GEN_55)) & ~issue_slots_18_in_uop_valid} + {1'h0, (~_slots_19_io_will_be_valid | (|_GEN_57)) & ~issue_slots_19_in_uop_valid}}}}}
    + {1'h0, {1'h0, {1'h0, {1'h0, {1'h0, (~_slots_20_io_will_be_valid | (|_GEN_59)) & ~issue_slots_20_in_uop_valid} + {1'h0, (~_slots_21_io_will_be_valid | (|_GEN_61)) & ~issue_slots_21_in_uop_valid}} + {1'h0, {1'h0, (~_slots_22_io_will_be_valid | (|_GEN_63)) & ~issue_slots_22_in_uop_valid} + {1'h0, (~_slots_23_io_will_be_valid | (|_GEN_65)) & ~issue_slots_23_in_uop_valid} + {1'h0, (~_slots_24_io_will_be_valid | (|_GEN_67)) & ~issue_slots_24_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_25_io_will_be_valid | (|_GEN_69)) & ~issue_slots_25_in_uop_valid} + {1'h0, (~_slots_26_io_will_be_valid | (|_GEN_71)) & ~issue_slots_26_in_uop_valid}} + {1'h0, {1'h0, (~_slots_27_io_will_be_valid | (|_GEN_73)) & ~issue_slots_27_in_uop_valid} + {1'h0, (~_slots_28_io_will_be_valid | (|_GEN_75)) & ~issue_slots_28_in_uop_valid} + {1'h0, (~_slots_29_io_will_be_valid | (|_GEN_77)) & ~issue_slots_29_in_uop_valid}}}} + {1'h0, {1'h0, {1'h0, {1'h0, (~_slots_30_io_will_be_valid | (|_GEN_79)) & ~issue_slots_30_in_uop_valid} + {1'h0, (~_slots_31_io_will_be_valid | (|_GEN_81)) & ~issue_slots_31_in_uop_valid}} + {1'h0, {1'h0, (~_slots_32_io_will_be_valid | (|_GEN_83)) & ~issue_slots_32_in_uop_valid} + {1'h0, (~_slots_33_io_will_be_valid | (|_GEN_85)) & ~issue_slots_33_in_uop_valid} + {1'h0, (~_slots_34_io_will_be_valid | (|_GEN_87)) & ~issue_slots_34_in_uop_valid}}} + {1'h0, {1'h0, {1'h0, (~_slots_35_io_will_be_valid | (|_GEN_89)) & ~issue_slots_35_in_uop_valid} + {1'h0, (~_slots_36_io_will_be_valid | (|_GEN_91)) & ~issue_slots_36_in_uop_valid}} + {1'h0, {1'h0, (~_slots_37_io_will_be_valid | (|_GEN_93)) & ~issue_slots_37_in_uop_valid} + {1'h0, (~_slots_38_io_will_be_valid | (|_GEN_95)) & ~issue_slots_38_in_uop_valid} + {1'h0, (~_slots_39_io_will_be_valid | (|_GEN_97)) & ~issue_slots_39_in_uop_valid}}}}};
  always @(posedge clock) begin
    io_dis_uops_0_ready_REG <= |num_available;
    io_dis_uops_1_ready_REG <= |(num_available[5:1]);
    io_dis_uops_2_ready_REG <= num_available > 6'h2;
    io_dis_uops_3_ready_REG <= |(num_available[5:2]);
  end // always @(posedge)
  IssueSlot_32 slots_0 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_0_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (1'h0),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_0_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_602 ? _slots_4_io_out_uop_uopc : _GEN_601 ? _slots_3_io_out_uop_uopc : _GEN_600 ? _slots_2_io_out_uop_uopc : _slots_1_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_602 ? _slots_4_io_out_uop_is_rvc : _GEN_601 ? _slots_3_io_out_uop_is_rvc : _GEN_600 ? _slots_2_io_out_uop_is_rvc : _slots_1_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_602 ? _slots_4_io_out_uop_fu_code : _GEN_601 ? _slots_3_io_out_uop_fu_code : _GEN_600 ? _slots_2_io_out_uop_fu_code : _slots_1_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_602 ? _slots_4_io_out_uop_iw_state : _GEN_601 ? _slots_3_io_out_uop_iw_state : _GEN_600 ? _slots_2_io_out_uop_iw_state : _slots_1_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_602 ? _slots_4_io_out_uop_iw_p1_poisoned : _GEN_601 ? _slots_3_io_out_uop_iw_p1_poisoned : _GEN_600 ? _slots_2_io_out_uop_iw_p1_poisoned : _slots_1_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_602 ? _slots_4_io_out_uop_iw_p2_poisoned : _GEN_601 ? _slots_3_io_out_uop_iw_p2_poisoned : _GEN_600 ? _slots_2_io_out_uop_iw_p2_poisoned : _slots_1_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_602 ? _slots_4_io_out_uop_is_br : _GEN_601 ? _slots_3_io_out_uop_is_br : _GEN_600 ? _slots_2_io_out_uop_is_br : _slots_1_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_602 ? _slots_4_io_out_uop_is_jalr : _GEN_601 ? _slots_3_io_out_uop_is_jalr : _GEN_600 ? _slots_2_io_out_uop_is_jalr : _slots_1_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_602 ? _slots_4_io_out_uop_is_jal : _GEN_601 ? _slots_3_io_out_uop_is_jal : _GEN_600 ? _slots_2_io_out_uop_is_jal : _slots_1_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_602 ? _slots_4_io_out_uop_is_sfb : _GEN_601 ? _slots_3_io_out_uop_is_sfb : _GEN_600 ? _slots_2_io_out_uop_is_sfb : _slots_1_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_602 ? _slots_4_io_out_uop_br_mask : _GEN_601 ? _slots_3_io_out_uop_br_mask : _GEN_600 ? _slots_2_io_out_uop_br_mask : _slots_1_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_602 ? _slots_4_io_out_uop_br_tag : _GEN_601 ? _slots_3_io_out_uop_br_tag : _GEN_600 ? _slots_2_io_out_uop_br_tag : _slots_1_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_602 ? _slots_4_io_out_uop_ftq_idx : _GEN_601 ? _slots_3_io_out_uop_ftq_idx : _GEN_600 ? _slots_2_io_out_uop_ftq_idx : _slots_1_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_602 ? _slots_4_io_out_uop_edge_inst : _GEN_601 ? _slots_3_io_out_uop_edge_inst : _GEN_600 ? _slots_2_io_out_uop_edge_inst : _slots_1_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_602 ? _slots_4_io_out_uop_pc_lob : _GEN_601 ? _slots_3_io_out_uop_pc_lob : _GEN_600 ? _slots_2_io_out_uop_pc_lob : _slots_1_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_602 ? _slots_4_io_out_uop_taken : _GEN_601 ? _slots_3_io_out_uop_taken : _GEN_600 ? _slots_2_io_out_uop_taken : _slots_1_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_602 ? _slots_4_io_out_uop_imm_packed : _GEN_601 ? _slots_3_io_out_uop_imm_packed : _GEN_600 ? _slots_2_io_out_uop_imm_packed : _slots_1_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_602 ? _slots_4_io_out_uop_rob_idx : _GEN_601 ? _slots_3_io_out_uop_rob_idx : _GEN_600 ? _slots_2_io_out_uop_rob_idx : _slots_1_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_602 ? _slots_4_io_out_uop_ldq_idx : _GEN_601 ? _slots_3_io_out_uop_ldq_idx : _GEN_600 ? _slots_2_io_out_uop_ldq_idx : _slots_1_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_602 ? _slots_4_io_out_uop_stq_idx : _GEN_601 ? _slots_3_io_out_uop_stq_idx : _GEN_600 ? _slots_2_io_out_uop_stq_idx : _slots_1_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_602 ? _slots_4_io_out_uop_pdst : _GEN_601 ? _slots_3_io_out_uop_pdst : _GEN_600 ? _slots_2_io_out_uop_pdst : _slots_1_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_602 ? _slots_4_io_out_uop_prs1 : _GEN_601 ? _slots_3_io_out_uop_prs1 : _GEN_600 ? _slots_2_io_out_uop_prs1 : _slots_1_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_602 ? _slots_4_io_out_uop_prs2 : _GEN_601 ? _slots_3_io_out_uop_prs2 : _GEN_600 ? _slots_2_io_out_uop_prs2 : _slots_1_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_602 ? _slots_4_io_out_uop_prs3 : _GEN_601 ? _slots_3_io_out_uop_prs3 : _GEN_600 ? _slots_2_io_out_uop_prs3 : _slots_1_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_602 ? _slots_4_io_out_uop_prs1_busy : _GEN_601 ? _slots_3_io_out_uop_prs1_busy : _GEN_600 ? _slots_2_io_out_uop_prs1_busy : _slots_1_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_602 ? _slots_4_io_out_uop_prs2_busy : _GEN_601 ? _slots_3_io_out_uop_prs2_busy : _GEN_600 ? _slots_2_io_out_uop_prs2_busy : _slots_1_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_602 ? _slots_4_io_out_uop_prs3_busy : _GEN_601 ? _slots_3_io_out_uop_prs3_busy : _GEN_600 ? _slots_2_io_out_uop_prs3_busy : _slots_1_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_602 ? _slots_4_io_out_uop_ppred_busy : _GEN_601 ? _slots_3_io_out_uop_ppred_busy : _GEN_600 ? _slots_2_io_out_uop_ppred_busy : _slots_1_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_602 ? _slots_4_io_out_uop_bypassable : _GEN_601 ? _slots_3_io_out_uop_bypassable : _GEN_600 ? _slots_2_io_out_uop_bypassable : _slots_1_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_602 ? _slots_4_io_out_uop_mem_cmd : _GEN_601 ? _slots_3_io_out_uop_mem_cmd : _GEN_600 ? _slots_2_io_out_uop_mem_cmd : _slots_1_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_602 ? _slots_4_io_out_uop_mem_size : _GEN_601 ? _slots_3_io_out_uop_mem_size : _GEN_600 ? _slots_2_io_out_uop_mem_size : _slots_1_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_602 ? _slots_4_io_out_uop_mem_signed : _GEN_601 ? _slots_3_io_out_uop_mem_signed : _GEN_600 ? _slots_2_io_out_uop_mem_signed : _slots_1_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_602 ? _slots_4_io_out_uop_is_fence : _GEN_601 ? _slots_3_io_out_uop_is_fence : _GEN_600 ? _slots_2_io_out_uop_is_fence : _slots_1_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_602 ? _slots_4_io_out_uop_is_amo : _GEN_601 ? _slots_3_io_out_uop_is_amo : _GEN_600 ? _slots_2_io_out_uop_is_amo : _slots_1_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_602 ? _slots_4_io_out_uop_uses_ldq : _GEN_601 ? _slots_3_io_out_uop_uses_ldq : _GEN_600 ? _slots_2_io_out_uop_uses_ldq : _slots_1_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_602 ? _slots_4_io_out_uop_uses_stq : _GEN_601 ? _slots_3_io_out_uop_uses_stq : _GEN_600 ? _slots_2_io_out_uop_uses_stq : _slots_1_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_602 ? _slots_4_io_out_uop_ldst_val : _GEN_601 ? _slots_3_io_out_uop_ldst_val : _GEN_600 ? _slots_2_io_out_uop_ldst_val : _slots_1_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_602 ? _slots_4_io_out_uop_dst_rtype : _GEN_601 ? _slots_3_io_out_uop_dst_rtype : _GEN_600 ? _slots_2_io_out_uop_dst_rtype : _slots_1_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_602 ? _slots_4_io_out_uop_lrs1_rtype : _GEN_601 ? _slots_3_io_out_uop_lrs1_rtype : _GEN_600 ? _slots_2_io_out_uop_lrs1_rtype : _slots_1_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_602 ? _slots_4_io_out_uop_lrs2_rtype : _GEN_601 ? _slots_3_io_out_uop_lrs2_rtype : _GEN_600 ? _slots_2_io_out_uop_lrs2_rtype : _slots_1_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_602 ? _slots_4_io_out_uop_fp_val : _GEN_601 ? _slots_3_io_out_uop_fp_val : _GEN_600 ? _slots_2_io_out_uop_fp_val : _slots_1_io_out_uop_fp_val),
    .io_valid                       (_slots_0_io_valid),
    .io_will_be_valid               (_slots_0_io_will_be_valid),
    .io_request                     (_slots_0_io_request),
    .io_out_uop_uopc                (/* unused */),
    .io_out_uop_is_rvc              (/* unused */),
    .io_out_uop_fu_code             (/* unused */),
    .io_out_uop_iw_state            (/* unused */),
    .io_out_uop_iw_p1_poisoned      (/* unused */),
    .io_out_uop_iw_p2_poisoned      (/* unused */),
    .io_out_uop_is_br               (/* unused */),
    .io_out_uop_is_jalr             (/* unused */),
    .io_out_uop_is_jal              (/* unused */),
    .io_out_uop_is_sfb              (/* unused */),
    .io_out_uop_br_mask             (/* unused */),
    .io_out_uop_br_tag              (/* unused */),
    .io_out_uop_ftq_idx             (/* unused */),
    .io_out_uop_edge_inst           (/* unused */),
    .io_out_uop_pc_lob              (/* unused */),
    .io_out_uop_taken               (/* unused */),
    .io_out_uop_imm_packed          (/* unused */),
    .io_out_uop_rob_idx             (/* unused */),
    .io_out_uop_ldq_idx             (/* unused */),
    .io_out_uop_stq_idx             (/* unused */),
    .io_out_uop_pdst                (/* unused */),
    .io_out_uop_prs1                (/* unused */),
    .io_out_uop_prs2                (/* unused */),
    .io_out_uop_prs3                (/* unused */),
    .io_out_uop_prs1_busy           (/* unused */),
    .io_out_uop_prs2_busy           (/* unused */),
    .io_out_uop_prs3_busy           (/* unused */),
    .io_out_uop_ppred_busy          (/* unused */),
    .io_out_uop_bypassable          (/* unused */),
    .io_out_uop_mem_cmd             (/* unused */),
    .io_out_uop_mem_size            (/* unused */),
    .io_out_uop_mem_signed          (/* unused */),
    .io_out_uop_is_fence            (/* unused */),
    .io_out_uop_is_amo              (/* unused */),
    .io_out_uop_uses_ldq            (/* unused */),
    .io_out_uop_uses_stq            (/* unused */),
    .io_out_uop_ldst_val            (/* unused */),
    .io_out_uop_dst_rtype           (/* unused */),
    .io_out_uop_lrs1_rtype          (/* unused */),
    .io_out_uop_lrs2_rtype          (/* unused */),
    .io_out_uop_fp_val              (/* unused */),
    .io_uop_uopc                    (_slots_0_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_0_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_0_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_0_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_0_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_0_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_0_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_0_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_0_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_0_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_0_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_0_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_0_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_0_io_uop_pc_lob),
    .io_uop_taken                   (_slots_0_io_uop_taken),
    .io_uop_imm_packed              (_slots_0_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_0_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_0_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_0_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_0_io_uop_pdst),
    .io_uop_prs1                    (_slots_0_io_uop_prs1),
    .io_uop_prs2                    (_slots_0_io_uop_prs2),
    .io_uop_bypassable              (_slots_0_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_0_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_0_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_0_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_0_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_0_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_0_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_0_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_0_io_uop_fp_val)
  );
  IssueSlot_32 slots_1 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_1_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (~_slots_0_io_valid),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_1_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_605 ? _slots_5_io_out_uop_uopc : _GEN_604 ? _slots_4_io_out_uop_uopc : _GEN_603 ? _slots_3_io_out_uop_uopc : _slots_2_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_605 ? _slots_5_io_out_uop_is_rvc : _GEN_604 ? _slots_4_io_out_uop_is_rvc : _GEN_603 ? _slots_3_io_out_uop_is_rvc : _slots_2_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_605 ? _slots_5_io_out_uop_fu_code : _GEN_604 ? _slots_4_io_out_uop_fu_code : _GEN_603 ? _slots_3_io_out_uop_fu_code : _slots_2_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_605 ? _slots_5_io_out_uop_iw_state : _GEN_604 ? _slots_4_io_out_uop_iw_state : _GEN_603 ? _slots_3_io_out_uop_iw_state : _slots_2_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_605 ? _slots_5_io_out_uop_iw_p1_poisoned : _GEN_604 ? _slots_4_io_out_uop_iw_p1_poisoned : _GEN_603 ? _slots_3_io_out_uop_iw_p1_poisoned : _slots_2_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_605 ? _slots_5_io_out_uop_iw_p2_poisoned : _GEN_604 ? _slots_4_io_out_uop_iw_p2_poisoned : _GEN_603 ? _slots_3_io_out_uop_iw_p2_poisoned : _slots_2_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_605 ? _slots_5_io_out_uop_is_br : _GEN_604 ? _slots_4_io_out_uop_is_br : _GEN_603 ? _slots_3_io_out_uop_is_br : _slots_2_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_605 ? _slots_5_io_out_uop_is_jalr : _GEN_604 ? _slots_4_io_out_uop_is_jalr : _GEN_603 ? _slots_3_io_out_uop_is_jalr : _slots_2_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_605 ? _slots_5_io_out_uop_is_jal : _GEN_604 ? _slots_4_io_out_uop_is_jal : _GEN_603 ? _slots_3_io_out_uop_is_jal : _slots_2_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_605 ? _slots_5_io_out_uop_is_sfb : _GEN_604 ? _slots_4_io_out_uop_is_sfb : _GEN_603 ? _slots_3_io_out_uop_is_sfb : _slots_2_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_605 ? _slots_5_io_out_uop_br_mask : _GEN_604 ? _slots_4_io_out_uop_br_mask : _GEN_603 ? _slots_3_io_out_uop_br_mask : _slots_2_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_605 ? _slots_5_io_out_uop_br_tag : _GEN_604 ? _slots_4_io_out_uop_br_tag : _GEN_603 ? _slots_3_io_out_uop_br_tag : _slots_2_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_605 ? _slots_5_io_out_uop_ftq_idx : _GEN_604 ? _slots_4_io_out_uop_ftq_idx : _GEN_603 ? _slots_3_io_out_uop_ftq_idx : _slots_2_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_605 ? _slots_5_io_out_uop_edge_inst : _GEN_604 ? _slots_4_io_out_uop_edge_inst : _GEN_603 ? _slots_3_io_out_uop_edge_inst : _slots_2_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_605 ? _slots_5_io_out_uop_pc_lob : _GEN_604 ? _slots_4_io_out_uop_pc_lob : _GEN_603 ? _slots_3_io_out_uop_pc_lob : _slots_2_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_605 ? _slots_5_io_out_uop_taken : _GEN_604 ? _slots_4_io_out_uop_taken : _GEN_603 ? _slots_3_io_out_uop_taken : _slots_2_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_605 ? _slots_5_io_out_uop_imm_packed : _GEN_604 ? _slots_4_io_out_uop_imm_packed : _GEN_603 ? _slots_3_io_out_uop_imm_packed : _slots_2_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_605 ? _slots_5_io_out_uop_rob_idx : _GEN_604 ? _slots_4_io_out_uop_rob_idx : _GEN_603 ? _slots_3_io_out_uop_rob_idx : _slots_2_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_605 ? _slots_5_io_out_uop_ldq_idx : _GEN_604 ? _slots_4_io_out_uop_ldq_idx : _GEN_603 ? _slots_3_io_out_uop_ldq_idx : _slots_2_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_605 ? _slots_5_io_out_uop_stq_idx : _GEN_604 ? _slots_4_io_out_uop_stq_idx : _GEN_603 ? _slots_3_io_out_uop_stq_idx : _slots_2_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_605 ? _slots_5_io_out_uop_pdst : _GEN_604 ? _slots_4_io_out_uop_pdst : _GEN_603 ? _slots_3_io_out_uop_pdst : _slots_2_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_605 ? _slots_5_io_out_uop_prs1 : _GEN_604 ? _slots_4_io_out_uop_prs1 : _GEN_603 ? _slots_3_io_out_uop_prs1 : _slots_2_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_605 ? _slots_5_io_out_uop_prs2 : _GEN_604 ? _slots_4_io_out_uop_prs2 : _GEN_603 ? _slots_3_io_out_uop_prs2 : _slots_2_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_605 ? _slots_5_io_out_uop_prs3 : _GEN_604 ? _slots_4_io_out_uop_prs3 : _GEN_603 ? _slots_3_io_out_uop_prs3 : _slots_2_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_605 ? _slots_5_io_out_uop_prs1_busy : _GEN_604 ? _slots_4_io_out_uop_prs1_busy : _GEN_603 ? _slots_3_io_out_uop_prs1_busy : _slots_2_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_605 ? _slots_5_io_out_uop_prs2_busy : _GEN_604 ? _slots_4_io_out_uop_prs2_busy : _GEN_603 ? _slots_3_io_out_uop_prs2_busy : _slots_2_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_605 ? _slots_5_io_out_uop_prs3_busy : _GEN_604 ? _slots_4_io_out_uop_prs3_busy : _GEN_603 ? _slots_3_io_out_uop_prs3_busy : _slots_2_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_605 ? _slots_5_io_out_uop_ppred_busy : _GEN_604 ? _slots_4_io_out_uop_ppred_busy : _GEN_603 ? _slots_3_io_out_uop_ppred_busy : _slots_2_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_605 ? _slots_5_io_out_uop_bypassable : _GEN_604 ? _slots_4_io_out_uop_bypassable : _GEN_603 ? _slots_3_io_out_uop_bypassable : _slots_2_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_605 ? _slots_5_io_out_uop_mem_cmd : _GEN_604 ? _slots_4_io_out_uop_mem_cmd : _GEN_603 ? _slots_3_io_out_uop_mem_cmd : _slots_2_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_605 ? _slots_5_io_out_uop_mem_size : _GEN_604 ? _slots_4_io_out_uop_mem_size : _GEN_603 ? _slots_3_io_out_uop_mem_size : _slots_2_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_605 ? _slots_5_io_out_uop_mem_signed : _GEN_604 ? _slots_4_io_out_uop_mem_signed : _GEN_603 ? _slots_3_io_out_uop_mem_signed : _slots_2_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_605 ? _slots_5_io_out_uop_is_fence : _GEN_604 ? _slots_4_io_out_uop_is_fence : _GEN_603 ? _slots_3_io_out_uop_is_fence : _slots_2_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_605 ? _slots_5_io_out_uop_is_amo : _GEN_604 ? _slots_4_io_out_uop_is_amo : _GEN_603 ? _slots_3_io_out_uop_is_amo : _slots_2_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_605 ? _slots_5_io_out_uop_uses_ldq : _GEN_604 ? _slots_4_io_out_uop_uses_ldq : _GEN_603 ? _slots_3_io_out_uop_uses_ldq : _slots_2_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_605 ? _slots_5_io_out_uop_uses_stq : _GEN_604 ? _slots_4_io_out_uop_uses_stq : _GEN_603 ? _slots_3_io_out_uop_uses_stq : _slots_2_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_605 ? _slots_5_io_out_uop_ldst_val : _GEN_604 ? _slots_4_io_out_uop_ldst_val : _GEN_603 ? _slots_3_io_out_uop_ldst_val : _slots_2_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_605 ? _slots_5_io_out_uop_dst_rtype : _GEN_604 ? _slots_4_io_out_uop_dst_rtype : _GEN_603 ? _slots_3_io_out_uop_dst_rtype : _slots_2_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_605 ? _slots_5_io_out_uop_lrs1_rtype : _GEN_604 ? _slots_4_io_out_uop_lrs1_rtype : _GEN_603 ? _slots_3_io_out_uop_lrs1_rtype : _slots_2_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_605 ? _slots_5_io_out_uop_lrs2_rtype : _GEN_604 ? _slots_4_io_out_uop_lrs2_rtype : _GEN_603 ? _slots_3_io_out_uop_lrs2_rtype : _slots_2_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_605 ? _slots_5_io_out_uop_fp_val : _GEN_604 ? _slots_4_io_out_uop_fp_val : _GEN_603 ? _slots_3_io_out_uop_fp_val : _slots_2_io_out_uop_fp_val),
    .io_valid                       (_slots_1_io_valid),
    .io_will_be_valid               (_slots_1_io_will_be_valid),
    .io_request                     (_slots_1_io_request),
    .io_out_uop_uopc                (_slots_1_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_1_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_1_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_1_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_1_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_1_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_1_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_1_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_1_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_1_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_1_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_1_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_1_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_1_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_1_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_1_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_1_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_1_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_1_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_1_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_1_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_1_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_1_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_1_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_1_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_1_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_1_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_1_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_1_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_1_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_1_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_1_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_1_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_1_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_1_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_1_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_1_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_1_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_1_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_1_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_1_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_1_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_1_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_1_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_1_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_1_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_1_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_1_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_1_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_1_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_1_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_1_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_1_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_1_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_1_io_uop_pc_lob),
    .io_uop_taken                   (_slots_1_io_uop_taken),
    .io_uop_imm_packed              (_slots_1_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_1_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_1_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_1_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_1_io_uop_pdst),
    .io_uop_prs1                    (_slots_1_io_uop_prs1),
    .io_uop_prs2                    (_slots_1_io_uop_prs2),
    .io_uop_bypassable              (_slots_1_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_1_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_1_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_1_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_1_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_1_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_1_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_1_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_1_io_uop_fp_val)
  );
  IssueSlot_32 slots_2 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_2_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_23_1to0),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_2_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_608 ? _slots_6_io_out_uop_uopc : _GEN_607 ? _slots_5_io_out_uop_uopc : _GEN_606 ? _slots_4_io_out_uop_uopc : _slots_3_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_608 ? _slots_6_io_out_uop_is_rvc : _GEN_607 ? _slots_5_io_out_uop_is_rvc : _GEN_606 ? _slots_4_io_out_uop_is_rvc : _slots_3_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_608 ? _slots_6_io_out_uop_fu_code : _GEN_607 ? _slots_5_io_out_uop_fu_code : _GEN_606 ? _slots_4_io_out_uop_fu_code : _slots_3_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_608 ? _slots_6_io_out_uop_iw_state : _GEN_607 ? _slots_5_io_out_uop_iw_state : _GEN_606 ? _slots_4_io_out_uop_iw_state : _slots_3_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_608 ? _slots_6_io_out_uop_iw_p1_poisoned : _GEN_607 ? _slots_5_io_out_uop_iw_p1_poisoned : _GEN_606 ? _slots_4_io_out_uop_iw_p1_poisoned : _slots_3_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_608 ? _slots_6_io_out_uop_iw_p2_poisoned : _GEN_607 ? _slots_5_io_out_uop_iw_p2_poisoned : _GEN_606 ? _slots_4_io_out_uop_iw_p2_poisoned : _slots_3_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_608 ? _slots_6_io_out_uop_is_br : _GEN_607 ? _slots_5_io_out_uop_is_br : _GEN_606 ? _slots_4_io_out_uop_is_br : _slots_3_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_608 ? _slots_6_io_out_uop_is_jalr : _GEN_607 ? _slots_5_io_out_uop_is_jalr : _GEN_606 ? _slots_4_io_out_uop_is_jalr : _slots_3_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_608 ? _slots_6_io_out_uop_is_jal : _GEN_607 ? _slots_5_io_out_uop_is_jal : _GEN_606 ? _slots_4_io_out_uop_is_jal : _slots_3_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_608 ? _slots_6_io_out_uop_is_sfb : _GEN_607 ? _slots_5_io_out_uop_is_sfb : _GEN_606 ? _slots_4_io_out_uop_is_sfb : _slots_3_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_608 ? _slots_6_io_out_uop_br_mask : _GEN_607 ? _slots_5_io_out_uop_br_mask : _GEN_606 ? _slots_4_io_out_uop_br_mask : _slots_3_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_608 ? _slots_6_io_out_uop_br_tag : _GEN_607 ? _slots_5_io_out_uop_br_tag : _GEN_606 ? _slots_4_io_out_uop_br_tag : _slots_3_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_608 ? _slots_6_io_out_uop_ftq_idx : _GEN_607 ? _slots_5_io_out_uop_ftq_idx : _GEN_606 ? _slots_4_io_out_uop_ftq_idx : _slots_3_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_608 ? _slots_6_io_out_uop_edge_inst : _GEN_607 ? _slots_5_io_out_uop_edge_inst : _GEN_606 ? _slots_4_io_out_uop_edge_inst : _slots_3_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_608 ? _slots_6_io_out_uop_pc_lob : _GEN_607 ? _slots_5_io_out_uop_pc_lob : _GEN_606 ? _slots_4_io_out_uop_pc_lob : _slots_3_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_608 ? _slots_6_io_out_uop_taken : _GEN_607 ? _slots_5_io_out_uop_taken : _GEN_606 ? _slots_4_io_out_uop_taken : _slots_3_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_608 ? _slots_6_io_out_uop_imm_packed : _GEN_607 ? _slots_5_io_out_uop_imm_packed : _GEN_606 ? _slots_4_io_out_uop_imm_packed : _slots_3_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_608 ? _slots_6_io_out_uop_rob_idx : _GEN_607 ? _slots_5_io_out_uop_rob_idx : _GEN_606 ? _slots_4_io_out_uop_rob_idx : _slots_3_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_608 ? _slots_6_io_out_uop_ldq_idx : _GEN_607 ? _slots_5_io_out_uop_ldq_idx : _GEN_606 ? _slots_4_io_out_uop_ldq_idx : _slots_3_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_608 ? _slots_6_io_out_uop_stq_idx : _GEN_607 ? _slots_5_io_out_uop_stq_idx : _GEN_606 ? _slots_4_io_out_uop_stq_idx : _slots_3_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_608 ? _slots_6_io_out_uop_pdst : _GEN_607 ? _slots_5_io_out_uop_pdst : _GEN_606 ? _slots_4_io_out_uop_pdst : _slots_3_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_608 ? _slots_6_io_out_uop_prs1 : _GEN_607 ? _slots_5_io_out_uop_prs1 : _GEN_606 ? _slots_4_io_out_uop_prs1 : _slots_3_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_608 ? _slots_6_io_out_uop_prs2 : _GEN_607 ? _slots_5_io_out_uop_prs2 : _GEN_606 ? _slots_4_io_out_uop_prs2 : _slots_3_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_608 ? _slots_6_io_out_uop_prs3 : _GEN_607 ? _slots_5_io_out_uop_prs3 : _GEN_606 ? _slots_4_io_out_uop_prs3 : _slots_3_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_608 ? _slots_6_io_out_uop_prs1_busy : _GEN_607 ? _slots_5_io_out_uop_prs1_busy : _GEN_606 ? _slots_4_io_out_uop_prs1_busy : _slots_3_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_608 ? _slots_6_io_out_uop_prs2_busy : _GEN_607 ? _slots_5_io_out_uop_prs2_busy : _GEN_606 ? _slots_4_io_out_uop_prs2_busy : _slots_3_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_608 ? _slots_6_io_out_uop_prs3_busy : _GEN_607 ? _slots_5_io_out_uop_prs3_busy : _GEN_606 ? _slots_4_io_out_uop_prs3_busy : _slots_3_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_608 ? _slots_6_io_out_uop_ppred_busy : _GEN_607 ? _slots_5_io_out_uop_ppred_busy : _GEN_606 ? _slots_4_io_out_uop_ppred_busy : _slots_3_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_608 ? _slots_6_io_out_uop_bypassable : _GEN_607 ? _slots_5_io_out_uop_bypassable : _GEN_606 ? _slots_4_io_out_uop_bypassable : _slots_3_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_608 ? _slots_6_io_out_uop_mem_cmd : _GEN_607 ? _slots_5_io_out_uop_mem_cmd : _GEN_606 ? _slots_4_io_out_uop_mem_cmd : _slots_3_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_608 ? _slots_6_io_out_uop_mem_size : _GEN_607 ? _slots_5_io_out_uop_mem_size : _GEN_606 ? _slots_4_io_out_uop_mem_size : _slots_3_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_608 ? _slots_6_io_out_uop_mem_signed : _GEN_607 ? _slots_5_io_out_uop_mem_signed : _GEN_606 ? _slots_4_io_out_uop_mem_signed : _slots_3_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_608 ? _slots_6_io_out_uop_is_fence : _GEN_607 ? _slots_5_io_out_uop_is_fence : _GEN_606 ? _slots_4_io_out_uop_is_fence : _slots_3_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_608 ? _slots_6_io_out_uop_is_amo : _GEN_607 ? _slots_5_io_out_uop_is_amo : _GEN_606 ? _slots_4_io_out_uop_is_amo : _slots_3_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_608 ? _slots_6_io_out_uop_uses_ldq : _GEN_607 ? _slots_5_io_out_uop_uses_ldq : _GEN_606 ? _slots_4_io_out_uop_uses_ldq : _slots_3_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_608 ? _slots_6_io_out_uop_uses_stq : _GEN_607 ? _slots_5_io_out_uop_uses_stq : _GEN_606 ? _slots_4_io_out_uop_uses_stq : _slots_3_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_608 ? _slots_6_io_out_uop_ldst_val : _GEN_607 ? _slots_5_io_out_uop_ldst_val : _GEN_606 ? _slots_4_io_out_uop_ldst_val : _slots_3_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_608 ? _slots_6_io_out_uop_dst_rtype : _GEN_607 ? _slots_5_io_out_uop_dst_rtype : _GEN_606 ? _slots_4_io_out_uop_dst_rtype : _slots_3_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_608 ? _slots_6_io_out_uop_lrs1_rtype : _GEN_607 ? _slots_5_io_out_uop_lrs1_rtype : _GEN_606 ? _slots_4_io_out_uop_lrs1_rtype : _slots_3_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_608 ? _slots_6_io_out_uop_lrs2_rtype : _GEN_607 ? _slots_5_io_out_uop_lrs2_rtype : _GEN_606 ? _slots_4_io_out_uop_lrs2_rtype : _slots_3_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_608 ? _slots_6_io_out_uop_fp_val : _GEN_607 ? _slots_5_io_out_uop_fp_val : _GEN_606 ? _slots_4_io_out_uop_fp_val : _slots_3_io_out_uop_fp_val),
    .io_valid                       (_slots_2_io_valid),
    .io_will_be_valid               (_slots_2_io_will_be_valid),
    .io_request                     (_slots_2_io_request),
    .io_out_uop_uopc                (_slots_2_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_2_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_2_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_2_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_2_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_2_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_2_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_2_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_2_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_2_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_2_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_2_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_2_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_2_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_2_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_2_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_2_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_2_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_2_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_2_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_2_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_2_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_2_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_2_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_2_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_2_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_2_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_2_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_2_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_2_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_2_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_2_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_2_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_2_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_2_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_2_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_2_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_2_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_2_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_2_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_2_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_2_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_2_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_2_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_2_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_2_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_2_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_2_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_2_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_2_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_2_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_2_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_2_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_2_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_2_io_uop_pc_lob),
    .io_uop_taken                   (_slots_2_io_uop_taken),
    .io_uop_imm_packed              (_slots_2_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_2_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_2_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_2_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_2_io_uop_pdst),
    .io_uop_prs1                    (_slots_2_io_uop_prs1),
    .io_uop_prs2                    (_slots_2_io_uop_prs2),
    .io_uop_bypassable              (_slots_2_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_2_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_2_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_2_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_2_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_2_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_2_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_2_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_2_io_uop_fp_val)
  );
  IssueSlot_32 slots_3 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_3_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_25),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_3_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_611 ? _slots_7_io_out_uop_uopc : _GEN_610 ? _slots_6_io_out_uop_uopc : _GEN_609 ? _slots_5_io_out_uop_uopc : _slots_4_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_611 ? _slots_7_io_out_uop_is_rvc : _GEN_610 ? _slots_6_io_out_uop_is_rvc : _GEN_609 ? _slots_5_io_out_uop_is_rvc : _slots_4_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_611 ? _slots_7_io_out_uop_fu_code : _GEN_610 ? _slots_6_io_out_uop_fu_code : _GEN_609 ? _slots_5_io_out_uop_fu_code : _slots_4_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_611 ? _slots_7_io_out_uop_iw_state : _GEN_610 ? _slots_6_io_out_uop_iw_state : _GEN_609 ? _slots_5_io_out_uop_iw_state : _slots_4_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_611 ? _slots_7_io_out_uop_iw_p1_poisoned : _GEN_610 ? _slots_6_io_out_uop_iw_p1_poisoned : _GEN_609 ? _slots_5_io_out_uop_iw_p1_poisoned : _slots_4_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_611 ? _slots_7_io_out_uop_iw_p2_poisoned : _GEN_610 ? _slots_6_io_out_uop_iw_p2_poisoned : _GEN_609 ? _slots_5_io_out_uop_iw_p2_poisoned : _slots_4_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_611 ? _slots_7_io_out_uop_is_br : _GEN_610 ? _slots_6_io_out_uop_is_br : _GEN_609 ? _slots_5_io_out_uop_is_br : _slots_4_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_611 ? _slots_7_io_out_uop_is_jalr : _GEN_610 ? _slots_6_io_out_uop_is_jalr : _GEN_609 ? _slots_5_io_out_uop_is_jalr : _slots_4_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_611 ? _slots_7_io_out_uop_is_jal : _GEN_610 ? _slots_6_io_out_uop_is_jal : _GEN_609 ? _slots_5_io_out_uop_is_jal : _slots_4_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_611 ? _slots_7_io_out_uop_is_sfb : _GEN_610 ? _slots_6_io_out_uop_is_sfb : _GEN_609 ? _slots_5_io_out_uop_is_sfb : _slots_4_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_611 ? _slots_7_io_out_uop_br_mask : _GEN_610 ? _slots_6_io_out_uop_br_mask : _GEN_609 ? _slots_5_io_out_uop_br_mask : _slots_4_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_611 ? _slots_7_io_out_uop_br_tag : _GEN_610 ? _slots_6_io_out_uop_br_tag : _GEN_609 ? _slots_5_io_out_uop_br_tag : _slots_4_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_611 ? _slots_7_io_out_uop_ftq_idx : _GEN_610 ? _slots_6_io_out_uop_ftq_idx : _GEN_609 ? _slots_5_io_out_uop_ftq_idx : _slots_4_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_611 ? _slots_7_io_out_uop_edge_inst : _GEN_610 ? _slots_6_io_out_uop_edge_inst : _GEN_609 ? _slots_5_io_out_uop_edge_inst : _slots_4_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_611 ? _slots_7_io_out_uop_pc_lob : _GEN_610 ? _slots_6_io_out_uop_pc_lob : _GEN_609 ? _slots_5_io_out_uop_pc_lob : _slots_4_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_611 ? _slots_7_io_out_uop_taken : _GEN_610 ? _slots_6_io_out_uop_taken : _GEN_609 ? _slots_5_io_out_uop_taken : _slots_4_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_611 ? _slots_7_io_out_uop_imm_packed : _GEN_610 ? _slots_6_io_out_uop_imm_packed : _GEN_609 ? _slots_5_io_out_uop_imm_packed : _slots_4_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_611 ? _slots_7_io_out_uop_rob_idx : _GEN_610 ? _slots_6_io_out_uop_rob_idx : _GEN_609 ? _slots_5_io_out_uop_rob_idx : _slots_4_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_611 ? _slots_7_io_out_uop_ldq_idx : _GEN_610 ? _slots_6_io_out_uop_ldq_idx : _GEN_609 ? _slots_5_io_out_uop_ldq_idx : _slots_4_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_611 ? _slots_7_io_out_uop_stq_idx : _GEN_610 ? _slots_6_io_out_uop_stq_idx : _GEN_609 ? _slots_5_io_out_uop_stq_idx : _slots_4_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_611 ? _slots_7_io_out_uop_pdst : _GEN_610 ? _slots_6_io_out_uop_pdst : _GEN_609 ? _slots_5_io_out_uop_pdst : _slots_4_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_611 ? _slots_7_io_out_uop_prs1 : _GEN_610 ? _slots_6_io_out_uop_prs1 : _GEN_609 ? _slots_5_io_out_uop_prs1 : _slots_4_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_611 ? _slots_7_io_out_uop_prs2 : _GEN_610 ? _slots_6_io_out_uop_prs2 : _GEN_609 ? _slots_5_io_out_uop_prs2 : _slots_4_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_611 ? _slots_7_io_out_uop_prs3 : _GEN_610 ? _slots_6_io_out_uop_prs3 : _GEN_609 ? _slots_5_io_out_uop_prs3 : _slots_4_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_611 ? _slots_7_io_out_uop_prs1_busy : _GEN_610 ? _slots_6_io_out_uop_prs1_busy : _GEN_609 ? _slots_5_io_out_uop_prs1_busy : _slots_4_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_611 ? _slots_7_io_out_uop_prs2_busy : _GEN_610 ? _slots_6_io_out_uop_prs2_busy : _GEN_609 ? _slots_5_io_out_uop_prs2_busy : _slots_4_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_611 ? _slots_7_io_out_uop_prs3_busy : _GEN_610 ? _slots_6_io_out_uop_prs3_busy : _GEN_609 ? _slots_5_io_out_uop_prs3_busy : _slots_4_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_611 ? _slots_7_io_out_uop_ppred_busy : _GEN_610 ? _slots_6_io_out_uop_ppred_busy : _GEN_609 ? _slots_5_io_out_uop_ppred_busy : _slots_4_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_611 ? _slots_7_io_out_uop_bypassable : _GEN_610 ? _slots_6_io_out_uop_bypassable : _GEN_609 ? _slots_5_io_out_uop_bypassable : _slots_4_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_611 ? _slots_7_io_out_uop_mem_cmd : _GEN_610 ? _slots_6_io_out_uop_mem_cmd : _GEN_609 ? _slots_5_io_out_uop_mem_cmd : _slots_4_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_611 ? _slots_7_io_out_uop_mem_size : _GEN_610 ? _slots_6_io_out_uop_mem_size : _GEN_609 ? _slots_5_io_out_uop_mem_size : _slots_4_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_611 ? _slots_7_io_out_uop_mem_signed : _GEN_610 ? _slots_6_io_out_uop_mem_signed : _GEN_609 ? _slots_5_io_out_uop_mem_signed : _slots_4_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_611 ? _slots_7_io_out_uop_is_fence : _GEN_610 ? _slots_6_io_out_uop_is_fence : _GEN_609 ? _slots_5_io_out_uop_is_fence : _slots_4_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_611 ? _slots_7_io_out_uop_is_amo : _GEN_610 ? _slots_6_io_out_uop_is_amo : _GEN_609 ? _slots_5_io_out_uop_is_amo : _slots_4_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_611 ? _slots_7_io_out_uop_uses_ldq : _GEN_610 ? _slots_6_io_out_uop_uses_ldq : _GEN_609 ? _slots_5_io_out_uop_uses_ldq : _slots_4_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_611 ? _slots_7_io_out_uop_uses_stq : _GEN_610 ? _slots_6_io_out_uop_uses_stq : _GEN_609 ? _slots_5_io_out_uop_uses_stq : _slots_4_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_611 ? _slots_7_io_out_uop_ldst_val : _GEN_610 ? _slots_6_io_out_uop_ldst_val : _GEN_609 ? _slots_5_io_out_uop_ldst_val : _slots_4_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_611 ? _slots_7_io_out_uop_dst_rtype : _GEN_610 ? _slots_6_io_out_uop_dst_rtype : _GEN_609 ? _slots_5_io_out_uop_dst_rtype : _slots_4_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_611 ? _slots_7_io_out_uop_lrs1_rtype : _GEN_610 ? _slots_6_io_out_uop_lrs1_rtype : _GEN_609 ? _slots_5_io_out_uop_lrs1_rtype : _slots_4_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_611 ? _slots_7_io_out_uop_lrs2_rtype : _GEN_610 ? _slots_6_io_out_uop_lrs2_rtype : _GEN_609 ? _slots_5_io_out_uop_lrs2_rtype : _slots_4_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_611 ? _slots_7_io_out_uop_fp_val : _GEN_610 ? _slots_6_io_out_uop_fp_val : _GEN_609 ? _slots_5_io_out_uop_fp_val : _slots_4_io_out_uop_fp_val),
    .io_valid                       (_slots_3_io_valid),
    .io_will_be_valid               (_slots_3_io_will_be_valid),
    .io_request                     (_slots_3_io_request),
    .io_out_uop_uopc                (_slots_3_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_3_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_3_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_3_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_3_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_3_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_3_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_3_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_3_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_3_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_3_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_3_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_3_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_3_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_3_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_3_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_3_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_3_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_3_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_3_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_3_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_3_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_3_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_3_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_3_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_3_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_3_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_3_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_3_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_3_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_3_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_3_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_3_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_3_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_3_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_3_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_3_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_3_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_3_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_3_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_3_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_3_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_3_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_3_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_3_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_3_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_3_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_3_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_3_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_3_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_3_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_3_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_3_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_3_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_3_io_uop_pc_lob),
    .io_uop_taken                   (_slots_3_io_uop_taken),
    .io_uop_imm_packed              (_slots_3_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_3_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_3_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_3_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_3_io_uop_pdst),
    .io_uop_prs1                    (_slots_3_io_uop_prs1),
    .io_uop_prs2                    (_slots_3_io_uop_prs2),
    .io_uop_bypassable              (_slots_3_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_3_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_3_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_3_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_3_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_3_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_3_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_3_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_3_io_uop_fp_val)
  );
  IssueSlot_32 slots_4 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_4_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_27),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_4_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_614 ? _slots_8_io_out_uop_uopc : _GEN_613 ? _slots_7_io_out_uop_uopc : _GEN_612 ? _slots_6_io_out_uop_uopc : _slots_5_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_614 ? _slots_8_io_out_uop_is_rvc : _GEN_613 ? _slots_7_io_out_uop_is_rvc : _GEN_612 ? _slots_6_io_out_uop_is_rvc : _slots_5_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_614 ? _slots_8_io_out_uop_fu_code : _GEN_613 ? _slots_7_io_out_uop_fu_code : _GEN_612 ? _slots_6_io_out_uop_fu_code : _slots_5_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_614 ? _slots_8_io_out_uop_iw_state : _GEN_613 ? _slots_7_io_out_uop_iw_state : _GEN_612 ? _slots_6_io_out_uop_iw_state : _slots_5_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_614 ? _slots_8_io_out_uop_iw_p1_poisoned : _GEN_613 ? _slots_7_io_out_uop_iw_p1_poisoned : _GEN_612 ? _slots_6_io_out_uop_iw_p1_poisoned : _slots_5_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_614 ? _slots_8_io_out_uop_iw_p2_poisoned : _GEN_613 ? _slots_7_io_out_uop_iw_p2_poisoned : _GEN_612 ? _slots_6_io_out_uop_iw_p2_poisoned : _slots_5_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_614 ? _slots_8_io_out_uop_is_br : _GEN_613 ? _slots_7_io_out_uop_is_br : _GEN_612 ? _slots_6_io_out_uop_is_br : _slots_5_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_614 ? _slots_8_io_out_uop_is_jalr : _GEN_613 ? _slots_7_io_out_uop_is_jalr : _GEN_612 ? _slots_6_io_out_uop_is_jalr : _slots_5_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_614 ? _slots_8_io_out_uop_is_jal : _GEN_613 ? _slots_7_io_out_uop_is_jal : _GEN_612 ? _slots_6_io_out_uop_is_jal : _slots_5_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_614 ? _slots_8_io_out_uop_is_sfb : _GEN_613 ? _slots_7_io_out_uop_is_sfb : _GEN_612 ? _slots_6_io_out_uop_is_sfb : _slots_5_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_614 ? _slots_8_io_out_uop_br_mask : _GEN_613 ? _slots_7_io_out_uop_br_mask : _GEN_612 ? _slots_6_io_out_uop_br_mask : _slots_5_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_614 ? _slots_8_io_out_uop_br_tag : _GEN_613 ? _slots_7_io_out_uop_br_tag : _GEN_612 ? _slots_6_io_out_uop_br_tag : _slots_5_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_614 ? _slots_8_io_out_uop_ftq_idx : _GEN_613 ? _slots_7_io_out_uop_ftq_idx : _GEN_612 ? _slots_6_io_out_uop_ftq_idx : _slots_5_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_614 ? _slots_8_io_out_uop_edge_inst : _GEN_613 ? _slots_7_io_out_uop_edge_inst : _GEN_612 ? _slots_6_io_out_uop_edge_inst : _slots_5_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_614 ? _slots_8_io_out_uop_pc_lob : _GEN_613 ? _slots_7_io_out_uop_pc_lob : _GEN_612 ? _slots_6_io_out_uop_pc_lob : _slots_5_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_614 ? _slots_8_io_out_uop_taken : _GEN_613 ? _slots_7_io_out_uop_taken : _GEN_612 ? _slots_6_io_out_uop_taken : _slots_5_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_614 ? _slots_8_io_out_uop_imm_packed : _GEN_613 ? _slots_7_io_out_uop_imm_packed : _GEN_612 ? _slots_6_io_out_uop_imm_packed : _slots_5_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_614 ? _slots_8_io_out_uop_rob_idx : _GEN_613 ? _slots_7_io_out_uop_rob_idx : _GEN_612 ? _slots_6_io_out_uop_rob_idx : _slots_5_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_614 ? _slots_8_io_out_uop_ldq_idx : _GEN_613 ? _slots_7_io_out_uop_ldq_idx : _GEN_612 ? _slots_6_io_out_uop_ldq_idx : _slots_5_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_614 ? _slots_8_io_out_uop_stq_idx : _GEN_613 ? _slots_7_io_out_uop_stq_idx : _GEN_612 ? _slots_6_io_out_uop_stq_idx : _slots_5_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_614 ? _slots_8_io_out_uop_pdst : _GEN_613 ? _slots_7_io_out_uop_pdst : _GEN_612 ? _slots_6_io_out_uop_pdst : _slots_5_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_614 ? _slots_8_io_out_uop_prs1 : _GEN_613 ? _slots_7_io_out_uop_prs1 : _GEN_612 ? _slots_6_io_out_uop_prs1 : _slots_5_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_614 ? _slots_8_io_out_uop_prs2 : _GEN_613 ? _slots_7_io_out_uop_prs2 : _GEN_612 ? _slots_6_io_out_uop_prs2 : _slots_5_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_614 ? _slots_8_io_out_uop_prs3 : _GEN_613 ? _slots_7_io_out_uop_prs3 : _GEN_612 ? _slots_6_io_out_uop_prs3 : _slots_5_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_614 ? _slots_8_io_out_uop_prs1_busy : _GEN_613 ? _slots_7_io_out_uop_prs1_busy : _GEN_612 ? _slots_6_io_out_uop_prs1_busy : _slots_5_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_614 ? _slots_8_io_out_uop_prs2_busy : _GEN_613 ? _slots_7_io_out_uop_prs2_busy : _GEN_612 ? _slots_6_io_out_uop_prs2_busy : _slots_5_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_614 ? _slots_8_io_out_uop_prs3_busy : _GEN_613 ? _slots_7_io_out_uop_prs3_busy : _GEN_612 ? _slots_6_io_out_uop_prs3_busy : _slots_5_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_614 ? _slots_8_io_out_uop_ppred_busy : _GEN_613 ? _slots_7_io_out_uop_ppred_busy : _GEN_612 ? _slots_6_io_out_uop_ppred_busy : _slots_5_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_614 ? _slots_8_io_out_uop_bypassable : _GEN_613 ? _slots_7_io_out_uop_bypassable : _GEN_612 ? _slots_6_io_out_uop_bypassable : _slots_5_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_614 ? _slots_8_io_out_uop_mem_cmd : _GEN_613 ? _slots_7_io_out_uop_mem_cmd : _GEN_612 ? _slots_6_io_out_uop_mem_cmd : _slots_5_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_614 ? _slots_8_io_out_uop_mem_size : _GEN_613 ? _slots_7_io_out_uop_mem_size : _GEN_612 ? _slots_6_io_out_uop_mem_size : _slots_5_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_614 ? _slots_8_io_out_uop_mem_signed : _GEN_613 ? _slots_7_io_out_uop_mem_signed : _GEN_612 ? _slots_6_io_out_uop_mem_signed : _slots_5_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_614 ? _slots_8_io_out_uop_is_fence : _GEN_613 ? _slots_7_io_out_uop_is_fence : _GEN_612 ? _slots_6_io_out_uop_is_fence : _slots_5_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_614 ? _slots_8_io_out_uop_is_amo : _GEN_613 ? _slots_7_io_out_uop_is_amo : _GEN_612 ? _slots_6_io_out_uop_is_amo : _slots_5_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_614 ? _slots_8_io_out_uop_uses_ldq : _GEN_613 ? _slots_7_io_out_uop_uses_ldq : _GEN_612 ? _slots_6_io_out_uop_uses_ldq : _slots_5_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_614 ? _slots_8_io_out_uop_uses_stq : _GEN_613 ? _slots_7_io_out_uop_uses_stq : _GEN_612 ? _slots_6_io_out_uop_uses_stq : _slots_5_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_614 ? _slots_8_io_out_uop_ldst_val : _GEN_613 ? _slots_7_io_out_uop_ldst_val : _GEN_612 ? _slots_6_io_out_uop_ldst_val : _slots_5_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_614 ? _slots_8_io_out_uop_dst_rtype : _GEN_613 ? _slots_7_io_out_uop_dst_rtype : _GEN_612 ? _slots_6_io_out_uop_dst_rtype : _slots_5_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_614 ? _slots_8_io_out_uop_lrs1_rtype : _GEN_613 ? _slots_7_io_out_uop_lrs1_rtype : _GEN_612 ? _slots_6_io_out_uop_lrs1_rtype : _slots_5_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_614 ? _slots_8_io_out_uop_lrs2_rtype : _GEN_613 ? _slots_7_io_out_uop_lrs2_rtype : _GEN_612 ? _slots_6_io_out_uop_lrs2_rtype : _slots_5_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_614 ? _slots_8_io_out_uop_fp_val : _GEN_613 ? _slots_7_io_out_uop_fp_val : _GEN_612 ? _slots_6_io_out_uop_fp_val : _slots_5_io_out_uop_fp_val),
    .io_valid                       (_slots_4_io_valid),
    .io_will_be_valid               (_slots_4_io_will_be_valid),
    .io_request                     (_slots_4_io_request),
    .io_out_uop_uopc                (_slots_4_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_4_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_4_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_4_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_4_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_4_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_4_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_4_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_4_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_4_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_4_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_4_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_4_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_4_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_4_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_4_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_4_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_4_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_4_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_4_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_4_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_4_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_4_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_4_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_4_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_4_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_4_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_4_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_4_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_4_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_4_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_4_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_4_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_4_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_4_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_4_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_4_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_4_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_4_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_4_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_4_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_4_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_4_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_4_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_4_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_4_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_4_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_4_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_4_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_4_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_4_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_4_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_4_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_4_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_4_io_uop_pc_lob),
    .io_uop_taken                   (_slots_4_io_uop_taken),
    .io_uop_imm_packed              (_slots_4_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_4_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_4_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_4_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_4_io_uop_pdst),
    .io_uop_prs1                    (_slots_4_io_uop_prs1),
    .io_uop_prs2                    (_slots_4_io_uop_prs2),
    .io_uop_bypassable              (_slots_4_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_4_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_4_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_4_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_4_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_4_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_4_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_4_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_4_io_uop_fp_val)
  );
  IssueSlot_32 slots_5 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_5_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_29),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_5_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_617 ? _slots_9_io_out_uop_uopc : _GEN_616 ? _slots_8_io_out_uop_uopc : _GEN_615 ? _slots_7_io_out_uop_uopc : _slots_6_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_617 ? _slots_9_io_out_uop_is_rvc : _GEN_616 ? _slots_8_io_out_uop_is_rvc : _GEN_615 ? _slots_7_io_out_uop_is_rvc : _slots_6_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_617 ? _slots_9_io_out_uop_fu_code : _GEN_616 ? _slots_8_io_out_uop_fu_code : _GEN_615 ? _slots_7_io_out_uop_fu_code : _slots_6_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_617 ? _slots_9_io_out_uop_iw_state : _GEN_616 ? _slots_8_io_out_uop_iw_state : _GEN_615 ? _slots_7_io_out_uop_iw_state : _slots_6_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_617 ? _slots_9_io_out_uop_iw_p1_poisoned : _GEN_616 ? _slots_8_io_out_uop_iw_p1_poisoned : _GEN_615 ? _slots_7_io_out_uop_iw_p1_poisoned : _slots_6_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_617 ? _slots_9_io_out_uop_iw_p2_poisoned : _GEN_616 ? _slots_8_io_out_uop_iw_p2_poisoned : _GEN_615 ? _slots_7_io_out_uop_iw_p2_poisoned : _slots_6_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_617 ? _slots_9_io_out_uop_is_br : _GEN_616 ? _slots_8_io_out_uop_is_br : _GEN_615 ? _slots_7_io_out_uop_is_br : _slots_6_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_617 ? _slots_9_io_out_uop_is_jalr : _GEN_616 ? _slots_8_io_out_uop_is_jalr : _GEN_615 ? _slots_7_io_out_uop_is_jalr : _slots_6_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_617 ? _slots_9_io_out_uop_is_jal : _GEN_616 ? _slots_8_io_out_uop_is_jal : _GEN_615 ? _slots_7_io_out_uop_is_jal : _slots_6_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_617 ? _slots_9_io_out_uop_is_sfb : _GEN_616 ? _slots_8_io_out_uop_is_sfb : _GEN_615 ? _slots_7_io_out_uop_is_sfb : _slots_6_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_617 ? _slots_9_io_out_uop_br_mask : _GEN_616 ? _slots_8_io_out_uop_br_mask : _GEN_615 ? _slots_7_io_out_uop_br_mask : _slots_6_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_617 ? _slots_9_io_out_uop_br_tag : _GEN_616 ? _slots_8_io_out_uop_br_tag : _GEN_615 ? _slots_7_io_out_uop_br_tag : _slots_6_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_617 ? _slots_9_io_out_uop_ftq_idx : _GEN_616 ? _slots_8_io_out_uop_ftq_idx : _GEN_615 ? _slots_7_io_out_uop_ftq_idx : _slots_6_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_617 ? _slots_9_io_out_uop_edge_inst : _GEN_616 ? _slots_8_io_out_uop_edge_inst : _GEN_615 ? _slots_7_io_out_uop_edge_inst : _slots_6_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_617 ? _slots_9_io_out_uop_pc_lob : _GEN_616 ? _slots_8_io_out_uop_pc_lob : _GEN_615 ? _slots_7_io_out_uop_pc_lob : _slots_6_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_617 ? _slots_9_io_out_uop_taken : _GEN_616 ? _slots_8_io_out_uop_taken : _GEN_615 ? _slots_7_io_out_uop_taken : _slots_6_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_617 ? _slots_9_io_out_uop_imm_packed : _GEN_616 ? _slots_8_io_out_uop_imm_packed : _GEN_615 ? _slots_7_io_out_uop_imm_packed : _slots_6_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_617 ? _slots_9_io_out_uop_rob_idx : _GEN_616 ? _slots_8_io_out_uop_rob_idx : _GEN_615 ? _slots_7_io_out_uop_rob_idx : _slots_6_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_617 ? _slots_9_io_out_uop_ldq_idx : _GEN_616 ? _slots_8_io_out_uop_ldq_idx : _GEN_615 ? _slots_7_io_out_uop_ldq_idx : _slots_6_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_617 ? _slots_9_io_out_uop_stq_idx : _GEN_616 ? _slots_8_io_out_uop_stq_idx : _GEN_615 ? _slots_7_io_out_uop_stq_idx : _slots_6_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_617 ? _slots_9_io_out_uop_pdst : _GEN_616 ? _slots_8_io_out_uop_pdst : _GEN_615 ? _slots_7_io_out_uop_pdst : _slots_6_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_617 ? _slots_9_io_out_uop_prs1 : _GEN_616 ? _slots_8_io_out_uop_prs1 : _GEN_615 ? _slots_7_io_out_uop_prs1 : _slots_6_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_617 ? _slots_9_io_out_uop_prs2 : _GEN_616 ? _slots_8_io_out_uop_prs2 : _GEN_615 ? _slots_7_io_out_uop_prs2 : _slots_6_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_617 ? _slots_9_io_out_uop_prs3 : _GEN_616 ? _slots_8_io_out_uop_prs3 : _GEN_615 ? _slots_7_io_out_uop_prs3 : _slots_6_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_617 ? _slots_9_io_out_uop_prs1_busy : _GEN_616 ? _slots_8_io_out_uop_prs1_busy : _GEN_615 ? _slots_7_io_out_uop_prs1_busy : _slots_6_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_617 ? _slots_9_io_out_uop_prs2_busy : _GEN_616 ? _slots_8_io_out_uop_prs2_busy : _GEN_615 ? _slots_7_io_out_uop_prs2_busy : _slots_6_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_617 ? _slots_9_io_out_uop_prs3_busy : _GEN_616 ? _slots_8_io_out_uop_prs3_busy : _GEN_615 ? _slots_7_io_out_uop_prs3_busy : _slots_6_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_617 ? _slots_9_io_out_uop_ppred_busy : _GEN_616 ? _slots_8_io_out_uop_ppred_busy : _GEN_615 ? _slots_7_io_out_uop_ppred_busy : _slots_6_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_617 ? _slots_9_io_out_uop_bypassable : _GEN_616 ? _slots_8_io_out_uop_bypassable : _GEN_615 ? _slots_7_io_out_uop_bypassable : _slots_6_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_617 ? _slots_9_io_out_uop_mem_cmd : _GEN_616 ? _slots_8_io_out_uop_mem_cmd : _GEN_615 ? _slots_7_io_out_uop_mem_cmd : _slots_6_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_617 ? _slots_9_io_out_uop_mem_size : _GEN_616 ? _slots_8_io_out_uop_mem_size : _GEN_615 ? _slots_7_io_out_uop_mem_size : _slots_6_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_617 ? _slots_9_io_out_uop_mem_signed : _GEN_616 ? _slots_8_io_out_uop_mem_signed : _GEN_615 ? _slots_7_io_out_uop_mem_signed : _slots_6_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_617 ? _slots_9_io_out_uop_is_fence : _GEN_616 ? _slots_8_io_out_uop_is_fence : _GEN_615 ? _slots_7_io_out_uop_is_fence : _slots_6_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_617 ? _slots_9_io_out_uop_is_amo : _GEN_616 ? _slots_8_io_out_uop_is_amo : _GEN_615 ? _slots_7_io_out_uop_is_amo : _slots_6_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_617 ? _slots_9_io_out_uop_uses_ldq : _GEN_616 ? _slots_8_io_out_uop_uses_ldq : _GEN_615 ? _slots_7_io_out_uop_uses_ldq : _slots_6_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_617 ? _slots_9_io_out_uop_uses_stq : _GEN_616 ? _slots_8_io_out_uop_uses_stq : _GEN_615 ? _slots_7_io_out_uop_uses_stq : _slots_6_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_617 ? _slots_9_io_out_uop_ldst_val : _GEN_616 ? _slots_8_io_out_uop_ldst_val : _GEN_615 ? _slots_7_io_out_uop_ldst_val : _slots_6_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_617 ? _slots_9_io_out_uop_dst_rtype : _GEN_616 ? _slots_8_io_out_uop_dst_rtype : _GEN_615 ? _slots_7_io_out_uop_dst_rtype : _slots_6_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_617 ? _slots_9_io_out_uop_lrs1_rtype : _GEN_616 ? _slots_8_io_out_uop_lrs1_rtype : _GEN_615 ? _slots_7_io_out_uop_lrs1_rtype : _slots_6_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_617 ? _slots_9_io_out_uop_lrs2_rtype : _GEN_616 ? _slots_8_io_out_uop_lrs2_rtype : _GEN_615 ? _slots_7_io_out_uop_lrs2_rtype : _slots_6_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_617 ? _slots_9_io_out_uop_fp_val : _GEN_616 ? _slots_8_io_out_uop_fp_val : _GEN_615 ? _slots_7_io_out_uop_fp_val : _slots_6_io_out_uop_fp_val),
    .io_valid                       (_slots_5_io_valid),
    .io_will_be_valid               (_slots_5_io_will_be_valid),
    .io_request                     (_slots_5_io_request),
    .io_out_uop_uopc                (_slots_5_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_5_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_5_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_5_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_5_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_5_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_5_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_5_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_5_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_5_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_5_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_5_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_5_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_5_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_5_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_5_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_5_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_5_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_5_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_5_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_5_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_5_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_5_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_5_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_5_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_5_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_5_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_5_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_5_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_5_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_5_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_5_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_5_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_5_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_5_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_5_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_5_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_5_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_5_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_5_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_5_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_5_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_5_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_5_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_5_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_5_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_5_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_5_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_5_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_5_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_5_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_5_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_5_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_5_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_5_io_uop_pc_lob),
    .io_uop_taken                   (_slots_5_io_uop_taken),
    .io_uop_imm_packed              (_slots_5_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_5_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_5_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_5_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_5_io_uop_pdst),
    .io_uop_prs1                    (_slots_5_io_uop_prs1),
    .io_uop_prs2                    (_slots_5_io_uop_prs2),
    .io_uop_bypassable              (_slots_5_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_5_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_5_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_5_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_5_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_5_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_5_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_5_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_5_io_uop_fp_val)
  );
  IssueSlot_32 slots_6 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_6_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_31),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_6_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_620 ? _slots_10_io_out_uop_uopc : _GEN_619 ? _slots_9_io_out_uop_uopc : _GEN_618 ? _slots_8_io_out_uop_uopc : _slots_7_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_620 ? _slots_10_io_out_uop_is_rvc : _GEN_619 ? _slots_9_io_out_uop_is_rvc : _GEN_618 ? _slots_8_io_out_uop_is_rvc : _slots_7_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_620 ? _slots_10_io_out_uop_fu_code : _GEN_619 ? _slots_9_io_out_uop_fu_code : _GEN_618 ? _slots_8_io_out_uop_fu_code : _slots_7_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_620 ? _slots_10_io_out_uop_iw_state : _GEN_619 ? _slots_9_io_out_uop_iw_state : _GEN_618 ? _slots_8_io_out_uop_iw_state : _slots_7_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_620 ? _slots_10_io_out_uop_iw_p1_poisoned : _GEN_619 ? _slots_9_io_out_uop_iw_p1_poisoned : _GEN_618 ? _slots_8_io_out_uop_iw_p1_poisoned : _slots_7_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_620 ? _slots_10_io_out_uop_iw_p2_poisoned : _GEN_619 ? _slots_9_io_out_uop_iw_p2_poisoned : _GEN_618 ? _slots_8_io_out_uop_iw_p2_poisoned : _slots_7_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_620 ? _slots_10_io_out_uop_is_br : _GEN_619 ? _slots_9_io_out_uop_is_br : _GEN_618 ? _slots_8_io_out_uop_is_br : _slots_7_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_620 ? _slots_10_io_out_uop_is_jalr : _GEN_619 ? _slots_9_io_out_uop_is_jalr : _GEN_618 ? _slots_8_io_out_uop_is_jalr : _slots_7_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_620 ? _slots_10_io_out_uop_is_jal : _GEN_619 ? _slots_9_io_out_uop_is_jal : _GEN_618 ? _slots_8_io_out_uop_is_jal : _slots_7_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_620 ? _slots_10_io_out_uop_is_sfb : _GEN_619 ? _slots_9_io_out_uop_is_sfb : _GEN_618 ? _slots_8_io_out_uop_is_sfb : _slots_7_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_620 ? _slots_10_io_out_uop_br_mask : _GEN_619 ? _slots_9_io_out_uop_br_mask : _GEN_618 ? _slots_8_io_out_uop_br_mask : _slots_7_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_620 ? _slots_10_io_out_uop_br_tag : _GEN_619 ? _slots_9_io_out_uop_br_tag : _GEN_618 ? _slots_8_io_out_uop_br_tag : _slots_7_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_620 ? _slots_10_io_out_uop_ftq_idx : _GEN_619 ? _slots_9_io_out_uop_ftq_idx : _GEN_618 ? _slots_8_io_out_uop_ftq_idx : _slots_7_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_620 ? _slots_10_io_out_uop_edge_inst : _GEN_619 ? _slots_9_io_out_uop_edge_inst : _GEN_618 ? _slots_8_io_out_uop_edge_inst : _slots_7_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_620 ? _slots_10_io_out_uop_pc_lob : _GEN_619 ? _slots_9_io_out_uop_pc_lob : _GEN_618 ? _slots_8_io_out_uop_pc_lob : _slots_7_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_620 ? _slots_10_io_out_uop_taken : _GEN_619 ? _slots_9_io_out_uop_taken : _GEN_618 ? _slots_8_io_out_uop_taken : _slots_7_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_620 ? _slots_10_io_out_uop_imm_packed : _GEN_619 ? _slots_9_io_out_uop_imm_packed : _GEN_618 ? _slots_8_io_out_uop_imm_packed : _slots_7_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_620 ? _slots_10_io_out_uop_rob_idx : _GEN_619 ? _slots_9_io_out_uop_rob_idx : _GEN_618 ? _slots_8_io_out_uop_rob_idx : _slots_7_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_620 ? _slots_10_io_out_uop_ldq_idx : _GEN_619 ? _slots_9_io_out_uop_ldq_idx : _GEN_618 ? _slots_8_io_out_uop_ldq_idx : _slots_7_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_620 ? _slots_10_io_out_uop_stq_idx : _GEN_619 ? _slots_9_io_out_uop_stq_idx : _GEN_618 ? _slots_8_io_out_uop_stq_idx : _slots_7_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_620 ? _slots_10_io_out_uop_pdst : _GEN_619 ? _slots_9_io_out_uop_pdst : _GEN_618 ? _slots_8_io_out_uop_pdst : _slots_7_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_620 ? _slots_10_io_out_uop_prs1 : _GEN_619 ? _slots_9_io_out_uop_prs1 : _GEN_618 ? _slots_8_io_out_uop_prs1 : _slots_7_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_620 ? _slots_10_io_out_uop_prs2 : _GEN_619 ? _slots_9_io_out_uop_prs2 : _GEN_618 ? _slots_8_io_out_uop_prs2 : _slots_7_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_620 ? _slots_10_io_out_uop_prs3 : _GEN_619 ? _slots_9_io_out_uop_prs3 : _GEN_618 ? _slots_8_io_out_uop_prs3 : _slots_7_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_620 ? _slots_10_io_out_uop_prs1_busy : _GEN_619 ? _slots_9_io_out_uop_prs1_busy : _GEN_618 ? _slots_8_io_out_uop_prs1_busy : _slots_7_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_620 ? _slots_10_io_out_uop_prs2_busy : _GEN_619 ? _slots_9_io_out_uop_prs2_busy : _GEN_618 ? _slots_8_io_out_uop_prs2_busy : _slots_7_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_620 ? _slots_10_io_out_uop_prs3_busy : _GEN_619 ? _slots_9_io_out_uop_prs3_busy : _GEN_618 ? _slots_8_io_out_uop_prs3_busy : _slots_7_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_620 ? _slots_10_io_out_uop_ppred_busy : _GEN_619 ? _slots_9_io_out_uop_ppred_busy : _GEN_618 ? _slots_8_io_out_uop_ppred_busy : _slots_7_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_620 ? _slots_10_io_out_uop_bypassable : _GEN_619 ? _slots_9_io_out_uop_bypassable : _GEN_618 ? _slots_8_io_out_uop_bypassable : _slots_7_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_620 ? _slots_10_io_out_uop_mem_cmd : _GEN_619 ? _slots_9_io_out_uop_mem_cmd : _GEN_618 ? _slots_8_io_out_uop_mem_cmd : _slots_7_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_620 ? _slots_10_io_out_uop_mem_size : _GEN_619 ? _slots_9_io_out_uop_mem_size : _GEN_618 ? _slots_8_io_out_uop_mem_size : _slots_7_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_620 ? _slots_10_io_out_uop_mem_signed : _GEN_619 ? _slots_9_io_out_uop_mem_signed : _GEN_618 ? _slots_8_io_out_uop_mem_signed : _slots_7_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_620 ? _slots_10_io_out_uop_is_fence : _GEN_619 ? _slots_9_io_out_uop_is_fence : _GEN_618 ? _slots_8_io_out_uop_is_fence : _slots_7_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_620 ? _slots_10_io_out_uop_is_amo : _GEN_619 ? _slots_9_io_out_uop_is_amo : _GEN_618 ? _slots_8_io_out_uop_is_amo : _slots_7_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_620 ? _slots_10_io_out_uop_uses_ldq : _GEN_619 ? _slots_9_io_out_uop_uses_ldq : _GEN_618 ? _slots_8_io_out_uop_uses_ldq : _slots_7_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_620 ? _slots_10_io_out_uop_uses_stq : _GEN_619 ? _slots_9_io_out_uop_uses_stq : _GEN_618 ? _slots_8_io_out_uop_uses_stq : _slots_7_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_620 ? _slots_10_io_out_uop_ldst_val : _GEN_619 ? _slots_9_io_out_uop_ldst_val : _GEN_618 ? _slots_8_io_out_uop_ldst_val : _slots_7_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_620 ? _slots_10_io_out_uop_dst_rtype : _GEN_619 ? _slots_9_io_out_uop_dst_rtype : _GEN_618 ? _slots_8_io_out_uop_dst_rtype : _slots_7_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_620 ? _slots_10_io_out_uop_lrs1_rtype : _GEN_619 ? _slots_9_io_out_uop_lrs1_rtype : _GEN_618 ? _slots_8_io_out_uop_lrs1_rtype : _slots_7_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_620 ? _slots_10_io_out_uop_lrs2_rtype : _GEN_619 ? _slots_9_io_out_uop_lrs2_rtype : _GEN_618 ? _slots_8_io_out_uop_lrs2_rtype : _slots_7_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_620 ? _slots_10_io_out_uop_fp_val : _GEN_619 ? _slots_9_io_out_uop_fp_val : _GEN_618 ? _slots_8_io_out_uop_fp_val : _slots_7_io_out_uop_fp_val),
    .io_valid                       (_slots_6_io_valid),
    .io_will_be_valid               (_slots_6_io_will_be_valid),
    .io_request                     (_slots_6_io_request),
    .io_out_uop_uopc                (_slots_6_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_6_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_6_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_6_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_6_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_6_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_6_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_6_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_6_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_6_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_6_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_6_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_6_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_6_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_6_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_6_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_6_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_6_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_6_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_6_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_6_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_6_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_6_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_6_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_6_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_6_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_6_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_6_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_6_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_6_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_6_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_6_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_6_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_6_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_6_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_6_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_6_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_6_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_6_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_6_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_6_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_6_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_6_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_6_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_6_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_6_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_6_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_6_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_6_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_6_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_6_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_6_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_6_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_6_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_6_io_uop_pc_lob),
    .io_uop_taken                   (_slots_6_io_uop_taken),
    .io_uop_imm_packed              (_slots_6_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_6_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_6_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_6_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_6_io_uop_pdst),
    .io_uop_prs1                    (_slots_6_io_uop_prs1),
    .io_uop_prs2                    (_slots_6_io_uop_prs2),
    .io_uop_bypassable              (_slots_6_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_6_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_6_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_6_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_6_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_6_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_6_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_6_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_6_io_uop_fp_val)
  );
  IssueSlot_32 slots_7 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_7_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_33),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_7_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_623 ? _slots_11_io_out_uop_uopc : _GEN_622 ? _slots_10_io_out_uop_uopc : _GEN_621 ? _slots_9_io_out_uop_uopc : _slots_8_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_623 ? _slots_11_io_out_uop_is_rvc : _GEN_622 ? _slots_10_io_out_uop_is_rvc : _GEN_621 ? _slots_9_io_out_uop_is_rvc : _slots_8_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_623 ? _slots_11_io_out_uop_fu_code : _GEN_622 ? _slots_10_io_out_uop_fu_code : _GEN_621 ? _slots_9_io_out_uop_fu_code : _slots_8_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_623 ? _slots_11_io_out_uop_iw_state : _GEN_622 ? _slots_10_io_out_uop_iw_state : _GEN_621 ? _slots_9_io_out_uop_iw_state : _slots_8_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_623 ? _slots_11_io_out_uop_iw_p1_poisoned : _GEN_622 ? _slots_10_io_out_uop_iw_p1_poisoned : _GEN_621 ? _slots_9_io_out_uop_iw_p1_poisoned : _slots_8_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_623 ? _slots_11_io_out_uop_iw_p2_poisoned : _GEN_622 ? _slots_10_io_out_uop_iw_p2_poisoned : _GEN_621 ? _slots_9_io_out_uop_iw_p2_poisoned : _slots_8_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_623 ? _slots_11_io_out_uop_is_br : _GEN_622 ? _slots_10_io_out_uop_is_br : _GEN_621 ? _slots_9_io_out_uop_is_br : _slots_8_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_623 ? _slots_11_io_out_uop_is_jalr : _GEN_622 ? _slots_10_io_out_uop_is_jalr : _GEN_621 ? _slots_9_io_out_uop_is_jalr : _slots_8_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_623 ? _slots_11_io_out_uop_is_jal : _GEN_622 ? _slots_10_io_out_uop_is_jal : _GEN_621 ? _slots_9_io_out_uop_is_jal : _slots_8_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_623 ? _slots_11_io_out_uop_is_sfb : _GEN_622 ? _slots_10_io_out_uop_is_sfb : _GEN_621 ? _slots_9_io_out_uop_is_sfb : _slots_8_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_623 ? _slots_11_io_out_uop_br_mask : _GEN_622 ? _slots_10_io_out_uop_br_mask : _GEN_621 ? _slots_9_io_out_uop_br_mask : _slots_8_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_623 ? _slots_11_io_out_uop_br_tag : _GEN_622 ? _slots_10_io_out_uop_br_tag : _GEN_621 ? _slots_9_io_out_uop_br_tag : _slots_8_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_623 ? _slots_11_io_out_uop_ftq_idx : _GEN_622 ? _slots_10_io_out_uop_ftq_idx : _GEN_621 ? _slots_9_io_out_uop_ftq_idx : _slots_8_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_623 ? _slots_11_io_out_uop_edge_inst : _GEN_622 ? _slots_10_io_out_uop_edge_inst : _GEN_621 ? _slots_9_io_out_uop_edge_inst : _slots_8_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_623 ? _slots_11_io_out_uop_pc_lob : _GEN_622 ? _slots_10_io_out_uop_pc_lob : _GEN_621 ? _slots_9_io_out_uop_pc_lob : _slots_8_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_623 ? _slots_11_io_out_uop_taken : _GEN_622 ? _slots_10_io_out_uop_taken : _GEN_621 ? _slots_9_io_out_uop_taken : _slots_8_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_623 ? _slots_11_io_out_uop_imm_packed : _GEN_622 ? _slots_10_io_out_uop_imm_packed : _GEN_621 ? _slots_9_io_out_uop_imm_packed : _slots_8_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_623 ? _slots_11_io_out_uop_rob_idx : _GEN_622 ? _slots_10_io_out_uop_rob_idx : _GEN_621 ? _slots_9_io_out_uop_rob_idx : _slots_8_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_623 ? _slots_11_io_out_uop_ldq_idx : _GEN_622 ? _slots_10_io_out_uop_ldq_idx : _GEN_621 ? _slots_9_io_out_uop_ldq_idx : _slots_8_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_623 ? _slots_11_io_out_uop_stq_idx : _GEN_622 ? _slots_10_io_out_uop_stq_idx : _GEN_621 ? _slots_9_io_out_uop_stq_idx : _slots_8_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_623 ? _slots_11_io_out_uop_pdst : _GEN_622 ? _slots_10_io_out_uop_pdst : _GEN_621 ? _slots_9_io_out_uop_pdst : _slots_8_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_623 ? _slots_11_io_out_uop_prs1 : _GEN_622 ? _slots_10_io_out_uop_prs1 : _GEN_621 ? _slots_9_io_out_uop_prs1 : _slots_8_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_623 ? _slots_11_io_out_uop_prs2 : _GEN_622 ? _slots_10_io_out_uop_prs2 : _GEN_621 ? _slots_9_io_out_uop_prs2 : _slots_8_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_623 ? _slots_11_io_out_uop_prs3 : _GEN_622 ? _slots_10_io_out_uop_prs3 : _GEN_621 ? _slots_9_io_out_uop_prs3 : _slots_8_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_623 ? _slots_11_io_out_uop_prs1_busy : _GEN_622 ? _slots_10_io_out_uop_prs1_busy : _GEN_621 ? _slots_9_io_out_uop_prs1_busy : _slots_8_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_623 ? _slots_11_io_out_uop_prs2_busy : _GEN_622 ? _slots_10_io_out_uop_prs2_busy : _GEN_621 ? _slots_9_io_out_uop_prs2_busy : _slots_8_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_623 ? _slots_11_io_out_uop_prs3_busy : _GEN_622 ? _slots_10_io_out_uop_prs3_busy : _GEN_621 ? _slots_9_io_out_uop_prs3_busy : _slots_8_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_623 ? _slots_11_io_out_uop_ppred_busy : _GEN_622 ? _slots_10_io_out_uop_ppred_busy : _GEN_621 ? _slots_9_io_out_uop_ppred_busy : _slots_8_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_623 ? _slots_11_io_out_uop_bypassable : _GEN_622 ? _slots_10_io_out_uop_bypassable : _GEN_621 ? _slots_9_io_out_uop_bypassable : _slots_8_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_623 ? _slots_11_io_out_uop_mem_cmd : _GEN_622 ? _slots_10_io_out_uop_mem_cmd : _GEN_621 ? _slots_9_io_out_uop_mem_cmd : _slots_8_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_623 ? _slots_11_io_out_uop_mem_size : _GEN_622 ? _slots_10_io_out_uop_mem_size : _GEN_621 ? _slots_9_io_out_uop_mem_size : _slots_8_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_623 ? _slots_11_io_out_uop_mem_signed : _GEN_622 ? _slots_10_io_out_uop_mem_signed : _GEN_621 ? _slots_9_io_out_uop_mem_signed : _slots_8_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_623 ? _slots_11_io_out_uop_is_fence : _GEN_622 ? _slots_10_io_out_uop_is_fence : _GEN_621 ? _slots_9_io_out_uop_is_fence : _slots_8_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_623 ? _slots_11_io_out_uop_is_amo : _GEN_622 ? _slots_10_io_out_uop_is_amo : _GEN_621 ? _slots_9_io_out_uop_is_amo : _slots_8_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_623 ? _slots_11_io_out_uop_uses_ldq : _GEN_622 ? _slots_10_io_out_uop_uses_ldq : _GEN_621 ? _slots_9_io_out_uop_uses_ldq : _slots_8_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_623 ? _slots_11_io_out_uop_uses_stq : _GEN_622 ? _slots_10_io_out_uop_uses_stq : _GEN_621 ? _slots_9_io_out_uop_uses_stq : _slots_8_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_623 ? _slots_11_io_out_uop_ldst_val : _GEN_622 ? _slots_10_io_out_uop_ldst_val : _GEN_621 ? _slots_9_io_out_uop_ldst_val : _slots_8_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_623 ? _slots_11_io_out_uop_dst_rtype : _GEN_622 ? _slots_10_io_out_uop_dst_rtype : _GEN_621 ? _slots_9_io_out_uop_dst_rtype : _slots_8_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_623 ? _slots_11_io_out_uop_lrs1_rtype : _GEN_622 ? _slots_10_io_out_uop_lrs1_rtype : _GEN_621 ? _slots_9_io_out_uop_lrs1_rtype : _slots_8_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_623 ? _slots_11_io_out_uop_lrs2_rtype : _GEN_622 ? _slots_10_io_out_uop_lrs2_rtype : _GEN_621 ? _slots_9_io_out_uop_lrs2_rtype : _slots_8_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_623 ? _slots_11_io_out_uop_fp_val : _GEN_622 ? _slots_10_io_out_uop_fp_val : _GEN_621 ? _slots_9_io_out_uop_fp_val : _slots_8_io_out_uop_fp_val),
    .io_valid                       (_slots_7_io_valid),
    .io_will_be_valid               (_slots_7_io_will_be_valid),
    .io_request                     (_slots_7_io_request),
    .io_out_uop_uopc                (_slots_7_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_7_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_7_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_7_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_7_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_7_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_7_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_7_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_7_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_7_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_7_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_7_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_7_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_7_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_7_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_7_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_7_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_7_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_7_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_7_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_7_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_7_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_7_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_7_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_7_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_7_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_7_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_7_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_7_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_7_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_7_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_7_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_7_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_7_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_7_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_7_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_7_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_7_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_7_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_7_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_7_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_7_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_7_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_7_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_7_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_7_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_7_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_7_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_7_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_7_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_7_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_7_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_7_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_7_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_7_io_uop_pc_lob),
    .io_uop_taken                   (_slots_7_io_uop_taken),
    .io_uop_imm_packed              (_slots_7_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_7_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_7_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_7_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_7_io_uop_pdst),
    .io_uop_prs1                    (_slots_7_io_uop_prs1),
    .io_uop_prs2                    (_slots_7_io_uop_prs2),
    .io_uop_bypassable              (_slots_7_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_7_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_7_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_7_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_7_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_7_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_7_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_7_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_7_io_uop_fp_val)
  );
  IssueSlot_32 slots_8 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_8_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_35),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_8_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_626 ? _slots_12_io_out_uop_uopc : _GEN_625 ? _slots_11_io_out_uop_uopc : _GEN_624 ? _slots_10_io_out_uop_uopc : _slots_9_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_626 ? _slots_12_io_out_uop_is_rvc : _GEN_625 ? _slots_11_io_out_uop_is_rvc : _GEN_624 ? _slots_10_io_out_uop_is_rvc : _slots_9_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_626 ? _slots_12_io_out_uop_fu_code : _GEN_625 ? _slots_11_io_out_uop_fu_code : _GEN_624 ? _slots_10_io_out_uop_fu_code : _slots_9_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_626 ? _slots_12_io_out_uop_iw_state : _GEN_625 ? _slots_11_io_out_uop_iw_state : _GEN_624 ? _slots_10_io_out_uop_iw_state : _slots_9_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_626 ? _slots_12_io_out_uop_iw_p1_poisoned : _GEN_625 ? _slots_11_io_out_uop_iw_p1_poisoned : _GEN_624 ? _slots_10_io_out_uop_iw_p1_poisoned : _slots_9_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_626 ? _slots_12_io_out_uop_iw_p2_poisoned : _GEN_625 ? _slots_11_io_out_uop_iw_p2_poisoned : _GEN_624 ? _slots_10_io_out_uop_iw_p2_poisoned : _slots_9_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_626 ? _slots_12_io_out_uop_is_br : _GEN_625 ? _slots_11_io_out_uop_is_br : _GEN_624 ? _slots_10_io_out_uop_is_br : _slots_9_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_626 ? _slots_12_io_out_uop_is_jalr : _GEN_625 ? _slots_11_io_out_uop_is_jalr : _GEN_624 ? _slots_10_io_out_uop_is_jalr : _slots_9_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_626 ? _slots_12_io_out_uop_is_jal : _GEN_625 ? _slots_11_io_out_uop_is_jal : _GEN_624 ? _slots_10_io_out_uop_is_jal : _slots_9_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_626 ? _slots_12_io_out_uop_is_sfb : _GEN_625 ? _slots_11_io_out_uop_is_sfb : _GEN_624 ? _slots_10_io_out_uop_is_sfb : _slots_9_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_626 ? _slots_12_io_out_uop_br_mask : _GEN_625 ? _slots_11_io_out_uop_br_mask : _GEN_624 ? _slots_10_io_out_uop_br_mask : _slots_9_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_626 ? _slots_12_io_out_uop_br_tag : _GEN_625 ? _slots_11_io_out_uop_br_tag : _GEN_624 ? _slots_10_io_out_uop_br_tag : _slots_9_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_626 ? _slots_12_io_out_uop_ftq_idx : _GEN_625 ? _slots_11_io_out_uop_ftq_idx : _GEN_624 ? _slots_10_io_out_uop_ftq_idx : _slots_9_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_626 ? _slots_12_io_out_uop_edge_inst : _GEN_625 ? _slots_11_io_out_uop_edge_inst : _GEN_624 ? _slots_10_io_out_uop_edge_inst : _slots_9_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_626 ? _slots_12_io_out_uop_pc_lob : _GEN_625 ? _slots_11_io_out_uop_pc_lob : _GEN_624 ? _slots_10_io_out_uop_pc_lob : _slots_9_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_626 ? _slots_12_io_out_uop_taken : _GEN_625 ? _slots_11_io_out_uop_taken : _GEN_624 ? _slots_10_io_out_uop_taken : _slots_9_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_626 ? _slots_12_io_out_uop_imm_packed : _GEN_625 ? _slots_11_io_out_uop_imm_packed : _GEN_624 ? _slots_10_io_out_uop_imm_packed : _slots_9_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_626 ? _slots_12_io_out_uop_rob_idx : _GEN_625 ? _slots_11_io_out_uop_rob_idx : _GEN_624 ? _slots_10_io_out_uop_rob_idx : _slots_9_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_626 ? _slots_12_io_out_uop_ldq_idx : _GEN_625 ? _slots_11_io_out_uop_ldq_idx : _GEN_624 ? _slots_10_io_out_uop_ldq_idx : _slots_9_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_626 ? _slots_12_io_out_uop_stq_idx : _GEN_625 ? _slots_11_io_out_uop_stq_idx : _GEN_624 ? _slots_10_io_out_uop_stq_idx : _slots_9_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_626 ? _slots_12_io_out_uop_pdst : _GEN_625 ? _slots_11_io_out_uop_pdst : _GEN_624 ? _slots_10_io_out_uop_pdst : _slots_9_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_626 ? _slots_12_io_out_uop_prs1 : _GEN_625 ? _slots_11_io_out_uop_prs1 : _GEN_624 ? _slots_10_io_out_uop_prs1 : _slots_9_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_626 ? _slots_12_io_out_uop_prs2 : _GEN_625 ? _slots_11_io_out_uop_prs2 : _GEN_624 ? _slots_10_io_out_uop_prs2 : _slots_9_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_626 ? _slots_12_io_out_uop_prs3 : _GEN_625 ? _slots_11_io_out_uop_prs3 : _GEN_624 ? _slots_10_io_out_uop_prs3 : _slots_9_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_626 ? _slots_12_io_out_uop_prs1_busy : _GEN_625 ? _slots_11_io_out_uop_prs1_busy : _GEN_624 ? _slots_10_io_out_uop_prs1_busy : _slots_9_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_626 ? _slots_12_io_out_uop_prs2_busy : _GEN_625 ? _slots_11_io_out_uop_prs2_busy : _GEN_624 ? _slots_10_io_out_uop_prs2_busy : _slots_9_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_626 ? _slots_12_io_out_uop_prs3_busy : _GEN_625 ? _slots_11_io_out_uop_prs3_busy : _GEN_624 ? _slots_10_io_out_uop_prs3_busy : _slots_9_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_626 ? _slots_12_io_out_uop_ppred_busy : _GEN_625 ? _slots_11_io_out_uop_ppred_busy : _GEN_624 ? _slots_10_io_out_uop_ppred_busy : _slots_9_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_626 ? _slots_12_io_out_uop_bypassable : _GEN_625 ? _slots_11_io_out_uop_bypassable : _GEN_624 ? _slots_10_io_out_uop_bypassable : _slots_9_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_626 ? _slots_12_io_out_uop_mem_cmd : _GEN_625 ? _slots_11_io_out_uop_mem_cmd : _GEN_624 ? _slots_10_io_out_uop_mem_cmd : _slots_9_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_626 ? _slots_12_io_out_uop_mem_size : _GEN_625 ? _slots_11_io_out_uop_mem_size : _GEN_624 ? _slots_10_io_out_uop_mem_size : _slots_9_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_626 ? _slots_12_io_out_uop_mem_signed : _GEN_625 ? _slots_11_io_out_uop_mem_signed : _GEN_624 ? _slots_10_io_out_uop_mem_signed : _slots_9_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_626 ? _slots_12_io_out_uop_is_fence : _GEN_625 ? _slots_11_io_out_uop_is_fence : _GEN_624 ? _slots_10_io_out_uop_is_fence : _slots_9_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_626 ? _slots_12_io_out_uop_is_amo : _GEN_625 ? _slots_11_io_out_uop_is_amo : _GEN_624 ? _slots_10_io_out_uop_is_amo : _slots_9_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_626 ? _slots_12_io_out_uop_uses_ldq : _GEN_625 ? _slots_11_io_out_uop_uses_ldq : _GEN_624 ? _slots_10_io_out_uop_uses_ldq : _slots_9_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_626 ? _slots_12_io_out_uop_uses_stq : _GEN_625 ? _slots_11_io_out_uop_uses_stq : _GEN_624 ? _slots_10_io_out_uop_uses_stq : _slots_9_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_626 ? _slots_12_io_out_uop_ldst_val : _GEN_625 ? _slots_11_io_out_uop_ldst_val : _GEN_624 ? _slots_10_io_out_uop_ldst_val : _slots_9_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_626 ? _slots_12_io_out_uop_dst_rtype : _GEN_625 ? _slots_11_io_out_uop_dst_rtype : _GEN_624 ? _slots_10_io_out_uop_dst_rtype : _slots_9_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_626 ? _slots_12_io_out_uop_lrs1_rtype : _GEN_625 ? _slots_11_io_out_uop_lrs1_rtype : _GEN_624 ? _slots_10_io_out_uop_lrs1_rtype : _slots_9_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_626 ? _slots_12_io_out_uop_lrs2_rtype : _GEN_625 ? _slots_11_io_out_uop_lrs2_rtype : _GEN_624 ? _slots_10_io_out_uop_lrs2_rtype : _slots_9_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_626 ? _slots_12_io_out_uop_fp_val : _GEN_625 ? _slots_11_io_out_uop_fp_val : _GEN_624 ? _slots_10_io_out_uop_fp_val : _slots_9_io_out_uop_fp_val),
    .io_valid                       (_slots_8_io_valid),
    .io_will_be_valid               (_slots_8_io_will_be_valid),
    .io_request                     (_slots_8_io_request),
    .io_out_uop_uopc                (_slots_8_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_8_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_8_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_8_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_8_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_8_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_8_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_8_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_8_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_8_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_8_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_8_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_8_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_8_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_8_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_8_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_8_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_8_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_8_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_8_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_8_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_8_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_8_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_8_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_8_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_8_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_8_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_8_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_8_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_8_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_8_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_8_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_8_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_8_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_8_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_8_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_8_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_8_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_8_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_8_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_8_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_8_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_8_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_8_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_8_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_8_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_8_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_8_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_8_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_8_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_8_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_8_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_8_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_8_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_8_io_uop_pc_lob),
    .io_uop_taken                   (_slots_8_io_uop_taken),
    .io_uop_imm_packed              (_slots_8_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_8_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_8_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_8_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_8_io_uop_pdst),
    .io_uop_prs1                    (_slots_8_io_uop_prs1),
    .io_uop_prs2                    (_slots_8_io_uop_prs2),
    .io_uop_bypassable              (_slots_8_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_8_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_8_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_8_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_8_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_8_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_8_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_8_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_8_io_uop_fp_val)
  );
  IssueSlot_32 slots_9 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_9_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_37),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_9_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_629 ? _slots_13_io_out_uop_uopc : _GEN_628 ? _slots_12_io_out_uop_uopc : _GEN_627 ? _slots_11_io_out_uop_uopc : _slots_10_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_629 ? _slots_13_io_out_uop_is_rvc : _GEN_628 ? _slots_12_io_out_uop_is_rvc : _GEN_627 ? _slots_11_io_out_uop_is_rvc : _slots_10_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_629 ? _slots_13_io_out_uop_fu_code : _GEN_628 ? _slots_12_io_out_uop_fu_code : _GEN_627 ? _slots_11_io_out_uop_fu_code : _slots_10_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_629 ? _slots_13_io_out_uop_iw_state : _GEN_628 ? _slots_12_io_out_uop_iw_state : _GEN_627 ? _slots_11_io_out_uop_iw_state : _slots_10_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_629 ? _slots_13_io_out_uop_iw_p1_poisoned : _GEN_628 ? _slots_12_io_out_uop_iw_p1_poisoned : _GEN_627 ? _slots_11_io_out_uop_iw_p1_poisoned : _slots_10_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_629 ? _slots_13_io_out_uop_iw_p2_poisoned : _GEN_628 ? _slots_12_io_out_uop_iw_p2_poisoned : _GEN_627 ? _slots_11_io_out_uop_iw_p2_poisoned : _slots_10_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_629 ? _slots_13_io_out_uop_is_br : _GEN_628 ? _slots_12_io_out_uop_is_br : _GEN_627 ? _slots_11_io_out_uop_is_br : _slots_10_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_629 ? _slots_13_io_out_uop_is_jalr : _GEN_628 ? _slots_12_io_out_uop_is_jalr : _GEN_627 ? _slots_11_io_out_uop_is_jalr : _slots_10_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_629 ? _slots_13_io_out_uop_is_jal : _GEN_628 ? _slots_12_io_out_uop_is_jal : _GEN_627 ? _slots_11_io_out_uop_is_jal : _slots_10_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_629 ? _slots_13_io_out_uop_is_sfb : _GEN_628 ? _slots_12_io_out_uop_is_sfb : _GEN_627 ? _slots_11_io_out_uop_is_sfb : _slots_10_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_629 ? _slots_13_io_out_uop_br_mask : _GEN_628 ? _slots_12_io_out_uop_br_mask : _GEN_627 ? _slots_11_io_out_uop_br_mask : _slots_10_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_629 ? _slots_13_io_out_uop_br_tag : _GEN_628 ? _slots_12_io_out_uop_br_tag : _GEN_627 ? _slots_11_io_out_uop_br_tag : _slots_10_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_629 ? _slots_13_io_out_uop_ftq_idx : _GEN_628 ? _slots_12_io_out_uop_ftq_idx : _GEN_627 ? _slots_11_io_out_uop_ftq_idx : _slots_10_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_629 ? _slots_13_io_out_uop_edge_inst : _GEN_628 ? _slots_12_io_out_uop_edge_inst : _GEN_627 ? _slots_11_io_out_uop_edge_inst : _slots_10_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_629 ? _slots_13_io_out_uop_pc_lob : _GEN_628 ? _slots_12_io_out_uop_pc_lob : _GEN_627 ? _slots_11_io_out_uop_pc_lob : _slots_10_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_629 ? _slots_13_io_out_uop_taken : _GEN_628 ? _slots_12_io_out_uop_taken : _GEN_627 ? _slots_11_io_out_uop_taken : _slots_10_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_629 ? _slots_13_io_out_uop_imm_packed : _GEN_628 ? _slots_12_io_out_uop_imm_packed : _GEN_627 ? _slots_11_io_out_uop_imm_packed : _slots_10_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_629 ? _slots_13_io_out_uop_rob_idx : _GEN_628 ? _slots_12_io_out_uop_rob_idx : _GEN_627 ? _slots_11_io_out_uop_rob_idx : _slots_10_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_629 ? _slots_13_io_out_uop_ldq_idx : _GEN_628 ? _slots_12_io_out_uop_ldq_idx : _GEN_627 ? _slots_11_io_out_uop_ldq_idx : _slots_10_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_629 ? _slots_13_io_out_uop_stq_idx : _GEN_628 ? _slots_12_io_out_uop_stq_idx : _GEN_627 ? _slots_11_io_out_uop_stq_idx : _slots_10_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_629 ? _slots_13_io_out_uop_pdst : _GEN_628 ? _slots_12_io_out_uop_pdst : _GEN_627 ? _slots_11_io_out_uop_pdst : _slots_10_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_629 ? _slots_13_io_out_uop_prs1 : _GEN_628 ? _slots_12_io_out_uop_prs1 : _GEN_627 ? _slots_11_io_out_uop_prs1 : _slots_10_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_629 ? _slots_13_io_out_uop_prs2 : _GEN_628 ? _slots_12_io_out_uop_prs2 : _GEN_627 ? _slots_11_io_out_uop_prs2 : _slots_10_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_629 ? _slots_13_io_out_uop_prs3 : _GEN_628 ? _slots_12_io_out_uop_prs3 : _GEN_627 ? _slots_11_io_out_uop_prs3 : _slots_10_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_629 ? _slots_13_io_out_uop_prs1_busy : _GEN_628 ? _slots_12_io_out_uop_prs1_busy : _GEN_627 ? _slots_11_io_out_uop_prs1_busy : _slots_10_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_629 ? _slots_13_io_out_uop_prs2_busy : _GEN_628 ? _slots_12_io_out_uop_prs2_busy : _GEN_627 ? _slots_11_io_out_uop_prs2_busy : _slots_10_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_629 ? _slots_13_io_out_uop_prs3_busy : _GEN_628 ? _slots_12_io_out_uop_prs3_busy : _GEN_627 ? _slots_11_io_out_uop_prs3_busy : _slots_10_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_629 ? _slots_13_io_out_uop_ppred_busy : _GEN_628 ? _slots_12_io_out_uop_ppred_busy : _GEN_627 ? _slots_11_io_out_uop_ppred_busy : _slots_10_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_629 ? _slots_13_io_out_uop_bypassable : _GEN_628 ? _slots_12_io_out_uop_bypassable : _GEN_627 ? _slots_11_io_out_uop_bypassable : _slots_10_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_629 ? _slots_13_io_out_uop_mem_cmd : _GEN_628 ? _slots_12_io_out_uop_mem_cmd : _GEN_627 ? _slots_11_io_out_uop_mem_cmd : _slots_10_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_629 ? _slots_13_io_out_uop_mem_size : _GEN_628 ? _slots_12_io_out_uop_mem_size : _GEN_627 ? _slots_11_io_out_uop_mem_size : _slots_10_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_629 ? _slots_13_io_out_uop_mem_signed : _GEN_628 ? _slots_12_io_out_uop_mem_signed : _GEN_627 ? _slots_11_io_out_uop_mem_signed : _slots_10_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_629 ? _slots_13_io_out_uop_is_fence : _GEN_628 ? _slots_12_io_out_uop_is_fence : _GEN_627 ? _slots_11_io_out_uop_is_fence : _slots_10_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_629 ? _slots_13_io_out_uop_is_amo : _GEN_628 ? _slots_12_io_out_uop_is_amo : _GEN_627 ? _slots_11_io_out_uop_is_amo : _slots_10_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_629 ? _slots_13_io_out_uop_uses_ldq : _GEN_628 ? _slots_12_io_out_uop_uses_ldq : _GEN_627 ? _slots_11_io_out_uop_uses_ldq : _slots_10_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_629 ? _slots_13_io_out_uop_uses_stq : _GEN_628 ? _slots_12_io_out_uop_uses_stq : _GEN_627 ? _slots_11_io_out_uop_uses_stq : _slots_10_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_629 ? _slots_13_io_out_uop_ldst_val : _GEN_628 ? _slots_12_io_out_uop_ldst_val : _GEN_627 ? _slots_11_io_out_uop_ldst_val : _slots_10_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_629 ? _slots_13_io_out_uop_dst_rtype : _GEN_628 ? _slots_12_io_out_uop_dst_rtype : _GEN_627 ? _slots_11_io_out_uop_dst_rtype : _slots_10_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_629 ? _slots_13_io_out_uop_lrs1_rtype : _GEN_628 ? _slots_12_io_out_uop_lrs1_rtype : _GEN_627 ? _slots_11_io_out_uop_lrs1_rtype : _slots_10_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_629 ? _slots_13_io_out_uop_lrs2_rtype : _GEN_628 ? _slots_12_io_out_uop_lrs2_rtype : _GEN_627 ? _slots_11_io_out_uop_lrs2_rtype : _slots_10_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_629 ? _slots_13_io_out_uop_fp_val : _GEN_628 ? _slots_12_io_out_uop_fp_val : _GEN_627 ? _slots_11_io_out_uop_fp_val : _slots_10_io_out_uop_fp_val),
    .io_valid                       (_slots_9_io_valid),
    .io_will_be_valid               (_slots_9_io_will_be_valid),
    .io_request                     (_slots_9_io_request),
    .io_out_uop_uopc                (_slots_9_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_9_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_9_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_9_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_9_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_9_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_9_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_9_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_9_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_9_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_9_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_9_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_9_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_9_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_9_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_9_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_9_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_9_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_9_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_9_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_9_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_9_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_9_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_9_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_9_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_9_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_9_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_9_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_9_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_9_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_9_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_9_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_9_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_9_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_9_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_9_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_9_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_9_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_9_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_9_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_9_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_9_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_9_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_9_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_9_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_9_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_9_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_9_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_9_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_9_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_9_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_9_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_9_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_9_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_9_io_uop_pc_lob),
    .io_uop_taken                   (_slots_9_io_uop_taken),
    .io_uop_imm_packed              (_slots_9_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_9_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_9_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_9_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_9_io_uop_pdst),
    .io_uop_prs1                    (_slots_9_io_uop_prs1),
    .io_uop_prs2                    (_slots_9_io_uop_prs2),
    .io_uop_bypassable              (_slots_9_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_9_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_9_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_9_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_9_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_9_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_9_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_9_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_9_io_uop_fp_val)
  );
  IssueSlot_32 slots_10 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_10_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_39),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_10_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_632 ? _slots_14_io_out_uop_uopc : _GEN_631 ? _slots_13_io_out_uop_uopc : _GEN_630 ? _slots_12_io_out_uop_uopc : _slots_11_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_632 ? _slots_14_io_out_uop_is_rvc : _GEN_631 ? _slots_13_io_out_uop_is_rvc : _GEN_630 ? _slots_12_io_out_uop_is_rvc : _slots_11_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_632 ? _slots_14_io_out_uop_fu_code : _GEN_631 ? _slots_13_io_out_uop_fu_code : _GEN_630 ? _slots_12_io_out_uop_fu_code : _slots_11_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_632 ? _slots_14_io_out_uop_iw_state : _GEN_631 ? _slots_13_io_out_uop_iw_state : _GEN_630 ? _slots_12_io_out_uop_iw_state : _slots_11_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_632 ? _slots_14_io_out_uop_iw_p1_poisoned : _GEN_631 ? _slots_13_io_out_uop_iw_p1_poisoned : _GEN_630 ? _slots_12_io_out_uop_iw_p1_poisoned : _slots_11_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_632 ? _slots_14_io_out_uop_iw_p2_poisoned : _GEN_631 ? _slots_13_io_out_uop_iw_p2_poisoned : _GEN_630 ? _slots_12_io_out_uop_iw_p2_poisoned : _slots_11_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_632 ? _slots_14_io_out_uop_is_br : _GEN_631 ? _slots_13_io_out_uop_is_br : _GEN_630 ? _slots_12_io_out_uop_is_br : _slots_11_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_632 ? _slots_14_io_out_uop_is_jalr : _GEN_631 ? _slots_13_io_out_uop_is_jalr : _GEN_630 ? _slots_12_io_out_uop_is_jalr : _slots_11_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_632 ? _slots_14_io_out_uop_is_jal : _GEN_631 ? _slots_13_io_out_uop_is_jal : _GEN_630 ? _slots_12_io_out_uop_is_jal : _slots_11_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_632 ? _slots_14_io_out_uop_is_sfb : _GEN_631 ? _slots_13_io_out_uop_is_sfb : _GEN_630 ? _slots_12_io_out_uop_is_sfb : _slots_11_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_632 ? _slots_14_io_out_uop_br_mask : _GEN_631 ? _slots_13_io_out_uop_br_mask : _GEN_630 ? _slots_12_io_out_uop_br_mask : _slots_11_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_632 ? _slots_14_io_out_uop_br_tag : _GEN_631 ? _slots_13_io_out_uop_br_tag : _GEN_630 ? _slots_12_io_out_uop_br_tag : _slots_11_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_632 ? _slots_14_io_out_uop_ftq_idx : _GEN_631 ? _slots_13_io_out_uop_ftq_idx : _GEN_630 ? _slots_12_io_out_uop_ftq_idx : _slots_11_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_632 ? _slots_14_io_out_uop_edge_inst : _GEN_631 ? _slots_13_io_out_uop_edge_inst : _GEN_630 ? _slots_12_io_out_uop_edge_inst : _slots_11_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_632 ? _slots_14_io_out_uop_pc_lob : _GEN_631 ? _slots_13_io_out_uop_pc_lob : _GEN_630 ? _slots_12_io_out_uop_pc_lob : _slots_11_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_632 ? _slots_14_io_out_uop_taken : _GEN_631 ? _slots_13_io_out_uop_taken : _GEN_630 ? _slots_12_io_out_uop_taken : _slots_11_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_632 ? _slots_14_io_out_uop_imm_packed : _GEN_631 ? _slots_13_io_out_uop_imm_packed : _GEN_630 ? _slots_12_io_out_uop_imm_packed : _slots_11_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_632 ? _slots_14_io_out_uop_rob_idx : _GEN_631 ? _slots_13_io_out_uop_rob_idx : _GEN_630 ? _slots_12_io_out_uop_rob_idx : _slots_11_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_632 ? _slots_14_io_out_uop_ldq_idx : _GEN_631 ? _slots_13_io_out_uop_ldq_idx : _GEN_630 ? _slots_12_io_out_uop_ldq_idx : _slots_11_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_632 ? _slots_14_io_out_uop_stq_idx : _GEN_631 ? _slots_13_io_out_uop_stq_idx : _GEN_630 ? _slots_12_io_out_uop_stq_idx : _slots_11_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_632 ? _slots_14_io_out_uop_pdst : _GEN_631 ? _slots_13_io_out_uop_pdst : _GEN_630 ? _slots_12_io_out_uop_pdst : _slots_11_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_632 ? _slots_14_io_out_uop_prs1 : _GEN_631 ? _slots_13_io_out_uop_prs1 : _GEN_630 ? _slots_12_io_out_uop_prs1 : _slots_11_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_632 ? _slots_14_io_out_uop_prs2 : _GEN_631 ? _slots_13_io_out_uop_prs2 : _GEN_630 ? _slots_12_io_out_uop_prs2 : _slots_11_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_632 ? _slots_14_io_out_uop_prs3 : _GEN_631 ? _slots_13_io_out_uop_prs3 : _GEN_630 ? _slots_12_io_out_uop_prs3 : _slots_11_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_632 ? _slots_14_io_out_uop_prs1_busy : _GEN_631 ? _slots_13_io_out_uop_prs1_busy : _GEN_630 ? _slots_12_io_out_uop_prs1_busy : _slots_11_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_632 ? _slots_14_io_out_uop_prs2_busy : _GEN_631 ? _slots_13_io_out_uop_prs2_busy : _GEN_630 ? _slots_12_io_out_uop_prs2_busy : _slots_11_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_632 ? _slots_14_io_out_uop_prs3_busy : _GEN_631 ? _slots_13_io_out_uop_prs3_busy : _GEN_630 ? _slots_12_io_out_uop_prs3_busy : _slots_11_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_632 ? _slots_14_io_out_uop_ppred_busy : _GEN_631 ? _slots_13_io_out_uop_ppred_busy : _GEN_630 ? _slots_12_io_out_uop_ppred_busy : _slots_11_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_632 ? _slots_14_io_out_uop_bypassable : _GEN_631 ? _slots_13_io_out_uop_bypassable : _GEN_630 ? _slots_12_io_out_uop_bypassable : _slots_11_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_632 ? _slots_14_io_out_uop_mem_cmd : _GEN_631 ? _slots_13_io_out_uop_mem_cmd : _GEN_630 ? _slots_12_io_out_uop_mem_cmd : _slots_11_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_632 ? _slots_14_io_out_uop_mem_size : _GEN_631 ? _slots_13_io_out_uop_mem_size : _GEN_630 ? _slots_12_io_out_uop_mem_size : _slots_11_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_632 ? _slots_14_io_out_uop_mem_signed : _GEN_631 ? _slots_13_io_out_uop_mem_signed : _GEN_630 ? _slots_12_io_out_uop_mem_signed : _slots_11_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_632 ? _slots_14_io_out_uop_is_fence : _GEN_631 ? _slots_13_io_out_uop_is_fence : _GEN_630 ? _slots_12_io_out_uop_is_fence : _slots_11_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_632 ? _slots_14_io_out_uop_is_amo : _GEN_631 ? _slots_13_io_out_uop_is_amo : _GEN_630 ? _slots_12_io_out_uop_is_amo : _slots_11_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_632 ? _slots_14_io_out_uop_uses_ldq : _GEN_631 ? _slots_13_io_out_uop_uses_ldq : _GEN_630 ? _slots_12_io_out_uop_uses_ldq : _slots_11_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_632 ? _slots_14_io_out_uop_uses_stq : _GEN_631 ? _slots_13_io_out_uop_uses_stq : _GEN_630 ? _slots_12_io_out_uop_uses_stq : _slots_11_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_632 ? _slots_14_io_out_uop_ldst_val : _GEN_631 ? _slots_13_io_out_uop_ldst_val : _GEN_630 ? _slots_12_io_out_uop_ldst_val : _slots_11_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_632 ? _slots_14_io_out_uop_dst_rtype : _GEN_631 ? _slots_13_io_out_uop_dst_rtype : _GEN_630 ? _slots_12_io_out_uop_dst_rtype : _slots_11_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_632 ? _slots_14_io_out_uop_lrs1_rtype : _GEN_631 ? _slots_13_io_out_uop_lrs1_rtype : _GEN_630 ? _slots_12_io_out_uop_lrs1_rtype : _slots_11_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_632 ? _slots_14_io_out_uop_lrs2_rtype : _GEN_631 ? _slots_13_io_out_uop_lrs2_rtype : _GEN_630 ? _slots_12_io_out_uop_lrs2_rtype : _slots_11_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_632 ? _slots_14_io_out_uop_fp_val : _GEN_631 ? _slots_13_io_out_uop_fp_val : _GEN_630 ? _slots_12_io_out_uop_fp_val : _slots_11_io_out_uop_fp_val),
    .io_valid                       (_slots_10_io_valid),
    .io_will_be_valid               (_slots_10_io_will_be_valid),
    .io_request                     (_slots_10_io_request),
    .io_out_uop_uopc                (_slots_10_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_10_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_10_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_10_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_10_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_10_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_10_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_10_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_10_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_10_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_10_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_10_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_10_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_10_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_10_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_10_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_10_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_10_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_10_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_10_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_10_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_10_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_10_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_10_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_10_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_10_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_10_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_10_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_10_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_10_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_10_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_10_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_10_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_10_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_10_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_10_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_10_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_10_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_10_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_10_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_10_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_10_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_10_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_10_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_10_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_10_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_10_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_10_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_10_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_10_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_10_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_10_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_10_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_10_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_10_io_uop_pc_lob),
    .io_uop_taken                   (_slots_10_io_uop_taken),
    .io_uop_imm_packed              (_slots_10_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_10_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_10_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_10_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_10_io_uop_pdst),
    .io_uop_prs1                    (_slots_10_io_uop_prs1),
    .io_uop_prs2                    (_slots_10_io_uop_prs2),
    .io_uop_bypassable              (_slots_10_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_10_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_10_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_10_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_10_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_10_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_10_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_10_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_10_io_uop_fp_val)
  );
  IssueSlot_32 slots_11 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_11_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_41),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_11_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_635 ? _slots_15_io_out_uop_uopc : _GEN_634 ? _slots_14_io_out_uop_uopc : _GEN_633 ? _slots_13_io_out_uop_uopc : _slots_12_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_635 ? _slots_15_io_out_uop_is_rvc : _GEN_634 ? _slots_14_io_out_uop_is_rvc : _GEN_633 ? _slots_13_io_out_uop_is_rvc : _slots_12_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_635 ? _slots_15_io_out_uop_fu_code : _GEN_634 ? _slots_14_io_out_uop_fu_code : _GEN_633 ? _slots_13_io_out_uop_fu_code : _slots_12_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_635 ? _slots_15_io_out_uop_iw_state : _GEN_634 ? _slots_14_io_out_uop_iw_state : _GEN_633 ? _slots_13_io_out_uop_iw_state : _slots_12_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_635 ? _slots_15_io_out_uop_iw_p1_poisoned : _GEN_634 ? _slots_14_io_out_uop_iw_p1_poisoned : _GEN_633 ? _slots_13_io_out_uop_iw_p1_poisoned : _slots_12_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_635 ? _slots_15_io_out_uop_iw_p2_poisoned : _GEN_634 ? _slots_14_io_out_uop_iw_p2_poisoned : _GEN_633 ? _slots_13_io_out_uop_iw_p2_poisoned : _slots_12_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_635 ? _slots_15_io_out_uop_is_br : _GEN_634 ? _slots_14_io_out_uop_is_br : _GEN_633 ? _slots_13_io_out_uop_is_br : _slots_12_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_635 ? _slots_15_io_out_uop_is_jalr : _GEN_634 ? _slots_14_io_out_uop_is_jalr : _GEN_633 ? _slots_13_io_out_uop_is_jalr : _slots_12_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_635 ? _slots_15_io_out_uop_is_jal : _GEN_634 ? _slots_14_io_out_uop_is_jal : _GEN_633 ? _slots_13_io_out_uop_is_jal : _slots_12_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_635 ? _slots_15_io_out_uop_is_sfb : _GEN_634 ? _slots_14_io_out_uop_is_sfb : _GEN_633 ? _slots_13_io_out_uop_is_sfb : _slots_12_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_635 ? _slots_15_io_out_uop_br_mask : _GEN_634 ? _slots_14_io_out_uop_br_mask : _GEN_633 ? _slots_13_io_out_uop_br_mask : _slots_12_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_635 ? _slots_15_io_out_uop_br_tag : _GEN_634 ? _slots_14_io_out_uop_br_tag : _GEN_633 ? _slots_13_io_out_uop_br_tag : _slots_12_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_635 ? _slots_15_io_out_uop_ftq_idx : _GEN_634 ? _slots_14_io_out_uop_ftq_idx : _GEN_633 ? _slots_13_io_out_uop_ftq_idx : _slots_12_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_635 ? _slots_15_io_out_uop_edge_inst : _GEN_634 ? _slots_14_io_out_uop_edge_inst : _GEN_633 ? _slots_13_io_out_uop_edge_inst : _slots_12_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_635 ? _slots_15_io_out_uop_pc_lob : _GEN_634 ? _slots_14_io_out_uop_pc_lob : _GEN_633 ? _slots_13_io_out_uop_pc_lob : _slots_12_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_635 ? _slots_15_io_out_uop_taken : _GEN_634 ? _slots_14_io_out_uop_taken : _GEN_633 ? _slots_13_io_out_uop_taken : _slots_12_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_635 ? _slots_15_io_out_uop_imm_packed : _GEN_634 ? _slots_14_io_out_uop_imm_packed : _GEN_633 ? _slots_13_io_out_uop_imm_packed : _slots_12_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_635 ? _slots_15_io_out_uop_rob_idx : _GEN_634 ? _slots_14_io_out_uop_rob_idx : _GEN_633 ? _slots_13_io_out_uop_rob_idx : _slots_12_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_635 ? _slots_15_io_out_uop_ldq_idx : _GEN_634 ? _slots_14_io_out_uop_ldq_idx : _GEN_633 ? _slots_13_io_out_uop_ldq_idx : _slots_12_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_635 ? _slots_15_io_out_uop_stq_idx : _GEN_634 ? _slots_14_io_out_uop_stq_idx : _GEN_633 ? _slots_13_io_out_uop_stq_idx : _slots_12_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_635 ? _slots_15_io_out_uop_pdst : _GEN_634 ? _slots_14_io_out_uop_pdst : _GEN_633 ? _slots_13_io_out_uop_pdst : _slots_12_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_635 ? _slots_15_io_out_uop_prs1 : _GEN_634 ? _slots_14_io_out_uop_prs1 : _GEN_633 ? _slots_13_io_out_uop_prs1 : _slots_12_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_635 ? _slots_15_io_out_uop_prs2 : _GEN_634 ? _slots_14_io_out_uop_prs2 : _GEN_633 ? _slots_13_io_out_uop_prs2 : _slots_12_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_635 ? _slots_15_io_out_uop_prs3 : _GEN_634 ? _slots_14_io_out_uop_prs3 : _GEN_633 ? _slots_13_io_out_uop_prs3 : _slots_12_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_635 ? _slots_15_io_out_uop_prs1_busy : _GEN_634 ? _slots_14_io_out_uop_prs1_busy : _GEN_633 ? _slots_13_io_out_uop_prs1_busy : _slots_12_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_635 ? _slots_15_io_out_uop_prs2_busy : _GEN_634 ? _slots_14_io_out_uop_prs2_busy : _GEN_633 ? _slots_13_io_out_uop_prs2_busy : _slots_12_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_635 ? _slots_15_io_out_uop_prs3_busy : _GEN_634 ? _slots_14_io_out_uop_prs3_busy : _GEN_633 ? _slots_13_io_out_uop_prs3_busy : _slots_12_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_635 ? _slots_15_io_out_uop_ppred_busy : _GEN_634 ? _slots_14_io_out_uop_ppred_busy : _GEN_633 ? _slots_13_io_out_uop_ppred_busy : _slots_12_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_635 ? _slots_15_io_out_uop_bypassable : _GEN_634 ? _slots_14_io_out_uop_bypassable : _GEN_633 ? _slots_13_io_out_uop_bypassable : _slots_12_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_635 ? _slots_15_io_out_uop_mem_cmd : _GEN_634 ? _slots_14_io_out_uop_mem_cmd : _GEN_633 ? _slots_13_io_out_uop_mem_cmd : _slots_12_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_635 ? _slots_15_io_out_uop_mem_size : _GEN_634 ? _slots_14_io_out_uop_mem_size : _GEN_633 ? _slots_13_io_out_uop_mem_size : _slots_12_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_635 ? _slots_15_io_out_uop_mem_signed : _GEN_634 ? _slots_14_io_out_uop_mem_signed : _GEN_633 ? _slots_13_io_out_uop_mem_signed : _slots_12_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_635 ? _slots_15_io_out_uop_is_fence : _GEN_634 ? _slots_14_io_out_uop_is_fence : _GEN_633 ? _slots_13_io_out_uop_is_fence : _slots_12_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_635 ? _slots_15_io_out_uop_is_amo : _GEN_634 ? _slots_14_io_out_uop_is_amo : _GEN_633 ? _slots_13_io_out_uop_is_amo : _slots_12_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_635 ? _slots_15_io_out_uop_uses_ldq : _GEN_634 ? _slots_14_io_out_uop_uses_ldq : _GEN_633 ? _slots_13_io_out_uop_uses_ldq : _slots_12_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_635 ? _slots_15_io_out_uop_uses_stq : _GEN_634 ? _slots_14_io_out_uop_uses_stq : _GEN_633 ? _slots_13_io_out_uop_uses_stq : _slots_12_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_635 ? _slots_15_io_out_uop_ldst_val : _GEN_634 ? _slots_14_io_out_uop_ldst_val : _GEN_633 ? _slots_13_io_out_uop_ldst_val : _slots_12_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_635 ? _slots_15_io_out_uop_dst_rtype : _GEN_634 ? _slots_14_io_out_uop_dst_rtype : _GEN_633 ? _slots_13_io_out_uop_dst_rtype : _slots_12_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_635 ? _slots_15_io_out_uop_lrs1_rtype : _GEN_634 ? _slots_14_io_out_uop_lrs1_rtype : _GEN_633 ? _slots_13_io_out_uop_lrs1_rtype : _slots_12_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_635 ? _slots_15_io_out_uop_lrs2_rtype : _GEN_634 ? _slots_14_io_out_uop_lrs2_rtype : _GEN_633 ? _slots_13_io_out_uop_lrs2_rtype : _slots_12_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_635 ? _slots_15_io_out_uop_fp_val : _GEN_634 ? _slots_14_io_out_uop_fp_val : _GEN_633 ? _slots_13_io_out_uop_fp_val : _slots_12_io_out_uop_fp_val),
    .io_valid                       (_slots_11_io_valid),
    .io_will_be_valid               (_slots_11_io_will_be_valid),
    .io_request                     (_slots_11_io_request),
    .io_out_uop_uopc                (_slots_11_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_11_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_11_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_11_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_11_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_11_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_11_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_11_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_11_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_11_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_11_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_11_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_11_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_11_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_11_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_11_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_11_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_11_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_11_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_11_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_11_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_11_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_11_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_11_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_11_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_11_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_11_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_11_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_11_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_11_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_11_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_11_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_11_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_11_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_11_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_11_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_11_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_11_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_11_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_11_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_11_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_11_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_11_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_11_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_11_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_11_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_11_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_11_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_11_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_11_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_11_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_11_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_11_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_11_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_11_io_uop_pc_lob),
    .io_uop_taken                   (_slots_11_io_uop_taken),
    .io_uop_imm_packed              (_slots_11_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_11_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_11_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_11_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_11_io_uop_pdst),
    .io_uop_prs1                    (_slots_11_io_uop_prs1),
    .io_uop_prs2                    (_slots_11_io_uop_prs2),
    .io_uop_bypassable              (_slots_11_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_11_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_11_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_11_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_11_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_11_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_11_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_11_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_11_io_uop_fp_val)
  );
  IssueSlot_32 slots_12 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_12_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_43),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_12_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_638 ? _slots_16_io_out_uop_uopc : _GEN_637 ? _slots_15_io_out_uop_uopc : _GEN_636 ? _slots_14_io_out_uop_uopc : _slots_13_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_638 ? _slots_16_io_out_uop_is_rvc : _GEN_637 ? _slots_15_io_out_uop_is_rvc : _GEN_636 ? _slots_14_io_out_uop_is_rvc : _slots_13_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_638 ? _slots_16_io_out_uop_fu_code : _GEN_637 ? _slots_15_io_out_uop_fu_code : _GEN_636 ? _slots_14_io_out_uop_fu_code : _slots_13_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_638 ? _slots_16_io_out_uop_iw_state : _GEN_637 ? _slots_15_io_out_uop_iw_state : _GEN_636 ? _slots_14_io_out_uop_iw_state : _slots_13_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_638 ? _slots_16_io_out_uop_iw_p1_poisoned : _GEN_637 ? _slots_15_io_out_uop_iw_p1_poisoned : _GEN_636 ? _slots_14_io_out_uop_iw_p1_poisoned : _slots_13_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_638 ? _slots_16_io_out_uop_iw_p2_poisoned : _GEN_637 ? _slots_15_io_out_uop_iw_p2_poisoned : _GEN_636 ? _slots_14_io_out_uop_iw_p2_poisoned : _slots_13_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_638 ? _slots_16_io_out_uop_is_br : _GEN_637 ? _slots_15_io_out_uop_is_br : _GEN_636 ? _slots_14_io_out_uop_is_br : _slots_13_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_638 ? _slots_16_io_out_uop_is_jalr : _GEN_637 ? _slots_15_io_out_uop_is_jalr : _GEN_636 ? _slots_14_io_out_uop_is_jalr : _slots_13_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_638 ? _slots_16_io_out_uop_is_jal : _GEN_637 ? _slots_15_io_out_uop_is_jal : _GEN_636 ? _slots_14_io_out_uop_is_jal : _slots_13_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_638 ? _slots_16_io_out_uop_is_sfb : _GEN_637 ? _slots_15_io_out_uop_is_sfb : _GEN_636 ? _slots_14_io_out_uop_is_sfb : _slots_13_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_638 ? _slots_16_io_out_uop_br_mask : _GEN_637 ? _slots_15_io_out_uop_br_mask : _GEN_636 ? _slots_14_io_out_uop_br_mask : _slots_13_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_638 ? _slots_16_io_out_uop_br_tag : _GEN_637 ? _slots_15_io_out_uop_br_tag : _GEN_636 ? _slots_14_io_out_uop_br_tag : _slots_13_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_638 ? _slots_16_io_out_uop_ftq_idx : _GEN_637 ? _slots_15_io_out_uop_ftq_idx : _GEN_636 ? _slots_14_io_out_uop_ftq_idx : _slots_13_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_638 ? _slots_16_io_out_uop_edge_inst : _GEN_637 ? _slots_15_io_out_uop_edge_inst : _GEN_636 ? _slots_14_io_out_uop_edge_inst : _slots_13_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_638 ? _slots_16_io_out_uop_pc_lob : _GEN_637 ? _slots_15_io_out_uop_pc_lob : _GEN_636 ? _slots_14_io_out_uop_pc_lob : _slots_13_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_638 ? _slots_16_io_out_uop_taken : _GEN_637 ? _slots_15_io_out_uop_taken : _GEN_636 ? _slots_14_io_out_uop_taken : _slots_13_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_638 ? _slots_16_io_out_uop_imm_packed : _GEN_637 ? _slots_15_io_out_uop_imm_packed : _GEN_636 ? _slots_14_io_out_uop_imm_packed : _slots_13_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_638 ? _slots_16_io_out_uop_rob_idx : _GEN_637 ? _slots_15_io_out_uop_rob_idx : _GEN_636 ? _slots_14_io_out_uop_rob_idx : _slots_13_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_638 ? _slots_16_io_out_uop_ldq_idx : _GEN_637 ? _slots_15_io_out_uop_ldq_idx : _GEN_636 ? _slots_14_io_out_uop_ldq_idx : _slots_13_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_638 ? _slots_16_io_out_uop_stq_idx : _GEN_637 ? _slots_15_io_out_uop_stq_idx : _GEN_636 ? _slots_14_io_out_uop_stq_idx : _slots_13_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_638 ? _slots_16_io_out_uop_pdst : _GEN_637 ? _slots_15_io_out_uop_pdst : _GEN_636 ? _slots_14_io_out_uop_pdst : _slots_13_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_638 ? _slots_16_io_out_uop_prs1 : _GEN_637 ? _slots_15_io_out_uop_prs1 : _GEN_636 ? _slots_14_io_out_uop_prs1 : _slots_13_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_638 ? _slots_16_io_out_uop_prs2 : _GEN_637 ? _slots_15_io_out_uop_prs2 : _GEN_636 ? _slots_14_io_out_uop_prs2 : _slots_13_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_638 ? _slots_16_io_out_uop_prs3 : _GEN_637 ? _slots_15_io_out_uop_prs3 : _GEN_636 ? _slots_14_io_out_uop_prs3 : _slots_13_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_638 ? _slots_16_io_out_uop_prs1_busy : _GEN_637 ? _slots_15_io_out_uop_prs1_busy : _GEN_636 ? _slots_14_io_out_uop_prs1_busy : _slots_13_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_638 ? _slots_16_io_out_uop_prs2_busy : _GEN_637 ? _slots_15_io_out_uop_prs2_busy : _GEN_636 ? _slots_14_io_out_uop_prs2_busy : _slots_13_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_638 ? _slots_16_io_out_uop_prs3_busy : _GEN_637 ? _slots_15_io_out_uop_prs3_busy : _GEN_636 ? _slots_14_io_out_uop_prs3_busy : _slots_13_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_638 ? _slots_16_io_out_uop_ppred_busy : _GEN_637 ? _slots_15_io_out_uop_ppred_busy : _GEN_636 ? _slots_14_io_out_uop_ppred_busy : _slots_13_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_638 ? _slots_16_io_out_uop_bypassable : _GEN_637 ? _slots_15_io_out_uop_bypassable : _GEN_636 ? _slots_14_io_out_uop_bypassable : _slots_13_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_638 ? _slots_16_io_out_uop_mem_cmd : _GEN_637 ? _slots_15_io_out_uop_mem_cmd : _GEN_636 ? _slots_14_io_out_uop_mem_cmd : _slots_13_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_638 ? _slots_16_io_out_uop_mem_size : _GEN_637 ? _slots_15_io_out_uop_mem_size : _GEN_636 ? _slots_14_io_out_uop_mem_size : _slots_13_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_638 ? _slots_16_io_out_uop_mem_signed : _GEN_637 ? _slots_15_io_out_uop_mem_signed : _GEN_636 ? _slots_14_io_out_uop_mem_signed : _slots_13_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_638 ? _slots_16_io_out_uop_is_fence : _GEN_637 ? _slots_15_io_out_uop_is_fence : _GEN_636 ? _slots_14_io_out_uop_is_fence : _slots_13_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_638 ? _slots_16_io_out_uop_is_amo : _GEN_637 ? _slots_15_io_out_uop_is_amo : _GEN_636 ? _slots_14_io_out_uop_is_amo : _slots_13_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_638 ? _slots_16_io_out_uop_uses_ldq : _GEN_637 ? _slots_15_io_out_uop_uses_ldq : _GEN_636 ? _slots_14_io_out_uop_uses_ldq : _slots_13_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_638 ? _slots_16_io_out_uop_uses_stq : _GEN_637 ? _slots_15_io_out_uop_uses_stq : _GEN_636 ? _slots_14_io_out_uop_uses_stq : _slots_13_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_638 ? _slots_16_io_out_uop_ldst_val : _GEN_637 ? _slots_15_io_out_uop_ldst_val : _GEN_636 ? _slots_14_io_out_uop_ldst_val : _slots_13_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_638 ? _slots_16_io_out_uop_dst_rtype : _GEN_637 ? _slots_15_io_out_uop_dst_rtype : _GEN_636 ? _slots_14_io_out_uop_dst_rtype : _slots_13_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_638 ? _slots_16_io_out_uop_lrs1_rtype : _GEN_637 ? _slots_15_io_out_uop_lrs1_rtype : _GEN_636 ? _slots_14_io_out_uop_lrs1_rtype : _slots_13_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_638 ? _slots_16_io_out_uop_lrs2_rtype : _GEN_637 ? _slots_15_io_out_uop_lrs2_rtype : _GEN_636 ? _slots_14_io_out_uop_lrs2_rtype : _slots_13_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_638 ? _slots_16_io_out_uop_fp_val : _GEN_637 ? _slots_15_io_out_uop_fp_val : _GEN_636 ? _slots_14_io_out_uop_fp_val : _slots_13_io_out_uop_fp_val),
    .io_valid                       (_slots_12_io_valid),
    .io_will_be_valid               (_slots_12_io_will_be_valid),
    .io_request                     (_slots_12_io_request),
    .io_out_uop_uopc                (_slots_12_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_12_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_12_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_12_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_12_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_12_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_12_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_12_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_12_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_12_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_12_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_12_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_12_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_12_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_12_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_12_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_12_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_12_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_12_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_12_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_12_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_12_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_12_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_12_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_12_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_12_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_12_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_12_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_12_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_12_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_12_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_12_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_12_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_12_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_12_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_12_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_12_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_12_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_12_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_12_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_12_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_12_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_12_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_12_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_12_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_12_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_12_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_12_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_12_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_12_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_12_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_12_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_12_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_12_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_12_io_uop_pc_lob),
    .io_uop_taken                   (_slots_12_io_uop_taken),
    .io_uop_imm_packed              (_slots_12_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_12_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_12_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_12_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_12_io_uop_pdst),
    .io_uop_prs1                    (_slots_12_io_uop_prs1),
    .io_uop_prs2                    (_slots_12_io_uop_prs2),
    .io_uop_bypassable              (_slots_12_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_12_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_12_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_12_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_12_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_12_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_12_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_12_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_12_io_uop_fp_val)
  );
  IssueSlot_32 slots_13 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_13_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_45),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_13_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_641 ? _slots_17_io_out_uop_uopc : _GEN_640 ? _slots_16_io_out_uop_uopc : _GEN_639 ? _slots_15_io_out_uop_uopc : _slots_14_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_641 ? _slots_17_io_out_uop_is_rvc : _GEN_640 ? _slots_16_io_out_uop_is_rvc : _GEN_639 ? _slots_15_io_out_uop_is_rvc : _slots_14_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_641 ? _slots_17_io_out_uop_fu_code : _GEN_640 ? _slots_16_io_out_uop_fu_code : _GEN_639 ? _slots_15_io_out_uop_fu_code : _slots_14_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_641 ? _slots_17_io_out_uop_iw_state : _GEN_640 ? _slots_16_io_out_uop_iw_state : _GEN_639 ? _slots_15_io_out_uop_iw_state : _slots_14_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_641 ? _slots_17_io_out_uop_iw_p1_poisoned : _GEN_640 ? _slots_16_io_out_uop_iw_p1_poisoned : _GEN_639 ? _slots_15_io_out_uop_iw_p1_poisoned : _slots_14_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_641 ? _slots_17_io_out_uop_iw_p2_poisoned : _GEN_640 ? _slots_16_io_out_uop_iw_p2_poisoned : _GEN_639 ? _slots_15_io_out_uop_iw_p2_poisoned : _slots_14_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_641 ? _slots_17_io_out_uop_is_br : _GEN_640 ? _slots_16_io_out_uop_is_br : _GEN_639 ? _slots_15_io_out_uop_is_br : _slots_14_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_641 ? _slots_17_io_out_uop_is_jalr : _GEN_640 ? _slots_16_io_out_uop_is_jalr : _GEN_639 ? _slots_15_io_out_uop_is_jalr : _slots_14_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_641 ? _slots_17_io_out_uop_is_jal : _GEN_640 ? _slots_16_io_out_uop_is_jal : _GEN_639 ? _slots_15_io_out_uop_is_jal : _slots_14_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_641 ? _slots_17_io_out_uop_is_sfb : _GEN_640 ? _slots_16_io_out_uop_is_sfb : _GEN_639 ? _slots_15_io_out_uop_is_sfb : _slots_14_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_641 ? _slots_17_io_out_uop_br_mask : _GEN_640 ? _slots_16_io_out_uop_br_mask : _GEN_639 ? _slots_15_io_out_uop_br_mask : _slots_14_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_641 ? _slots_17_io_out_uop_br_tag : _GEN_640 ? _slots_16_io_out_uop_br_tag : _GEN_639 ? _slots_15_io_out_uop_br_tag : _slots_14_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_641 ? _slots_17_io_out_uop_ftq_idx : _GEN_640 ? _slots_16_io_out_uop_ftq_idx : _GEN_639 ? _slots_15_io_out_uop_ftq_idx : _slots_14_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_641 ? _slots_17_io_out_uop_edge_inst : _GEN_640 ? _slots_16_io_out_uop_edge_inst : _GEN_639 ? _slots_15_io_out_uop_edge_inst : _slots_14_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_641 ? _slots_17_io_out_uop_pc_lob : _GEN_640 ? _slots_16_io_out_uop_pc_lob : _GEN_639 ? _slots_15_io_out_uop_pc_lob : _slots_14_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_641 ? _slots_17_io_out_uop_taken : _GEN_640 ? _slots_16_io_out_uop_taken : _GEN_639 ? _slots_15_io_out_uop_taken : _slots_14_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_641 ? _slots_17_io_out_uop_imm_packed : _GEN_640 ? _slots_16_io_out_uop_imm_packed : _GEN_639 ? _slots_15_io_out_uop_imm_packed : _slots_14_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_641 ? _slots_17_io_out_uop_rob_idx : _GEN_640 ? _slots_16_io_out_uop_rob_idx : _GEN_639 ? _slots_15_io_out_uop_rob_idx : _slots_14_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_641 ? _slots_17_io_out_uop_ldq_idx : _GEN_640 ? _slots_16_io_out_uop_ldq_idx : _GEN_639 ? _slots_15_io_out_uop_ldq_idx : _slots_14_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_641 ? _slots_17_io_out_uop_stq_idx : _GEN_640 ? _slots_16_io_out_uop_stq_idx : _GEN_639 ? _slots_15_io_out_uop_stq_idx : _slots_14_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_641 ? _slots_17_io_out_uop_pdst : _GEN_640 ? _slots_16_io_out_uop_pdst : _GEN_639 ? _slots_15_io_out_uop_pdst : _slots_14_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_641 ? _slots_17_io_out_uop_prs1 : _GEN_640 ? _slots_16_io_out_uop_prs1 : _GEN_639 ? _slots_15_io_out_uop_prs1 : _slots_14_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_641 ? _slots_17_io_out_uop_prs2 : _GEN_640 ? _slots_16_io_out_uop_prs2 : _GEN_639 ? _slots_15_io_out_uop_prs2 : _slots_14_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_641 ? _slots_17_io_out_uop_prs3 : _GEN_640 ? _slots_16_io_out_uop_prs3 : _GEN_639 ? _slots_15_io_out_uop_prs3 : _slots_14_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_641 ? _slots_17_io_out_uop_prs1_busy : _GEN_640 ? _slots_16_io_out_uop_prs1_busy : _GEN_639 ? _slots_15_io_out_uop_prs1_busy : _slots_14_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_641 ? _slots_17_io_out_uop_prs2_busy : _GEN_640 ? _slots_16_io_out_uop_prs2_busy : _GEN_639 ? _slots_15_io_out_uop_prs2_busy : _slots_14_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_641 ? _slots_17_io_out_uop_prs3_busy : _GEN_640 ? _slots_16_io_out_uop_prs3_busy : _GEN_639 ? _slots_15_io_out_uop_prs3_busy : _slots_14_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_641 ? _slots_17_io_out_uop_ppred_busy : _GEN_640 ? _slots_16_io_out_uop_ppred_busy : _GEN_639 ? _slots_15_io_out_uop_ppred_busy : _slots_14_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_641 ? _slots_17_io_out_uop_bypassable : _GEN_640 ? _slots_16_io_out_uop_bypassable : _GEN_639 ? _slots_15_io_out_uop_bypassable : _slots_14_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_641 ? _slots_17_io_out_uop_mem_cmd : _GEN_640 ? _slots_16_io_out_uop_mem_cmd : _GEN_639 ? _slots_15_io_out_uop_mem_cmd : _slots_14_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_641 ? _slots_17_io_out_uop_mem_size : _GEN_640 ? _slots_16_io_out_uop_mem_size : _GEN_639 ? _slots_15_io_out_uop_mem_size : _slots_14_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_641 ? _slots_17_io_out_uop_mem_signed : _GEN_640 ? _slots_16_io_out_uop_mem_signed : _GEN_639 ? _slots_15_io_out_uop_mem_signed : _slots_14_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_641 ? _slots_17_io_out_uop_is_fence : _GEN_640 ? _slots_16_io_out_uop_is_fence : _GEN_639 ? _slots_15_io_out_uop_is_fence : _slots_14_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_641 ? _slots_17_io_out_uop_is_amo : _GEN_640 ? _slots_16_io_out_uop_is_amo : _GEN_639 ? _slots_15_io_out_uop_is_amo : _slots_14_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_641 ? _slots_17_io_out_uop_uses_ldq : _GEN_640 ? _slots_16_io_out_uop_uses_ldq : _GEN_639 ? _slots_15_io_out_uop_uses_ldq : _slots_14_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_641 ? _slots_17_io_out_uop_uses_stq : _GEN_640 ? _slots_16_io_out_uop_uses_stq : _GEN_639 ? _slots_15_io_out_uop_uses_stq : _slots_14_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_641 ? _slots_17_io_out_uop_ldst_val : _GEN_640 ? _slots_16_io_out_uop_ldst_val : _GEN_639 ? _slots_15_io_out_uop_ldst_val : _slots_14_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_641 ? _slots_17_io_out_uop_dst_rtype : _GEN_640 ? _slots_16_io_out_uop_dst_rtype : _GEN_639 ? _slots_15_io_out_uop_dst_rtype : _slots_14_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_641 ? _slots_17_io_out_uop_lrs1_rtype : _GEN_640 ? _slots_16_io_out_uop_lrs1_rtype : _GEN_639 ? _slots_15_io_out_uop_lrs1_rtype : _slots_14_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_641 ? _slots_17_io_out_uop_lrs2_rtype : _GEN_640 ? _slots_16_io_out_uop_lrs2_rtype : _GEN_639 ? _slots_15_io_out_uop_lrs2_rtype : _slots_14_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_641 ? _slots_17_io_out_uop_fp_val : _GEN_640 ? _slots_16_io_out_uop_fp_val : _GEN_639 ? _slots_15_io_out_uop_fp_val : _slots_14_io_out_uop_fp_val),
    .io_valid                       (_slots_13_io_valid),
    .io_will_be_valid               (_slots_13_io_will_be_valid),
    .io_request                     (_slots_13_io_request),
    .io_out_uop_uopc                (_slots_13_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_13_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_13_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_13_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_13_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_13_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_13_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_13_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_13_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_13_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_13_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_13_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_13_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_13_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_13_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_13_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_13_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_13_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_13_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_13_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_13_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_13_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_13_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_13_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_13_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_13_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_13_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_13_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_13_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_13_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_13_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_13_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_13_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_13_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_13_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_13_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_13_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_13_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_13_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_13_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_13_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_13_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_13_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_13_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_13_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_13_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_13_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_13_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_13_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_13_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_13_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_13_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_13_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_13_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_13_io_uop_pc_lob),
    .io_uop_taken                   (_slots_13_io_uop_taken),
    .io_uop_imm_packed              (_slots_13_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_13_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_13_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_13_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_13_io_uop_pdst),
    .io_uop_prs1                    (_slots_13_io_uop_prs1),
    .io_uop_prs2                    (_slots_13_io_uop_prs2),
    .io_uop_bypassable              (_slots_13_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_13_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_13_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_13_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_13_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_13_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_13_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_13_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_13_io_uop_fp_val)
  );
  IssueSlot_32 slots_14 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_14_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_47),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_14_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_644 ? _slots_18_io_out_uop_uopc : _GEN_643 ? _slots_17_io_out_uop_uopc : _GEN_642 ? _slots_16_io_out_uop_uopc : _slots_15_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_644 ? _slots_18_io_out_uop_is_rvc : _GEN_643 ? _slots_17_io_out_uop_is_rvc : _GEN_642 ? _slots_16_io_out_uop_is_rvc : _slots_15_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_644 ? _slots_18_io_out_uop_fu_code : _GEN_643 ? _slots_17_io_out_uop_fu_code : _GEN_642 ? _slots_16_io_out_uop_fu_code : _slots_15_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_644 ? _slots_18_io_out_uop_iw_state : _GEN_643 ? _slots_17_io_out_uop_iw_state : _GEN_642 ? _slots_16_io_out_uop_iw_state : _slots_15_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_644 ? _slots_18_io_out_uop_iw_p1_poisoned : _GEN_643 ? _slots_17_io_out_uop_iw_p1_poisoned : _GEN_642 ? _slots_16_io_out_uop_iw_p1_poisoned : _slots_15_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_644 ? _slots_18_io_out_uop_iw_p2_poisoned : _GEN_643 ? _slots_17_io_out_uop_iw_p2_poisoned : _GEN_642 ? _slots_16_io_out_uop_iw_p2_poisoned : _slots_15_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_644 ? _slots_18_io_out_uop_is_br : _GEN_643 ? _slots_17_io_out_uop_is_br : _GEN_642 ? _slots_16_io_out_uop_is_br : _slots_15_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_644 ? _slots_18_io_out_uop_is_jalr : _GEN_643 ? _slots_17_io_out_uop_is_jalr : _GEN_642 ? _slots_16_io_out_uop_is_jalr : _slots_15_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_644 ? _slots_18_io_out_uop_is_jal : _GEN_643 ? _slots_17_io_out_uop_is_jal : _GEN_642 ? _slots_16_io_out_uop_is_jal : _slots_15_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_644 ? _slots_18_io_out_uop_is_sfb : _GEN_643 ? _slots_17_io_out_uop_is_sfb : _GEN_642 ? _slots_16_io_out_uop_is_sfb : _slots_15_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_644 ? _slots_18_io_out_uop_br_mask : _GEN_643 ? _slots_17_io_out_uop_br_mask : _GEN_642 ? _slots_16_io_out_uop_br_mask : _slots_15_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_644 ? _slots_18_io_out_uop_br_tag : _GEN_643 ? _slots_17_io_out_uop_br_tag : _GEN_642 ? _slots_16_io_out_uop_br_tag : _slots_15_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_644 ? _slots_18_io_out_uop_ftq_idx : _GEN_643 ? _slots_17_io_out_uop_ftq_idx : _GEN_642 ? _slots_16_io_out_uop_ftq_idx : _slots_15_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_644 ? _slots_18_io_out_uop_edge_inst : _GEN_643 ? _slots_17_io_out_uop_edge_inst : _GEN_642 ? _slots_16_io_out_uop_edge_inst : _slots_15_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_644 ? _slots_18_io_out_uop_pc_lob : _GEN_643 ? _slots_17_io_out_uop_pc_lob : _GEN_642 ? _slots_16_io_out_uop_pc_lob : _slots_15_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_644 ? _slots_18_io_out_uop_taken : _GEN_643 ? _slots_17_io_out_uop_taken : _GEN_642 ? _slots_16_io_out_uop_taken : _slots_15_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_644 ? _slots_18_io_out_uop_imm_packed : _GEN_643 ? _slots_17_io_out_uop_imm_packed : _GEN_642 ? _slots_16_io_out_uop_imm_packed : _slots_15_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_644 ? _slots_18_io_out_uop_rob_idx : _GEN_643 ? _slots_17_io_out_uop_rob_idx : _GEN_642 ? _slots_16_io_out_uop_rob_idx : _slots_15_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_644 ? _slots_18_io_out_uop_ldq_idx : _GEN_643 ? _slots_17_io_out_uop_ldq_idx : _GEN_642 ? _slots_16_io_out_uop_ldq_idx : _slots_15_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_644 ? _slots_18_io_out_uop_stq_idx : _GEN_643 ? _slots_17_io_out_uop_stq_idx : _GEN_642 ? _slots_16_io_out_uop_stq_idx : _slots_15_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_644 ? _slots_18_io_out_uop_pdst : _GEN_643 ? _slots_17_io_out_uop_pdst : _GEN_642 ? _slots_16_io_out_uop_pdst : _slots_15_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_644 ? _slots_18_io_out_uop_prs1 : _GEN_643 ? _slots_17_io_out_uop_prs1 : _GEN_642 ? _slots_16_io_out_uop_prs1 : _slots_15_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_644 ? _slots_18_io_out_uop_prs2 : _GEN_643 ? _slots_17_io_out_uop_prs2 : _GEN_642 ? _slots_16_io_out_uop_prs2 : _slots_15_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_644 ? _slots_18_io_out_uop_prs3 : _GEN_643 ? _slots_17_io_out_uop_prs3 : _GEN_642 ? _slots_16_io_out_uop_prs3 : _slots_15_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_644 ? _slots_18_io_out_uop_prs1_busy : _GEN_643 ? _slots_17_io_out_uop_prs1_busy : _GEN_642 ? _slots_16_io_out_uop_prs1_busy : _slots_15_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_644 ? _slots_18_io_out_uop_prs2_busy : _GEN_643 ? _slots_17_io_out_uop_prs2_busy : _GEN_642 ? _slots_16_io_out_uop_prs2_busy : _slots_15_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_644 ? _slots_18_io_out_uop_prs3_busy : _GEN_643 ? _slots_17_io_out_uop_prs3_busy : _GEN_642 ? _slots_16_io_out_uop_prs3_busy : _slots_15_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_644 ? _slots_18_io_out_uop_ppred_busy : _GEN_643 ? _slots_17_io_out_uop_ppred_busy : _GEN_642 ? _slots_16_io_out_uop_ppred_busy : _slots_15_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_644 ? _slots_18_io_out_uop_bypassable : _GEN_643 ? _slots_17_io_out_uop_bypassable : _GEN_642 ? _slots_16_io_out_uop_bypassable : _slots_15_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_644 ? _slots_18_io_out_uop_mem_cmd : _GEN_643 ? _slots_17_io_out_uop_mem_cmd : _GEN_642 ? _slots_16_io_out_uop_mem_cmd : _slots_15_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_644 ? _slots_18_io_out_uop_mem_size : _GEN_643 ? _slots_17_io_out_uop_mem_size : _GEN_642 ? _slots_16_io_out_uop_mem_size : _slots_15_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_644 ? _slots_18_io_out_uop_mem_signed : _GEN_643 ? _slots_17_io_out_uop_mem_signed : _GEN_642 ? _slots_16_io_out_uop_mem_signed : _slots_15_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_644 ? _slots_18_io_out_uop_is_fence : _GEN_643 ? _slots_17_io_out_uop_is_fence : _GEN_642 ? _slots_16_io_out_uop_is_fence : _slots_15_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_644 ? _slots_18_io_out_uop_is_amo : _GEN_643 ? _slots_17_io_out_uop_is_amo : _GEN_642 ? _slots_16_io_out_uop_is_amo : _slots_15_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_644 ? _slots_18_io_out_uop_uses_ldq : _GEN_643 ? _slots_17_io_out_uop_uses_ldq : _GEN_642 ? _slots_16_io_out_uop_uses_ldq : _slots_15_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_644 ? _slots_18_io_out_uop_uses_stq : _GEN_643 ? _slots_17_io_out_uop_uses_stq : _GEN_642 ? _slots_16_io_out_uop_uses_stq : _slots_15_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_644 ? _slots_18_io_out_uop_ldst_val : _GEN_643 ? _slots_17_io_out_uop_ldst_val : _GEN_642 ? _slots_16_io_out_uop_ldst_val : _slots_15_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_644 ? _slots_18_io_out_uop_dst_rtype : _GEN_643 ? _slots_17_io_out_uop_dst_rtype : _GEN_642 ? _slots_16_io_out_uop_dst_rtype : _slots_15_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_644 ? _slots_18_io_out_uop_lrs1_rtype : _GEN_643 ? _slots_17_io_out_uop_lrs1_rtype : _GEN_642 ? _slots_16_io_out_uop_lrs1_rtype : _slots_15_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_644 ? _slots_18_io_out_uop_lrs2_rtype : _GEN_643 ? _slots_17_io_out_uop_lrs2_rtype : _GEN_642 ? _slots_16_io_out_uop_lrs2_rtype : _slots_15_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_644 ? _slots_18_io_out_uop_fp_val : _GEN_643 ? _slots_17_io_out_uop_fp_val : _GEN_642 ? _slots_16_io_out_uop_fp_val : _slots_15_io_out_uop_fp_val),
    .io_valid                       (_slots_14_io_valid),
    .io_will_be_valid               (_slots_14_io_will_be_valid),
    .io_request                     (_slots_14_io_request),
    .io_out_uop_uopc                (_slots_14_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_14_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_14_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_14_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_14_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_14_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_14_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_14_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_14_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_14_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_14_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_14_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_14_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_14_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_14_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_14_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_14_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_14_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_14_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_14_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_14_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_14_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_14_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_14_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_14_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_14_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_14_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_14_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_14_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_14_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_14_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_14_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_14_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_14_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_14_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_14_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_14_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_14_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_14_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_14_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_14_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_14_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_14_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_14_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_14_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_14_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_14_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_14_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_14_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_14_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_14_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_14_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_14_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_14_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_14_io_uop_pc_lob),
    .io_uop_taken                   (_slots_14_io_uop_taken),
    .io_uop_imm_packed              (_slots_14_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_14_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_14_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_14_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_14_io_uop_pdst),
    .io_uop_prs1                    (_slots_14_io_uop_prs1),
    .io_uop_prs2                    (_slots_14_io_uop_prs2),
    .io_uop_bypassable              (_slots_14_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_14_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_14_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_14_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_14_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_14_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_14_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_14_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_14_io_uop_fp_val)
  );
  IssueSlot_32 slots_15 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_15_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_49),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_15_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_647 ? _slots_19_io_out_uop_uopc : _GEN_646 ? _slots_18_io_out_uop_uopc : _GEN_645 ? _slots_17_io_out_uop_uopc : _slots_16_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_647 ? _slots_19_io_out_uop_is_rvc : _GEN_646 ? _slots_18_io_out_uop_is_rvc : _GEN_645 ? _slots_17_io_out_uop_is_rvc : _slots_16_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_647 ? _slots_19_io_out_uop_fu_code : _GEN_646 ? _slots_18_io_out_uop_fu_code : _GEN_645 ? _slots_17_io_out_uop_fu_code : _slots_16_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_647 ? _slots_19_io_out_uop_iw_state : _GEN_646 ? _slots_18_io_out_uop_iw_state : _GEN_645 ? _slots_17_io_out_uop_iw_state : _slots_16_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_647 ? _slots_19_io_out_uop_iw_p1_poisoned : _GEN_646 ? _slots_18_io_out_uop_iw_p1_poisoned : _GEN_645 ? _slots_17_io_out_uop_iw_p1_poisoned : _slots_16_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_647 ? _slots_19_io_out_uop_iw_p2_poisoned : _GEN_646 ? _slots_18_io_out_uop_iw_p2_poisoned : _GEN_645 ? _slots_17_io_out_uop_iw_p2_poisoned : _slots_16_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_647 ? _slots_19_io_out_uop_is_br : _GEN_646 ? _slots_18_io_out_uop_is_br : _GEN_645 ? _slots_17_io_out_uop_is_br : _slots_16_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_647 ? _slots_19_io_out_uop_is_jalr : _GEN_646 ? _slots_18_io_out_uop_is_jalr : _GEN_645 ? _slots_17_io_out_uop_is_jalr : _slots_16_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_647 ? _slots_19_io_out_uop_is_jal : _GEN_646 ? _slots_18_io_out_uop_is_jal : _GEN_645 ? _slots_17_io_out_uop_is_jal : _slots_16_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_647 ? _slots_19_io_out_uop_is_sfb : _GEN_646 ? _slots_18_io_out_uop_is_sfb : _GEN_645 ? _slots_17_io_out_uop_is_sfb : _slots_16_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_647 ? _slots_19_io_out_uop_br_mask : _GEN_646 ? _slots_18_io_out_uop_br_mask : _GEN_645 ? _slots_17_io_out_uop_br_mask : _slots_16_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_647 ? _slots_19_io_out_uop_br_tag : _GEN_646 ? _slots_18_io_out_uop_br_tag : _GEN_645 ? _slots_17_io_out_uop_br_tag : _slots_16_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_647 ? _slots_19_io_out_uop_ftq_idx : _GEN_646 ? _slots_18_io_out_uop_ftq_idx : _GEN_645 ? _slots_17_io_out_uop_ftq_idx : _slots_16_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_647 ? _slots_19_io_out_uop_edge_inst : _GEN_646 ? _slots_18_io_out_uop_edge_inst : _GEN_645 ? _slots_17_io_out_uop_edge_inst : _slots_16_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_647 ? _slots_19_io_out_uop_pc_lob : _GEN_646 ? _slots_18_io_out_uop_pc_lob : _GEN_645 ? _slots_17_io_out_uop_pc_lob : _slots_16_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_647 ? _slots_19_io_out_uop_taken : _GEN_646 ? _slots_18_io_out_uop_taken : _GEN_645 ? _slots_17_io_out_uop_taken : _slots_16_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_647 ? _slots_19_io_out_uop_imm_packed : _GEN_646 ? _slots_18_io_out_uop_imm_packed : _GEN_645 ? _slots_17_io_out_uop_imm_packed : _slots_16_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_647 ? _slots_19_io_out_uop_rob_idx : _GEN_646 ? _slots_18_io_out_uop_rob_idx : _GEN_645 ? _slots_17_io_out_uop_rob_idx : _slots_16_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_647 ? _slots_19_io_out_uop_ldq_idx : _GEN_646 ? _slots_18_io_out_uop_ldq_idx : _GEN_645 ? _slots_17_io_out_uop_ldq_idx : _slots_16_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_647 ? _slots_19_io_out_uop_stq_idx : _GEN_646 ? _slots_18_io_out_uop_stq_idx : _GEN_645 ? _slots_17_io_out_uop_stq_idx : _slots_16_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_647 ? _slots_19_io_out_uop_pdst : _GEN_646 ? _slots_18_io_out_uop_pdst : _GEN_645 ? _slots_17_io_out_uop_pdst : _slots_16_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_647 ? _slots_19_io_out_uop_prs1 : _GEN_646 ? _slots_18_io_out_uop_prs1 : _GEN_645 ? _slots_17_io_out_uop_prs1 : _slots_16_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_647 ? _slots_19_io_out_uop_prs2 : _GEN_646 ? _slots_18_io_out_uop_prs2 : _GEN_645 ? _slots_17_io_out_uop_prs2 : _slots_16_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_647 ? _slots_19_io_out_uop_prs3 : _GEN_646 ? _slots_18_io_out_uop_prs3 : _GEN_645 ? _slots_17_io_out_uop_prs3 : _slots_16_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_647 ? _slots_19_io_out_uop_prs1_busy : _GEN_646 ? _slots_18_io_out_uop_prs1_busy : _GEN_645 ? _slots_17_io_out_uop_prs1_busy : _slots_16_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_647 ? _slots_19_io_out_uop_prs2_busy : _GEN_646 ? _slots_18_io_out_uop_prs2_busy : _GEN_645 ? _slots_17_io_out_uop_prs2_busy : _slots_16_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_647 ? _slots_19_io_out_uop_prs3_busy : _GEN_646 ? _slots_18_io_out_uop_prs3_busy : _GEN_645 ? _slots_17_io_out_uop_prs3_busy : _slots_16_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_647 ? _slots_19_io_out_uop_ppred_busy : _GEN_646 ? _slots_18_io_out_uop_ppred_busy : _GEN_645 ? _slots_17_io_out_uop_ppred_busy : _slots_16_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_647 ? _slots_19_io_out_uop_bypassable : _GEN_646 ? _slots_18_io_out_uop_bypassable : _GEN_645 ? _slots_17_io_out_uop_bypassable : _slots_16_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_647 ? _slots_19_io_out_uop_mem_cmd : _GEN_646 ? _slots_18_io_out_uop_mem_cmd : _GEN_645 ? _slots_17_io_out_uop_mem_cmd : _slots_16_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_647 ? _slots_19_io_out_uop_mem_size : _GEN_646 ? _slots_18_io_out_uop_mem_size : _GEN_645 ? _slots_17_io_out_uop_mem_size : _slots_16_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_647 ? _slots_19_io_out_uop_mem_signed : _GEN_646 ? _slots_18_io_out_uop_mem_signed : _GEN_645 ? _slots_17_io_out_uop_mem_signed : _slots_16_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_647 ? _slots_19_io_out_uop_is_fence : _GEN_646 ? _slots_18_io_out_uop_is_fence : _GEN_645 ? _slots_17_io_out_uop_is_fence : _slots_16_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_647 ? _slots_19_io_out_uop_is_amo : _GEN_646 ? _slots_18_io_out_uop_is_amo : _GEN_645 ? _slots_17_io_out_uop_is_amo : _slots_16_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_647 ? _slots_19_io_out_uop_uses_ldq : _GEN_646 ? _slots_18_io_out_uop_uses_ldq : _GEN_645 ? _slots_17_io_out_uop_uses_ldq : _slots_16_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_647 ? _slots_19_io_out_uop_uses_stq : _GEN_646 ? _slots_18_io_out_uop_uses_stq : _GEN_645 ? _slots_17_io_out_uop_uses_stq : _slots_16_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_647 ? _slots_19_io_out_uop_ldst_val : _GEN_646 ? _slots_18_io_out_uop_ldst_val : _GEN_645 ? _slots_17_io_out_uop_ldst_val : _slots_16_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_647 ? _slots_19_io_out_uop_dst_rtype : _GEN_646 ? _slots_18_io_out_uop_dst_rtype : _GEN_645 ? _slots_17_io_out_uop_dst_rtype : _slots_16_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_647 ? _slots_19_io_out_uop_lrs1_rtype : _GEN_646 ? _slots_18_io_out_uop_lrs1_rtype : _GEN_645 ? _slots_17_io_out_uop_lrs1_rtype : _slots_16_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_647 ? _slots_19_io_out_uop_lrs2_rtype : _GEN_646 ? _slots_18_io_out_uop_lrs2_rtype : _GEN_645 ? _slots_17_io_out_uop_lrs2_rtype : _slots_16_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_647 ? _slots_19_io_out_uop_fp_val : _GEN_646 ? _slots_18_io_out_uop_fp_val : _GEN_645 ? _slots_17_io_out_uop_fp_val : _slots_16_io_out_uop_fp_val),
    .io_valid                       (_slots_15_io_valid),
    .io_will_be_valid               (_slots_15_io_will_be_valid),
    .io_request                     (_slots_15_io_request),
    .io_out_uop_uopc                (_slots_15_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_15_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_15_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_15_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_15_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_15_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_15_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_15_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_15_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_15_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_15_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_15_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_15_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_15_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_15_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_15_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_15_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_15_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_15_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_15_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_15_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_15_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_15_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_15_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_15_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_15_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_15_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_15_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_15_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_15_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_15_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_15_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_15_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_15_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_15_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_15_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_15_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_15_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_15_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_15_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_15_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_15_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_15_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_15_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_15_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_15_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_15_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_15_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_15_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_15_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_15_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_15_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_15_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_15_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_15_io_uop_pc_lob),
    .io_uop_taken                   (_slots_15_io_uop_taken),
    .io_uop_imm_packed              (_slots_15_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_15_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_15_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_15_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_15_io_uop_pdst),
    .io_uop_prs1                    (_slots_15_io_uop_prs1),
    .io_uop_prs2                    (_slots_15_io_uop_prs2),
    .io_uop_bypassable              (_slots_15_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_15_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_15_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_15_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_15_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_15_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_15_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_15_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_15_io_uop_fp_val)
  );
  IssueSlot_32 slots_16 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_16_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_51),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_16_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_650 ? _slots_20_io_out_uop_uopc : _GEN_649 ? _slots_19_io_out_uop_uopc : _GEN_648 ? _slots_18_io_out_uop_uopc : _slots_17_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_650 ? _slots_20_io_out_uop_is_rvc : _GEN_649 ? _slots_19_io_out_uop_is_rvc : _GEN_648 ? _slots_18_io_out_uop_is_rvc : _slots_17_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_650 ? _slots_20_io_out_uop_fu_code : _GEN_649 ? _slots_19_io_out_uop_fu_code : _GEN_648 ? _slots_18_io_out_uop_fu_code : _slots_17_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_650 ? _slots_20_io_out_uop_iw_state : _GEN_649 ? _slots_19_io_out_uop_iw_state : _GEN_648 ? _slots_18_io_out_uop_iw_state : _slots_17_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_650 ? _slots_20_io_out_uop_iw_p1_poisoned : _GEN_649 ? _slots_19_io_out_uop_iw_p1_poisoned : _GEN_648 ? _slots_18_io_out_uop_iw_p1_poisoned : _slots_17_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_650 ? _slots_20_io_out_uop_iw_p2_poisoned : _GEN_649 ? _slots_19_io_out_uop_iw_p2_poisoned : _GEN_648 ? _slots_18_io_out_uop_iw_p2_poisoned : _slots_17_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_650 ? _slots_20_io_out_uop_is_br : _GEN_649 ? _slots_19_io_out_uop_is_br : _GEN_648 ? _slots_18_io_out_uop_is_br : _slots_17_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_650 ? _slots_20_io_out_uop_is_jalr : _GEN_649 ? _slots_19_io_out_uop_is_jalr : _GEN_648 ? _slots_18_io_out_uop_is_jalr : _slots_17_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_650 ? _slots_20_io_out_uop_is_jal : _GEN_649 ? _slots_19_io_out_uop_is_jal : _GEN_648 ? _slots_18_io_out_uop_is_jal : _slots_17_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_650 ? _slots_20_io_out_uop_is_sfb : _GEN_649 ? _slots_19_io_out_uop_is_sfb : _GEN_648 ? _slots_18_io_out_uop_is_sfb : _slots_17_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_650 ? _slots_20_io_out_uop_br_mask : _GEN_649 ? _slots_19_io_out_uop_br_mask : _GEN_648 ? _slots_18_io_out_uop_br_mask : _slots_17_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_650 ? _slots_20_io_out_uop_br_tag : _GEN_649 ? _slots_19_io_out_uop_br_tag : _GEN_648 ? _slots_18_io_out_uop_br_tag : _slots_17_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_650 ? _slots_20_io_out_uop_ftq_idx : _GEN_649 ? _slots_19_io_out_uop_ftq_idx : _GEN_648 ? _slots_18_io_out_uop_ftq_idx : _slots_17_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_650 ? _slots_20_io_out_uop_edge_inst : _GEN_649 ? _slots_19_io_out_uop_edge_inst : _GEN_648 ? _slots_18_io_out_uop_edge_inst : _slots_17_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_650 ? _slots_20_io_out_uop_pc_lob : _GEN_649 ? _slots_19_io_out_uop_pc_lob : _GEN_648 ? _slots_18_io_out_uop_pc_lob : _slots_17_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_650 ? _slots_20_io_out_uop_taken : _GEN_649 ? _slots_19_io_out_uop_taken : _GEN_648 ? _slots_18_io_out_uop_taken : _slots_17_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_650 ? _slots_20_io_out_uop_imm_packed : _GEN_649 ? _slots_19_io_out_uop_imm_packed : _GEN_648 ? _slots_18_io_out_uop_imm_packed : _slots_17_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_650 ? _slots_20_io_out_uop_rob_idx : _GEN_649 ? _slots_19_io_out_uop_rob_idx : _GEN_648 ? _slots_18_io_out_uop_rob_idx : _slots_17_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_650 ? _slots_20_io_out_uop_ldq_idx : _GEN_649 ? _slots_19_io_out_uop_ldq_idx : _GEN_648 ? _slots_18_io_out_uop_ldq_idx : _slots_17_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_650 ? _slots_20_io_out_uop_stq_idx : _GEN_649 ? _slots_19_io_out_uop_stq_idx : _GEN_648 ? _slots_18_io_out_uop_stq_idx : _slots_17_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_650 ? _slots_20_io_out_uop_pdst : _GEN_649 ? _slots_19_io_out_uop_pdst : _GEN_648 ? _slots_18_io_out_uop_pdst : _slots_17_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_650 ? _slots_20_io_out_uop_prs1 : _GEN_649 ? _slots_19_io_out_uop_prs1 : _GEN_648 ? _slots_18_io_out_uop_prs1 : _slots_17_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_650 ? _slots_20_io_out_uop_prs2 : _GEN_649 ? _slots_19_io_out_uop_prs2 : _GEN_648 ? _slots_18_io_out_uop_prs2 : _slots_17_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_650 ? _slots_20_io_out_uop_prs3 : _GEN_649 ? _slots_19_io_out_uop_prs3 : _GEN_648 ? _slots_18_io_out_uop_prs3 : _slots_17_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_650 ? _slots_20_io_out_uop_prs1_busy : _GEN_649 ? _slots_19_io_out_uop_prs1_busy : _GEN_648 ? _slots_18_io_out_uop_prs1_busy : _slots_17_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_650 ? _slots_20_io_out_uop_prs2_busy : _GEN_649 ? _slots_19_io_out_uop_prs2_busy : _GEN_648 ? _slots_18_io_out_uop_prs2_busy : _slots_17_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_650 ? _slots_20_io_out_uop_prs3_busy : _GEN_649 ? _slots_19_io_out_uop_prs3_busy : _GEN_648 ? _slots_18_io_out_uop_prs3_busy : _slots_17_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_650 ? _slots_20_io_out_uop_ppred_busy : _GEN_649 ? _slots_19_io_out_uop_ppred_busy : _GEN_648 ? _slots_18_io_out_uop_ppred_busy : _slots_17_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_650 ? _slots_20_io_out_uop_bypassable : _GEN_649 ? _slots_19_io_out_uop_bypassable : _GEN_648 ? _slots_18_io_out_uop_bypassable : _slots_17_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_650 ? _slots_20_io_out_uop_mem_cmd : _GEN_649 ? _slots_19_io_out_uop_mem_cmd : _GEN_648 ? _slots_18_io_out_uop_mem_cmd : _slots_17_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_650 ? _slots_20_io_out_uop_mem_size : _GEN_649 ? _slots_19_io_out_uop_mem_size : _GEN_648 ? _slots_18_io_out_uop_mem_size : _slots_17_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_650 ? _slots_20_io_out_uop_mem_signed : _GEN_649 ? _slots_19_io_out_uop_mem_signed : _GEN_648 ? _slots_18_io_out_uop_mem_signed : _slots_17_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_650 ? _slots_20_io_out_uop_is_fence : _GEN_649 ? _slots_19_io_out_uop_is_fence : _GEN_648 ? _slots_18_io_out_uop_is_fence : _slots_17_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_650 ? _slots_20_io_out_uop_is_amo : _GEN_649 ? _slots_19_io_out_uop_is_amo : _GEN_648 ? _slots_18_io_out_uop_is_amo : _slots_17_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_650 ? _slots_20_io_out_uop_uses_ldq : _GEN_649 ? _slots_19_io_out_uop_uses_ldq : _GEN_648 ? _slots_18_io_out_uop_uses_ldq : _slots_17_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_650 ? _slots_20_io_out_uop_uses_stq : _GEN_649 ? _slots_19_io_out_uop_uses_stq : _GEN_648 ? _slots_18_io_out_uop_uses_stq : _slots_17_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_650 ? _slots_20_io_out_uop_ldst_val : _GEN_649 ? _slots_19_io_out_uop_ldst_val : _GEN_648 ? _slots_18_io_out_uop_ldst_val : _slots_17_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_650 ? _slots_20_io_out_uop_dst_rtype : _GEN_649 ? _slots_19_io_out_uop_dst_rtype : _GEN_648 ? _slots_18_io_out_uop_dst_rtype : _slots_17_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_650 ? _slots_20_io_out_uop_lrs1_rtype : _GEN_649 ? _slots_19_io_out_uop_lrs1_rtype : _GEN_648 ? _slots_18_io_out_uop_lrs1_rtype : _slots_17_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_650 ? _slots_20_io_out_uop_lrs2_rtype : _GEN_649 ? _slots_19_io_out_uop_lrs2_rtype : _GEN_648 ? _slots_18_io_out_uop_lrs2_rtype : _slots_17_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_650 ? _slots_20_io_out_uop_fp_val : _GEN_649 ? _slots_19_io_out_uop_fp_val : _GEN_648 ? _slots_18_io_out_uop_fp_val : _slots_17_io_out_uop_fp_val),
    .io_valid                       (_slots_16_io_valid),
    .io_will_be_valid               (_slots_16_io_will_be_valid),
    .io_request                     (_slots_16_io_request),
    .io_out_uop_uopc                (_slots_16_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_16_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_16_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_16_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_16_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_16_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_16_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_16_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_16_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_16_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_16_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_16_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_16_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_16_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_16_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_16_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_16_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_16_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_16_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_16_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_16_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_16_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_16_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_16_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_16_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_16_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_16_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_16_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_16_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_16_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_16_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_16_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_16_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_16_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_16_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_16_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_16_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_16_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_16_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_16_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_16_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_16_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_16_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_16_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_16_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_16_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_16_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_16_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_16_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_16_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_16_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_16_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_16_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_16_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_16_io_uop_pc_lob),
    .io_uop_taken                   (_slots_16_io_uop_taken),
    .io_uop_imm_packed              (_slots_16_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_16_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_16_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_16_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_16_io_uop_pdst),
    .io_uop_prs1                    (_slots_16_io_uop_prs1),
    .io_uop_prs2                    (_slots_16_io_uop_prs2),
    .io_uop_bypassable              (_slots_16_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_16_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_16_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_16_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_16_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_16_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_16_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_16_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_16_io_uop_fp_val)
  );
  IssueSlot_32 slots_17 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_17_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_53),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_17_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_653 ? _slots_21_io_out_uop_uopc : _GEN_652 ? _slots_20_io_out_uop_uopc : _GEN_651 ? _slots_19_io_out_uop_uopc : _slots_18_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_653 ? _slots_21_io_out_uop_is_rvc : _GEN_652 ? _slots_20_io_out_uop_is_rvc : _GEN_651 ? _slots_19_io_out_uop_is_rvc : _slots_18_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_653 ? _slots_21_io_out_uop_fu_code : _GEN_652 ? _slots_20_io_out_uop_fu_code : _GEN_651 ? _slots_19_io_out_uop_fu_code : _slots_18_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_653 ? _slots_21_io_out_uop_iw_state : _GEN_652 ? _slots_20_io_out_uop_iw_state : _GEN_651 ? _slots_19_io_out_uop_iw_state : _slots_18_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_653 ? _slots_21_io_out_uop_iw_p1_poisoned : _GEN_652 ? _slots_20_io_out_uop_iw_p1_poisoned : _GEN_651 ? _slots_19_io_out_uop_iw_p1_poisoned : _slots_18_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_653 ? _slots_21_io_out_uop_iw_p2_poisoned : _GEN_652 ? _slots_20_io_out_uop_iw_p2_poisoned : _GEN_651 ? _slots_19_io_out_uop_iw_p2_poisoned : _slots_18_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_653 ? _slots_21_io_out_uop_is_br : _GEN_652 ? _slots_20_io_out_uop_is_br : _GEN_651 ? _slots_19_io_out_uop_is_br : _slots_18_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_653 ? _slots_21_io_out_uop_is_jalr : _GEN_652 ? _slots_20_io_out_uop_is_jalr : _GEN_651 ? _slots_19_io_out_uop_is_jalr : _slots_18_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_653 ? _slots_21_io_out_uop_is_jal : _GEN_652 ? _slots_20_io_out_uop_is_jal : _GEN_651 ? _slots_19_io_out_uop_is_jal : _slots_18_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_653 ? _slots_21_io_out_uop_is_sfb : _GEN_652 ? _slots_20_io_out_uop_is_sfb : _GEN_651 ? _slots_19_io_out_uop_is_sfb : _slots_18_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_653 ? _slots_21_io_out_uop_br_mask : _GEN_652 ? _slots_20_io_out_uop_br_mask : _GEN_651 ? _slots_19_io_out_uop_br_mask : _slots_18_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_653 ? _slots_21_io_out_uop_br_tag : _GEN_652 ? _slots_20_io_out_uop_br_tag : _GEN_651 ? _slots_19_io_out_uop_br_tag : _slots_18_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_653 ? _slots_21_io_out_uop_ftq_idx : _GEN_652 ? _slots_20_io_out_uop_ftq_idx : _GEN_651 ? _slots_19_io_out_uop_ftq_idx : _slots_18_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_653 ? _slots_21_io_out_uop_edge_inst : _GEN_652 ? _slots_20_io_out_uop_edge_inst : _GEN_651 ? _slots_19_io_out_uop_edge_inst : _slots_18_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_653 ? _slots_21_io_out_uop_pc_lob : _GEN_652 ? _slots_20_io_out_uop_pc_lob : _GEN_651 ? _slots_19_io_out_uop_pc_lob : _slots_18_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_653 ? _slots_21_io_out_uop_taken : _GEN_652 ? _slots_20_io_out_uop_taken : _GEN_651 ? _slots_19_io_out_uop_taken : _slots_18_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_653 ? _slots_21_io_out_uop_imm_packed : _GEN_652 ? _slots_20_io_out_uop_imm_packed : _GEN_651 ? _slots_19_io_out_uop_imm_packed : _slots_18_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_653 ? _slots_21_io_out_uop_rob_idx : _GEN_652 ? _slots_20_io_out_uop_rob_idx : _GEN_651 ? _slots_19_io_out_uop_rob_idx : _slots_18_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_653 ? _slots_21_io_out_uop_ldq_idx : _GEN_652 ? _slots_20_io_out_uop_ldq_idx : _GEN_651 ? _slots_19_io_out_uop_ldq_idx : _slots_18_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_653 ? _slots_21_io_out_uop_stq_idx : _GEN_652 ? _slots_20_io_out_uop_stq_idx : _GEN_651 ? _slots_19_io_out_uop_stq_idx : _slots_18_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_653 ? _slots_21_io_out_uop_pdst : _GEN_652 ? _slots_20_io_out_uop_pdst : _GEN_651 ? _slots_19_io_out_uop_pdst : _slots_18_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_653 ? _slots_21_io_out_uop_prs1 : _GEN_652 ? _slots_20_io_out_uop_prs1 : _GEN_651 ? _slots_19_io_out_uop_prs1 : _slots_18_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_653 ? _slots_21_io_out_uop_prs2 : _GEN_652 ? _slots_20_io_out_uop_prs2 : _GEN_651 ? _slots_19_io_out_uop_prs2 : _slots_18_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_653 ? _slots_21_io_out_uop_prs3 : _GEN_652 ? _slots_20_io_out_uop_prs3 : _GEN_651 ? _slots_19_io_out_uop_prs3 : _slots_18_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_653 ? _slots_21_io_out_uop_prs1_busy : _GEN_652 ? _slots_20_io_out_uop_prs1_busy : _GEN_651 ? _slots_19_io_out_uop_prs1_busy : _slots_18_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_653 ? _slots_21_io_out_uop_prs2_busy : _GEN_652 ? _slots_20_io_out_uop_prs2_busy : _GEN_651 ? _slots_19_io_out_uop_prs2_busy : _slots_18_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_653 ? _slots_21_io_out_uop_prs3_busy : _GEN_652 ? _slots_20_io_out_uop_prs3_busy : _GEN_651 ? _slots_19_io_out_uop_prs3_busy : _slots_18_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_653 ? _slots_21_io_out_uop_ppred_busy : _GEN_652 ? _slots_20_io_out_uop_ppred_busy : _GEN_651 ? _slots_19_io_out_uop_ppred_busy : _slots_18_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_653 ? _slots_21_io_out_uop_bypassable : _GEN_652 ? _slots_20_io_out_uop_bypassable : _GEN_651 ? _slots_19_io_out_uop_bypassable : _slots_18_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_653 ? _slots_21_io_out_uop_mem_cmd : _GEN_652 ? _slots_20_io_out_uop_mem_cmd : _GEN_651 ? _slots_19_io_out_uop_mem_cmd : _slots_18_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_653 ? _slots_21_io_out_uop_mem_size : _GEN_652 ? _slots_20_io_out_uop_mem_size : _GEN_651 ? _slots_19_io_out_uop_mem_size : _slots_18_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_653 ? _slots_21_io_out_uop_mem_signed : _GEN_652 ? _slots_20_io_out_uop_mem_signed : _GEN_651 ? _slots_19_io_out_uop_mem_signed : _slots_18_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_653 ? _slots_21_io_out_uop_is_fence : _GEN_652 ? _slots_20_io_out_uop_is_fence : _GEN_651 ? _slots_19_io_out_uop_is_fence : _slots_18_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_653 ? _slots_21_io_out_uop_is_amo : _GEN_652 ? _slots_20_io_out_uop_is_amo : _GEN_651 ? _slots_19_io_out_uop_is_amo : _slots_18_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_653 ? _slots_21_io_out_uop_uses_ldq : _GEN_652 ? _slots_20_io_out_uop_uses_ldq : _GEN_651 ? _slots_19_io_out_uop_uses_ldq : _slots_18_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_653 ? _slots_21_io_out_uop_uses_stq : _GEN_652 ? _slots_20_io_out_uop_uses_stq : _GEN_651 ? _slots_19_io_out_uop_uses_stq : _slots_18_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_653 ? _slots_21_io_out_uop_ldst_val : _GEN_652 ? _slots_20_io_out_uop_ldst_val : _GEN_651 ? _slots_19_io_out_uop_ldst_val : _slots_18_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_653 ? _slots_21_io_out_uop_dst_rtype : _GEN_652 ? _slots_20_io_out_uop_dst_rtype : _GEN_651 ? _slots_19_io_out_uop_dst_rtype : _slots_18_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_653 ? _slots_21_io_out_uop_lrs1_rtype : _GEN_652 ? _slots_20_io_out_uop_lrs1_rtype : _GEN_651 ? _slots_19_io_out_uop_lrs1_rtype : _slots_18_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_653 ? _slots_21_io_out_uop_lrs2_rtype : _GEN_652 ? _slots_20_io_out_uop_lrs2_rtype : _GEN_651 ? _slots_19_io_out_uop_lrs2_rtype : _slots_18_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_653 ? _slots_21_io_out_uop_fp_val : _GEN_652 ? _slots_20_io_out_uop_fp_val : _GEN_651 ? _slots_19_io_out_uop_fp_val : _slots_18_io_out_uop_fp_val),
    .io_valid                       (_slots_17_io_valid),
    .io_will_be_valid               (_slots_17_io_will_be_valid),
    .io_request                     (_slots_17_io_request),
    .io_out_uop_uopc                (_slots_17_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_17_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_17_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_17_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_17_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_17_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_17_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_17_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_17_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_17_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_17_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_17_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_17_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_17_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_17_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_17_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_17_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_17_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_17_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_17_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_17_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_17_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_17_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_17_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_17_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_17_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_17_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_17_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_17_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_17_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_17_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_17_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_17_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_17_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_17_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_17_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_17_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_17_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_17_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_17_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_17_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_17_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_17_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_17_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_17_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_17_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_17_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_17_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_17_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_17_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_17_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_17_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_17_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_17_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_17_io_uop_pc_lob),
    .io_uop_taken                   (_slots_17_io_uop_taken),
    .io_uop_imm_packed              (_slots_17_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_17_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_17_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_17_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_17_io_uop_pdst),
    .io_uop_prs1                    (_slots_17_io_uop_prs1),
    .io_uop_prs2                    (_slots_17_io_uop_prs2),
    .io_uop_bypassable              (_slots_17_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_17_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_17_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_17_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_17_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_17_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_17_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_17_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_17_io_uop_fp_val)
  );
  IssueSlot_32 slots_18 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_18_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_55),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_18_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_656 ? _slots_22_io_out_uop_uopc : _GEN_655 ? _slots_21_io_out_uop_uopc : _GEN_654 ? _slots_20_io_out_uop_uopc : _slots_19_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_656 ? _slots_22_io_out_uop_is_rvc : _GEN_655 ? _slots_21_io_out_uop_is_rvc : _GEN_654 ? _slots_20_io_out_uop_is_rvc : _slots_19_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_656 ? _slots_22_io_out_uop_fu_code : _GEN_655 ? _slots_21_io_out_uop_fu_code : _GEN_654 ? _slots_20_io_out_uop_fu_code : _slots_19_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_656 ? _slots_22_io_out_uop_iw_state : _GEN_655 ? _slots_21_io_out_uop_iw_state : _GEN_654 ? _slots_20_io_out_uop_iw_state : _slots_19_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_656 ? _slots_22_io_out_uop_iw_p1_poisoned : _GEN_655 ? _slots_21_io_out_uop_iw_p1_poisoned : _GEN_654 ? _slots_20_io_out_uop_iw_p1_poisoned : _slots_19_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_656 ? _slots_22_io_out_uop_iw_p2_poisoned : _GEN_655 ? _slots_21_io_out_uop_iw_p2_poisoned : _GEN_654 ? _slots_20_io_out_uop_iw_p2_poisoned : _slots_19_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_656 ? _slots_22_io_out_uop_is_br : _GEN_655 ? _slots_21_io_out_uop_is_br : _GEN_654 ? _slots_20_io_out_uop_is_br : _slots_19_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_656 ? _slots_22_io_out_uop_is_jalr : _GEN_655 ? _slots_21_io_out_uop_is_jalr : _GEN_654 ? _slots_20_io_out_uop_is_jalr : _slots_19_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_656 ? _slots_22_io_out_uop_is_jal : _GEN_655 ? _slots_21_io_out_uop_is_jal : _GEN_654 ? _slots_20_io_out_uop_is_jal : _slots_19_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_656 ? _slots_22_io_out_uop_is_sfb : _GEN_655 ? _slots_21_io_out_uop_is_sfb : _GEN_654 ? _slots_20_io_out_uop_is_sfb : _slots_19_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_656 ? _slots_22_io_out_uop_br_mask : _GEN_655 ? _slots_21_io_out_uop_br_mask : _GEN_654 ? _slots_20_io_out_uop_br_mask : _slots_19_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_656 ? _slots_22_io_out_uop_br_tag : _GEN_655 ? _slots_21_io_out_uop_br_tag : _GEN_654 ? _slots_20_io_out_uop_br_tag : _slots_19_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_656 ? _slots_22_io_out_uop_ftq_idx : _GEN_655 ? _slots_21_io_out_uop_ftq_idx : _GEN_654 ? _slots_20_io_out_uop_ftq_idx : _slots_19_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_656 ? _slots_22_io_out_uop_edge_inst : _GEN_655 ? _slots_21_io_out_uop_edge_inst : _GEN_654 ? _slots_20_io_out_uop_edge_inst : _slots_19_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_656 ? _slots_22_io_out_uop_pc_lob : _GEN_655 ? _slots_21_io_out_uop_pc_lob : _GEN_654 ? _slots_20_io_out_uop_pc_lob : _slots_19_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_656 ? _slots_22_io_out_uop_taken : _GEN_655 ? _slots_21_io_out_uop_taken : _GEN_654 ? _slots_20_io_out_uop_taken : _slots_19_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_656 ? _slots_22_io_out_uop_imm_packed : _GEN_655 ? _slots_21_io_out_uop_imm_packed : _GEN_654 ? _slots_20_io_out_uop_imm_packed : _slots_19_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_656 ? _slots_22_io_out_uop_rob_idx : _GEN_655 ? _slots_21_io_out_uop_rob_idx : _GEN_654 ? _slots_20_io_out_uop_rob_idx : _slots_19_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_656 ? _slots_22_io_out_uop_ldq_idx : _GEN_655 ? _slots_21_io_out_uop_ldq_idx : _GEN_654 ? _slots_20_io_out_uop_ldq_idx : _slots_19_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_656 ? _slots_22_io_out_uop_stq_idx : _GEN_655 ? _slots_21_io_out_uop_stq_idx : _GEN_654 ? _slots_20_io_out_uop_stq_idx : _slots_19_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_656 ? _slots_22_io_out_uop_pdst : _GEN_655 ? _slots_21_io_out_uop_pdst : _GEN_654 ? _slots_20_io_out_uop_pdst : _slots_19_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_656 ? _slots_22_io_out_uop_prs1 : _GEN_655 ? _slots_21_io_out_uop_prs1 : _GEN_654 ? _slots_20_io_out_uop_prs1 : _slots_19_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_656 ? _slots_22_io_out_uop_prs2 : _GEN_655 ? _slots_21_io_out_uop_prs2 : _GEN_654 ? _slots_20_io_out_uop_prs2 : _slots_19_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_656 ? _slots_22_io_out_uop_prs3 : _GEN_655 ? _slots_21_io_out_uop_prs3 : _GEN_654 ? _slots_20_io_out_uop_prs3 : _slots_19_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_656 ? _slots_22_io_out_uop_prs1_busy : _GEN_655 ? _slots_21_io_out_uop_prs1_busy : _GEN_654 ? _slots_20_io_out_uop_prs1_busy : _slots_19_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_656 ? _slots_22_io_out_uop_prs2_busy : _GEN_655 ? _slots_21_io_out_uop_prs2_busy : _GEN_654 ? _slots_20_io_out_uop_prs2_busy : _slots_19_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_656 ? _slots_22_io_out_uop_prs3_busy : _GEN_655 ? _slots_21_io_out_uop_prs3_busy : _GEN_654 ? _slots_20_io_out_uop_prs3_busy : _slots_19_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_656 ? _slots_22_io_out_uop_ppred_busy : _GEN_655 ? _slots_21_io_out_uop_ppred_busy : _GEN_654 ? _slots_20_io_out_uop_ppred_busy : _slots_19_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_656 ? _slots_22_io_out_uop_bypassable : _GEN_655 ? _slots_21_io_out_uop_bypassable : _GEN_654 ? _slots_20_io_out_uop_bypassable : _slots_19_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_656 ? _slots_22_io_out_uop_mem_cmd : _GEN_655 ? _slots_21_io_out_uop_mem_cmd : _GEN_654 ? _slots_20_io_out_uop_mem_cmd : _slots_19_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_656 ? _slots_22_io_out_uop_mem_size : _GEN_655 ? _slots_21_io_out_uop_mem_size : _GEN_654 ? _slots_20_io_out_uop_mem_size : _slots_19_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_656 ? _slots_22_io_out_uop_mem_signed : _GEN_655 ? _slots_21_io_out_uop_mem_signed : _GEN_654 ? _slots_20_io_out_uop_mem_signed : _slots_19_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_656 ? _slots_22_io_out_uop_is_fence : _GEN_655 ? _slots_21_io_out_uop_is_fence : _GEN_654 ? _slots_20_io_out_uop_is_fence : _slots_19_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_656 ? _slots_22_io_out_uop_is_amo : _GEN_655 ? _slots_21_io_out_uop_is_amo : _GEN_654 ? _slots_20_io_out_uop_is_amo : _slots_19_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_656 ? _slots_22_io_out_uop_uses_ldq : _GEN_655 ? _slots_21_io_out_uop_uses_ldq : _GEN_654 ? _slots_20_io_out_uop_uses_ldq : _slots_19_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_656 ? _slots_22_io_out_uop_uses_stq : _GEN_655 ? _slots_21_io_out_uop_uses_stq : _GEN_654 ? _slots_20_io_out_uop_uses_stq : _slots_19_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_656 ? _slots_22_io_out_uop_ldst_val : _GEN_655 ? _slots_21_io_out_uop_ldst_val : _GEN_654 ? _slots_20_io_out_uop_ldst_val : _slots_19_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_656 ? _slots_22_io_out_uop_dst_rtype : _GEN_655 ? _slots_21_io_out_uop_dst_rtype : _GEN_654 ? _slots_20_io_out_uop_dst_rtype : _slots_19_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_656 ? _slots_22_io_out_uop_lrs1_rtype : _GEN_655 ? _slots_21_io_out_uop_lrs1_rtype : _GEN_654 ? _slots_20_io_out_uop_lrs1_rtype : _slots_19_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_656 ? _slots_22_io_out_uop_lrs2_rtype : _GEN_655 ? _slots_21_io_out_uop_lrs2_rtype : _GEN_654 ? _slots_20_io_out_uop_lrs2_rtype : _slots_19_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_656 ? _slots_22_io_out_uop_fp_val : _GEN_655 ? _slots_21_io_out_uop_fp_val : _GEN_654 ? _slots_20_io_out_uop_fp_val : _slots_19_io_out_uop_fp_val),
    .io_valid                       (_slots_18_io_valid),
    .io_will_be_valid               (_slots_18_io_will_be_valid),
    .io_request                     (_slots_18_io_request),
    .io_out_uop_uopc                (_slots_18_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_18_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_18_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_18_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_18_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_18_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_18_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_18_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_18_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_18_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_18_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_18_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_18_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_18_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_18_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_18_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_18_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_18_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_18_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_18_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_18_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_18_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_18_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_18_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_18_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_18_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_18_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_18_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_18_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_18_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_18_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_18_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_18_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_18_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_18_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_18_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_18_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_18_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_18_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_18_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_18_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_18_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_18_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_18_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_18_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_18_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_18_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_18_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_18_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_18_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_18_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_18_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_18_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_18_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_18_io_uop_pc_lob),
    .io_uop_taken                   (_slots_18_io_uop_taken),
    .io_uop_imm_packed              (_slots_18_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_18_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_18_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_18_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_18_io_uop_pdst),
    .io_uop_prs1                    (_slots_18_io_uop_prs1),
    .io_uop_prs2                    (_slots_18_io_uop_prs2),
    .io_uop_bypassable              (_slots_18_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_18_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_18_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_18_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_18_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_18_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_18_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_18_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_18_io_uop_fp_val)
  );
  IssueSlot_32 slots_19 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_19_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_57),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_19_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_659 ? _slots_23_io_out_uop_uopc : _GEN_658 ? _slots_22_io_out_uop_uopc : _GEN_657 ? _slots_21_io_out_uop_uopc : _slots_20_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_659 ? _slots_23_io_out_uop_is_rvc : _GEN_658 ? _slots_22_io_out_uop_is_rvc : _GEN_657 ? _slots_21_io_out_uop_is_rvc : _slots_20_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_659 ? _slots_23_io_out_uop_fu_code : _GEN_658 ? _slots_22_io_out_uop_fu_code : _GEN_657 ? _slots_21_io_out_uop_fu_code : _slots_20_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_659 ? _slots_23_io_out_uop_iw_state : _GEN_658 ? _slots_22_io_out_uop_iw_state : _GEN_657 ? _slots_21_io_out_uop_iw_state : _slots_20_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_659 ? _slots_23_io_out_uop_iw_p1_poisoned : _GEN_658 ? _slots_22_io_out_uop_iw_p1_poisoned : _GEN_657 ? _slots_21_io_out_uop_iw_p1_poisoned : _slots_20_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_659 ? _slots_23_io_out_uop_iw_p2_poisoned : _GEN_658 ? _slots_22_io_out_uop_iw_p2_poisoned : _GEN_657 ? _slots_21_io_out_uop_iw_p2_poisoned : _slots_20_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_659 ? _slots_23_io_out_uop_is_br : _GEN_658 ? _slots_22_io_out_uop_is_br : _GEN_657 ? _slots_21_io_out_uop_is_br : _slots_20_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_659 ? _slots_23_io_out_uop_is_jalr : _GEN_658 ? _slots_22_io_out_uop_is_jalr : _GEN_657 ? _slots_21_io_out_uop_is_jalr : _slots_20_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_659 ? _slots_23_io_out_uop_is_jal : _GEN_658 ? _slots_22_io_out_uop_is_jal : _GEN_657 ? _slots_21_io_out_uop_is_jal : _slots_20_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_659 ? _slots_23_io_out_uop_is_sfb : _GEN_658 ? _slots_22_io_out_uop_is_sfb : _GEN_657 ? _slots_21_io_out_uop_is_sfb : _slots_20_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_659 ? _slots_23_io_out_uop_br_mask : _GEN_658 ? _slots_22_io_out_uop_br_mask : _GEN_657 ? _slots_21_io_out_uop_br_mask : _slots_20_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_659 ? _slots_23_io_out_uop_br_tag : _GEN_658 ? _slots_22_io_out_uop_br_tag : _GEN_657 ? _slots_21_io_out_uop_br_tag : _slots_20_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_659 ? _slots_23_io_out_uop_ftq_idx : _GEN_658 ? _slots_22_io_out_uop_ftq_idx : _GEN_657 ? _slots_21_io_out_uop_ftq_idx : _slots_20_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_659 ? _slots_23_io_out_uop_edge_inst : _GEN_658 ? _slots_22_io_out_uop_edge_inst : _GEN_657 ? _slots_21_io_out_uop_edge_inst : _slots_20_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_659 ? _slots_23_io_out_uop_pc_lob : _GEN_658 ? _slots_22_io_out_uop_pc_lob : _GEN_657 ? _slots_21_io_out_uop_pc_lob : _slots_20_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_659 ? _slots_23_io_out_uop_taken : _GEN_658 ? _slots_22_io_out_uop_taken : _GEN_657 ? _slots_21_io_out_uop_taken : _slots_20_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_659 ? _slots_23_io_out_uop_imm_packed : _GEN_658 ? _slots_22_io_out_uop_imm_packed : _GEN_657 ? _slots_21_io_out_uop_imm_packed : _slots_20_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_659 ? _slots_23_io_out_uop_rob_idx : _GEN_658 ? _slots_22_io_out_uop_rob_idx : _GEN_657 ? _slots_21_io_out_uop_rob_idx : _slots_20_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_659 ? _slots_23_io_out_uop_ldq_idx : _GEN_658 ? _slots_22_io_out_uop_ldq_idx : _GEN_657 ? _slots_21_io_out_uop_ldq_idx : _slots_20_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_659 ? _slots_23_io_out_uop_stq_idx : _GEN_658 ? _slots_22_io_out_uop_stq_idx : _GEN_657 ? _slots_21_io_out_uop_stq_idx : _slots_20_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_659 ? _slots_23_io_out_uop_pdst : _GEN_658 ? _slots_22_io_out_uop_pdst : _GEN_657 ? _slots_21_io_out_uop_pdst : _slots_20_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_659 ? _slots_23_io_out_uop_prs1 : _GEN_658 ? _slots_22_io_out_uop_prs1 : _GEN_657 ? _slots_21_io_out_uop_prs1 : _slots_20_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_659 ? _slots_23_io_out_uop_prs2 : _GEN_658 ? _slots_22_io_out_uop_prs2 : _GEN_657 ? _slots_21_io_out_uop_prs2 : _slots_20_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_659 ? _slots_23_io_out_uop_prs3 : _GEN_658 ? _slots_22_io_out_uop_prs3 : _GEN_657 ? _slots_21_io_out_uop_prs3 : _slots_20_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_659 ? _slots_23_io_out_uop_prs1_busy : _GEN_658 ? _slots_22_io_out_uop_prs1_busy : _GEN_657 ? _slots_21_io_out_uop_prs1_busy : _slots_20_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_659 ? _slots_23_io_out_uop_prs2_busy : _GEN_658 ? _slots_22_io_out_uop_prs2_busy : _GEN_657 ? _slots_21_io_out_uop_prs2_busy : _slots_20_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_659 ? _slots_23_io_out_uop_prs3_busy : _GEN_658 ? _slots_22_io_out_uop_prs3_busy : _GEN_657 ? _slots_21_io_out_uop_prs3_busy : _slots_20_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_659 ? _slots_23_io_out_uop_ppred_busy : _GEN_658 ? _slots_22_io_out_uop_ppred_busy : _GEN_657 ? _slots_21_io_out_uop_ppred_busy : _slots_20_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_659 ? _slots_23_io_out_uop_bypassable : _GEN_658 ? _slots_22_io_out_uop_bypassable : _GEN_657 ? _slots_21_io_out_uop_bypassable : _slots_20_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_659 ? _slots_23_io_out_uop_mem_cmd : _GEN_658 ? _slots_22_io_out_uop_mem_cmd : _GEN_657 ? _slots_21_io_out_uop_mem_cmd : _slots_20_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_659 ? _slots_23_io_out_uop_mem_size : _GEN_658 ? _slots_22_io_out_uop_mem_size : _GEN_657 ? _slots_21_io_out_uop_mem_size : _slots_20_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_659 ? _slots_23_io_out_uop_mem_signed : _GEN_658 ? _slots_22_io_out_uop_mem_signed : _GEN_657 ? _slots_21_io_out_uop_mem_signed : _slots_20_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_659 ? _slots_23_io_out_uop_is_fence : _GEN_658 ? _slots_22_io_out_uop_is_fence : _GEN_657 ? _slots_21_io_out_uop_is_fence : _slots_20_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_659 ? _slots_23_io_out_uop_is_amo : _GEN_658 ? _slots_22_io_out_uop_is_amo : _GEN_657 ? _slots_21_io_out_uop_is_amo : _slots_20_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_659 ? _slots_23_io_out_uop_uses_ldq : _GEN_658 ? _slots_22_io_out_uop_uses_ldq : _GEN_657 ? _slots_21_io_out_uop_uses_ldq : _slots_20_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_659 ? _slots_23_io_out_uop_uses_stq : _GEN_658 ? _slots_22_io_out_uop_uses_stq : _GEN_657 ? _slots_21_io_out_uop_uses_stq : _slots_20_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_659 ? _slots_23_io_out_uop_ldst_val : _GEN_658 ? _slots_22_io_out_uop_ldst_val : _GEN_657 ? _slots_21_io_out_uop_ldst_val : _slots_20_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_659 ? _slots_23_io_out_uop_dst_rtype : _GEN_658 ? _slots_22_io_out_uop_dst_rtype : _GEN_657 ? _slots_21_io_out_uop_dst_rtype : _slots_20_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_659 ? _slots_23_io_out_uop_lrs1_rtype : _GEN_658 ? _slots_22_io_out_uop_lrs1_rtype : _GEN_657 ? _slots_21_io_out_uop_lrs1_rtype : _slots_20_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_659 ? _slots_23_io_out_uop_lrs2_rtype : _GEN_658 ? _slots_22_io_out_uop_lrs2_rtype : _GEN_657 ? _slots_21_io_out_uop_lrs2_rtype : _slots_20_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_659 ? _slots_23_io_out_uop_fp_val : _GEN_658 ? _slots_22_io_out_uop_fp_val : _GEN_657 ? _slots_21_io_out_uop_fp_val : _slots_20_io_out_uop_fp_val),
    .io_valid                       (_slots_19_io_valid),
    .io_will_be_valid               (_slots_19_io_will_be_valid),
    .io_request                     (_slots_19_io_request),
    .io_out_uop_uopc                (_slots_19_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_19_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_19_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_19_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_19_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_19_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_19_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_19_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_19_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_19_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_19_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_19_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_19_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_19_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_19_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_19_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_19_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_19_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_19_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_19_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_19_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_19_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_19_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_19_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_19_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_19_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_19_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_19_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_19_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_19_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_19_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_19_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_19_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_19_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_19_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_19_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_19_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_19_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_19_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_19_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_19_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_19_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_19_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_19_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_19_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_19_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_19_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_19_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_19_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_19_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_19_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_19_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_19_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_19_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_19_io_uop_pc_lob),
    .io_uop_taken                   (_slots_19_io_uop_taken),
    .io_uop_imm_packed              (_slots_19_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_19_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_19_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_19_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_19_io_uop_pdst),
    .io_uop_prs1                    (_slots_19_io_uop_prs1),
    .io_uop_prs2                    (_slots_19_io_uop_prs2),
    .io_uop_bypassable              (_slots_19_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_19_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_19_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_19_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_19_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_19_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_19_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_19_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_19_io_uop_fp_val)
  );
  IssueSlot_32 slots_20 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_20_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_59),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_20_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_662 ? _slots_24_io_out_uop_uopc : _GEN_661 ? _slots_23_io_out_uop_uopc : _GEN_660 ? _slots_22_io_out_uop_uopc : _slots_21_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_662 ? _slots_24_io_out_uop_is_rvc : _GEN_661 ? _slots_23_io_out_uop_is_rvc : _GEN_660 ? _slots_22_io_out_uop_is_rvc : _slots_21_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_662 ? _slots_24_io_out_uop_fu_code : _GEN_661 ? _slots_23_io_out_uop_fu_code : _GEN_660 ? _slots_22_io_out_uop_fu_code : _slots_21_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_662 ? _slots_24_io_out_uop_iw_state : _GEN_661 ? _slots_23_io_out_uop_iw_state : _GEN_660 ? _slots_22_io_out_uop_iw_state : _slots_21_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_662 ? _slots_24_io_out_uop_iw_p1_poisoned : _GEN_661 ? _slots_23_io_out_uop_iw_p1_poisoned : _GEN_660 ? _slots_22_io_out_uop_iw_p1_poisoned : _slots_21_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_662 ? _slots_24_io_out_uop_iw_p2_poisoned : _GEN_661 ? _slots_23_io_out_uop_iw_p2_poisoned : _GEN_660 ? _slots_22_io_out_uop_iw_p2_poisoned : _slots_21_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_662 ? _slots_24_io_out_uop_is_br : _GEN_661 ? _slots_23_io_out_uop_is_br : _GEN_660 ? _slots_22_io_out_uop_is_br : _slots_21_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_662 ? _slots_24_io_out_uop_is_jalr : _GEN_661 ? _slots_23_io_out_uop_is_jalr : _GEN_660 ? _slots_22_io_out_uop_is_jalr : _slots_21_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_662 ? _slots_24_io_out_uop_is_jal : _GEN_661 ? _slots_23_io_out_uop_is_jal : _GEN_660 ? _slots_22_io_out_uop_is_jal : _slots_21_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_662 ? _slots_24_io_out_uop_is_sfb : _GEN_661 ? _slots_23_io_out_uop_is_sfb : _GEN_660 ? _slots_22_io_out_uop_is_sfb : _slots_21_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_662 ? _slots_24_io_out_uop_br_mask : _GEN_661 ? _slots_23_io_out_uop_br_mask : _GEN_660 ? _slots_22_io_out_uop_br_mask : _slots_21_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_662 ? _slots_24_io_out_uop_br_tag : _GEN_661 ? _slots_23_io_out_uop_br_tag : _GEN_660 ? _slots_22_io_out_uop_br_tag : _slots_21_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_662 ? _slots_24_io_out_uop_ftq_idx : _GEN_661 ? _slots_23_io_out_uop_ftq_idx : _GEN_660 ? _slots_22_io_out_uop_ftq_idx : _slots_21_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_662 ? _slots_24_io_out_uop_edge_inst : _GEN_661 ? _slots_23_io_out_uop_edge_inst : _GEN_660 ? _slots_22_io_out_uop_edge_inst : _slots_21_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_662 ? _slots_24_io_out_uop_pc_lob : _GEN_661 ? _slots_23_io_out_uop_pc_lob : _GEN_660 ? _slots_22_io_out_uop_pc_lob : _slots_21_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_662 ? _slots_24_io_out_uop_taken : _GEN_661 ? _slots_23_io_out_uop_taken : _GEN_660 ? _slots_22_io_out_uop_taken : _slots_21_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_662 ? _slots_24_io_out_uop_imm_packed : _GEN_661 ? _slots_23_io_out_uop_imm_packed : _GEN_660 ? _slots_22_io_out_uop_imm_packed : _slots_21_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_662 ? _slots_24_io_out_uop_rob_idx : _GEN_661 ? _slots_23_io_out_uop_rob_idx : _GEN_660 ? _slots_22_io_out_uop_rob_idx : _slots_21_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_662 ? _slots_24_io_out_uop_ldq_idx : _GEN_661 ? _slots_23_io_out_uop_ldq_idx : _GEN_660 ? _slots_22_io_out_uop_ldq_idx : _slots_21_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_662 ? _slots_24_io_out_uop_stq_idx : _GEN_661 ? _slots_23_io_out_uop_stq_idx : _GEN_660 ? _slots_22_io_out_uop_stq_idx : _slots_21_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_662 ? _slots_24_io_out_uop_pdst : _GEN_661 ? _slots_23_io_out_uop_pdst : _GEN_660 ? _slots_22_io_out_uop_pdst : _slots_21_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_662 ? _slots_24_io_out_uop_prs1 : _GEN_661 ? _slots_23_io_out_uop_prs1 : _GEN_660 ? _slots_22_io_out_uop_prs1 : _slots_21_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_662 ? _slots_24_io_out_uop_prs2 : _GEN_661 ? _slots_23_io_out_uop_prs2 : _GEN_660 ? _slots_22_io_out_uop_prs2 : _slots_21_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_662 ? _slots_24_io_out_uop_prs3 : _GEN_661 ? _slots_23_io_out_uop_prs3 : _GEN_660 ? _slots_22_io_out_uop_prs3 : _slots_21_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_662 ? _slots_24_io_out_uop_prs1_busy : _GEN_661 ? _slots_23_io_out_uop_prs1_busy : _GEN_660 ? _slots_22_io_out_uop_prs1_busy : _slots_21_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_662 ? _slots_24_io_out_uop_prs2_busy : _GEN_661 ? _slots_23_io_out_uop_prs2_busy : _GEN_660 ? _slots_22_io_out_uop_prs2_busy : _slots_21_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_662 ? _slots_24_io_out_uop_prs3_busy : _GEN_661 ? _slots_23_io_out_uop_prs3_busy : _GEN_660 ? _slots_22_io_out_uop_prs3_busy : _slots_21_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_662 ? _slots_24_io_out_uop_ppred_busy : _GEN_661 ? _slots_23_io_out_uop_ppred_busy : _GEN_660 ? _slots_22_io_out_uop_ppred_busy : _slots_21_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_662 ? _slots_24_io_out_uop_bypassable : _GEN_661 ? _slots_23_io_out_uop_bypassable : _GEN_660 ? _slots_22_io_out_uop_bypassable : _slots_21_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_662 ? _slots_24_io_out_uop_mem_cmd : _GEN_661 ? _slots_23_io_out_uop_mem_cmd : _GEN_660 ? _slots_22_io_out_uop_mem_cmd : _slots_21_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_662 ? _slots_24_io_out_uop_mem_size : _GEN_661 ? _slots_23_io_out_uop_mem_size : _GEN_660 ? _slots_22_io_out_uop_mem_size : _slots_21_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_662 ? _slots_24_io_out_uop_mem_signed : _GEN_661 ? _slots_23_io_out_uop_mem_signed : _GEN_660 ? _slots_22_io_out_uop_mem_signed : _slots_21_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_662 ? _slots_24_io_out_uop_is_fence : _GEN_661 ? _slots_23_io_out_uop_is_fence : _GEN_660 ? _slots_22_io_out_uop_is_fence : _slots_21_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_662 ? _slots_24_io_out_uop_is_amo : _GEN_661 ? _slots_23_io_out_uop_is_amo : _GEN_660 ? _slots_22_io_out_uop_is_amo : _slots_21_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_662 ? _slots_24_io_out_uop_uses_ldq : _GEN_661 ? _slots_23_io_out_uop_uses_ldq : _GEN_660 ? _slots_22_io_out_uop_uses_ldq : _slots_21_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_662 ? _slots_24_io_out_uop_uses_stq : _GEN_661 ? _slots_23_io_out_uop_uses_stq : _GEN_660 ? _slots_22_io_out_uop_uses_stq : _slots_21_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_662 ? _slots_24_io_out_uop_ldst_val : _GEN_661 ? _slots_23_io_out_uop_ldst_val : _GEN_660 ? _slots_22_io_out_uop_ldst_val : _slots_21_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_662 ? _slots_24_io_out_uop_dst_rtype : _GEN_661 ? _slots_23_io_out_uop_dst_rtype : _GEN_660 ? _slots_22_io_out_uop_dst_rtype : _slots_21_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_662 ? _slots_24_io_out_uop_lrs1_rtype : _GEN_661 ? _slots_23_io_out_uop_lrs1_rtype : _GEN_660 ? _slots_22_io_out_uop_lrs1_rtype : _slots_21_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_662 ? _slots_24_io_out_uop_lrs2_rtype : _GEN_661 ? _slots_23_io_out_uop_lrs2_rtype : _GEN_660 ? _slots_22_io_out_uop_lrs2_rtype : _slots_21_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_662 ? _slots_24_io_out_uop_fp_val : _GEN_661 ? _slots_23_io_out_uop_fp_val : _GEN_660 ? _slots_22_io_out_uop_fp_val : _slots_21_io_out_uop_fp_val),
    .io_valid                       (_slots_20_io_valid),
    .io_will_be_valid               (_slots_20_io_will_be_valid),
    .io_request                     (_slots_20_io_request),
    .io_out_uop_uopc                (_slots_20_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_20_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_20_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_20_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_20_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_20_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_20_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_20_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_20_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_20_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_20_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_20_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_20_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_20_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_20_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_20_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_20_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_20_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_20_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_20_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_20_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_20_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_20_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_20_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_20_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_20_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_20_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_20_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_20_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_20_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_20_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_20_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_20_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_20_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_20_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_20_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_20_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_20_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_20_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_20_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_20_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_20_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_20_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_20_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_20_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_20_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_20_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_20_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_20_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_20_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_20_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_20_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_20_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_20_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_20_io_uop_pc_lob),
    .io_uop_taken                   (_slots_20_io_uop_taken),
    .io_uop_imm_packed              (_slots_20_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_20_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_20_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_20_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_20_io_uop_pdst),
    .io_uop_prs1                    (_slots_20_io_uop_prs1),
    .io_uop_prs2                    (_slots_20_io_uop_prs2),
    .io_uop_bypassable              (_slots_20_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_20_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_20_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_20_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_20_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_20_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_20_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_20_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_20_io_uop_fp_val)
  );
  IssueSlot_32 slots_21 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_21_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_61),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_21_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_665 ? _slots_25_io_out_uop_uopc : _GEN_664 ? _slots_24_io_out_uop_uopc : _GEN_663 ? _slots_23_io_out_uop_uopc : _slots_22_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_665 ? _slots_25_io_out_uop_is_rvc : _GEN_664 ? _slots_24_io_out_uop_is_rvc : _GEN_663 ? _slots_23_io_out_uop_is_rvc : _slots_22_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_665 ? _slots_25_io_out_uop_fu_code : _GEN_664 ? _slots_24_io_out_uop_fu_code : _GEN_663 ? _slots_23_io_out_uop_fu_code : _slots_22_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_665 ? _slots_25_io_out_uop_iw_state : _GEN_664 ? _slots_24_io_out_uop_iw_state : _GEN_663 ? _slots_23_io_out_uop_iw_state : _slots_22_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_665 ? _slots_25_io_out_uop_iw_p1_poisoned : _GEN_664 ? _slots_24_io_out_uop_iw_p1_poisoned : _GEN_663 ? _slots_23_io_out_uop_iw_p1_poisoned : _slots_22_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_665 ? _slots_25_io_out_uop_iw_p2_poisoned : _GEN_664 ? _slots_24_io_out_uop_iw_p2_poisoned : _GEN_663 ? _slots_23_io_out_uop_iw_p2_poisoned : _slots_22_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_665 ? _slots_25_io_out_uop_is_br : _GEN_664 ? _slots_24_io_out_uop_is_br : _GEN_663 ? _slots_23_io_out_uop_is_br : _slots_22_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_665 ? _slots_25_io_out_uop_is_jalr : _GEN_664 ? _slots_24_io_out_uop_is_jalr : _GEN_663 ? _slots_23_io_out_uop_is_jalr : _slots_22_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_665 ? _slots_25_io_out_uop_is_jal : _GEN_664 ? _slots_24_io_out_uop_is_jal : _GEN_663 ? _slots_23_io_out_uop_is_jal : _slots_22_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_665 ? _slots_25_io_out_uop_is_sfb : _GEN_664 ? _slots_24_io_out_uop_is_sfb : _GEN_663 ? _slots_23_io_out_uop_is_sfb : _slots_22_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_665 ? _slots_25_io_out_uop_br_mask : _GEN_664 ? _slots_24_io_out_uop_br_mask : _GEN_663 ? _slots_23_io_out_uop_br_mask : _slots_22_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_665 ? _slots_25_io_out_uop_br_tag : _GEN_664 ? _slots_24_io_out_uop_br_tag : _GEN_663 ? _slots_23_io_out_uop_br_tag : _slots_22_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_665 ? _slots_25_io_out_uop_ftq_idx : _GEN_664 ? _slots_24_io_out_uop_ftq_idx : _GEN_663 ? _slots_23_io_out_uop_ftq_idx : _slots_22_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_665 ? _slots_25_io_out_uop_edge_inst : _GEN_664 ? _slots_24_io_out_uop_edge_inst : _GEN_663 ? _slots_23_io_out_uop_edge_inst : _slots_22_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_665 ? _slots_25_io_out_uop_pc_lob : _GEN_664 ? _slots_24_io_out_uop_pc_lob : _GEN_663 ? _slots_23_io_out_uop_pc_lob : _slots_22_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_665 ? _slots_25_io_out_uop_taken : _GEN_664 ? _slots_24_io_out_uop_taken : _GEN_663 ? _slots_23_io_out_uop_taken : _slots_22_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_665 ? _slots_25_io_out_uop_imm_packed : _GEN_664 ? _slots_24_io_out_uop_imm_packed : _GEN_663 ? _slots_23_io_out_uop_imm_packed : _slots_22_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_665 ? _slots_25_io_out_uop_rob_idx : _GEN_664 ? _slots_24_io_out_uop_rob_idx : _GEN_663 ? _slots_23_io_out_uop_rob_idx : _slots_22_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_665 ? _slots_25_io_out_uop_ldq_idx : _GEN_664 ? _slots_24_io_out_uop_ldq_idx : _GEN_663 ? _slots_23_io_out_uop_ldq_idx : _slots_22_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_665 ? _slots_25_io_out_uop_stq_idx : _GEN_664 ? _slots_24_io_out_uop_stq_idx : _GEN_663 ? _slots_23_io_out_uop_stq_idx : _slots_22_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_665 ? _slots_25_io_out_uop_pdst : _GEN_664 ? _slots_24_io_out_uop_pdst : _GEN_663 ? _slots_23_io_out_uop_pdst : _slots_22_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_665 ? _slots_25_io_out_uop_prs1 : _GEN_664 ? _slots_24_io_out_uop_prs1 : _GEN_663 ? _slots_23_io_out_uop_prs1 : _slots_22_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_665 ? _slots_25_io_out_uop_prs2 : _GEN_664 ? _slots_24_io_out_uop_prs2 : _GEN_663 ? _slots_23_io_out_uop_prs2 : _slots_22_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_665 ? _slots_25_io_out_uop_prs3 : _GEN_664 ? _slots_24_io_out_uop_prs3 : _GEN_663 ? _slots_23_io_out_uop_prs3 : _slots_22_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_665 ? _slots_25_io_out_uop_prs1_busy : _GEN_664 ? _slots_24_io_out_uop_prs1_busy : _GEN_663 ? _slots_23_io_out_uop_prs1_busy : _slots_22_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_665 ? _slots_25_io_out_uop_prs2_busy : _GEN_664 ? _slots_24_io_out_uop_prs2_busy : _GEN_663 ? _slots_23_io_out_uop_prs2_busy : _slots_22_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_665 ? _slots_25_io_out_uop_prs3_busy : _GEN_664 ? _slots_24_io_out_uop_prs3_busy : _GEN_663 ? _slots_23_io_out_uop_prs3_busy : _slots_22_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_665 ? _slots_25_io_out_uop_ppred_busy : _GEN_664 ? _slots_24_io_out_uop_ppred_busy : _GEN_663 ? _slots_23_io_out_uop_ppred_busy : _slots_22_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_665 ? _slots_25_io_out_uop_bypassable : _GEN_664 ? _slots_24_io_out_uop_bypassable : _GEN_663 ? _slots_23_io_out_uop_bypassable : _slots_22_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_665 ? _slots_25_io_out_uop_mem_cmd : _GEN_664 ? _slots_24_io_out_uop_mem_cmd : _GEN_663 ? _slots_23_io_out_uop_mem_cmd : _slots_22_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_665 ? _slots_25_io_out_uop_mem_size : _GEN_664 ? _slots_24_io_out_uop_mem_size : _GEN_663 ? _slots_23_io_out_uop_mem_size : _slots_22_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_665 ? _slots_25_io_out_uop_mem_signed : _GEN_664 ? _slots_24_io_out_uop_mem_signed : _GEN_663 ? _slots_23_io_out_uop_mem_signed : _slots_22_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_665 ? _slots_25_io_out_uop_is_fence : _GEN_664 ? _slots_24_io_out_uop_is_fence : _GEN_663 ? _slots_23_io_out_uop_is_fence : _slots_22_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_665 ? _slots_25_io_out_uop_is_amo : _GEN_664 ? _slots_24_io_out_uop_is_amo : _GEN_663 ? _slots_23_io_out_uop_is_amo : _slots_22_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_665 ? _slots_25_io_out_uop_uses_ldq : _GEN_664 ? _slots_24_io_out_uop_uses_ldq : _GEN_663 ? _slots_23_io_out_uop_uses_ldq : _slots_22_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_665 ? _slots_25_io_out_uop_uses_stq : _GEN_664 ? _slots_24_io_out_uop_uses_stq : _GEN_663 ? _slots_23_io_out_uop_uses_stq : _slots_22_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_665 ? _slots_25_io_out_uop_ldst_val : _GEN_664 ? _slots_24_io_out_uop_ldst_val : _GEN_663 ? _slots_23_io_out_uop_ldst_val : _slots_22_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_665 ? _slots_25_io_out_uop_dst_rtype : _GEN_664 ? _slots_24_io_out_uop_dst_rtype : _GEN_663 ? _slots_23_io_out_uop_dst_rtype : _slots_22_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_665 ? _slots_25_io_out_uop_lrs1_rtype : _GEN_664 ? _slots_24_io_out_uop_lrs1_rtype : _GEN_663 ? _slots_23_io_out_uop_lrs1_rtype : _slots_22_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_665 ? _slots_25_io_out_uop_lrs2_rtype : _GEN_664 ? _slots_24_io_out_uop_lrs2_rtype : _GEN_663 ? _slots_23_io_out_uop_lrs2_rtype : _slots_22_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_665 ? _slots_25_io_out_uop_fp_val : _GEN_664 ? _slots_24_io_out_uop_fp_val : _GEN_663 ? _slots_23_io_out_uop_fp_val : _slots_22_io_out_uop_fp_val),
    .io_valid                       (_slots_21_io_valid),
    .io_will_be_valid               (_slots_21_io_will_be_valid),
    .io_request                     (_slots_21_io_request),
    .io_out_uop_uopc                (_slots_21_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_21_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_21_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_21_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_21_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_21_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_21_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_21_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_21_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_21_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_21_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_21_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_21_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_21_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_21_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_21_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_21_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_21_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_21_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_21_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_21_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_21_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_21_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_21_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_21_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_21_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_21_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_21_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_21_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_21_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_21_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_21_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_21_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_21_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_21_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_21_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_21_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_21_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_21_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_21_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_21_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_21_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_21_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_21_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_21_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_21_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_21_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_21_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_21_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_21_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_21_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_21_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_21_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_21_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_21_io_uop_pc_lob),
    .io_uop_taken                   (_slots_21_io_uop_taken),
    .io_uop_imm_packed              (_slots_21_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_21_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_21_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_21_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_21_io_uop_pdst),
    .io_uop_prs1                    (_slots_21_io_uop_prs1),
    .io_uop_prs2                    (_slots_21_io_uop_prs2),
    .io_uop_bypassable              (_slots_21_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_21_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_21_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_21_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_21_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_21_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_21_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_21_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_21_io_uop_fp_val)
  );
  IssueSlot_32 slots_22 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_22_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_63),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_22_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_668 ? _slots_26_io_out_uop_uopc : _GEN_667 ? _slots_25_io_out_uop_uopc : _GEN_666 ? _slots_24_io_out_uop_uopc : _slots_23_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_668 ? _slots_26_io_out_uop_is_rvc : _GEN_667 ? _slots_25_io_out_uop_is_rvc : _GEN_666 ? _slots_24_io_out_uop_is_rvc : _slots_23_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_668 ? _slots_26_io_out_uop_fu_code : _GEN_667 ? _slots_25_io_out_uop_fu_code : _GEN_666 ? _slots_24_io_out_uop_fu_code : _slots_23_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_668 ? _slots_26_io_out_uop_iw_state : _GEN_667 ? _slots_25_io_out_uop_iw_state : _GEN_666 ? _slots_24_io_out_uop_iw_state : _slots_23_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_668 ? _slots_26_io_out_uop_iw_p1_poisoned : _GEN_667 ? _slots_25_io_out_uop_iw_p1_poisoned : _GEN_666 ? _slots_24_io_out_uop_iw_p1_poisoned : _slots_23_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_668 ? _slots_26_io_out_uop_iw_p2_poisoned : _GEN_667 ? _slots_25_io_out_uop_iw_p2_poisoned : _GEN_666 ? _slots_24_io_out_uop_iw_p2_poisoned : _slots_23_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_668 ? _slots_26_io_out_uop_is_br : _GEN_667 ? _slots_25_io_out_uop_is_br : _GEN_666 ? _slots_24_io_out_uop_is_br : _slots_23_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_668 ? _slots_26_io_out_uop_is_jalr : _GEN_667 ? _slots_25_io_out_uop_is_jalr : _GEN_666 ? _slots_24_io_out_uop_is_jalr : _slots_23_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_668 ? _slots_26_io_out_uop_is_jal : _GEN_667 ? _slots_25_io_out_uop_is_jal : _GEN_666 ? _slots_24_io_out_uop_is_jal : _slots_23_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_668 ? _slots_26_io_out_uop_is_sfb : _GEN_667 ? _slots_25_io_out_uop_is_sfb : _GEN_666 ? _slots_24_io_out_uop_is_sfb : _slots_23_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_668 ? _slots_26_io_out_uop_br_mask : _GEN_667 ? _slots_25_io_out_uop_br_mask : _GEN_666 ? _slots_24_io_out_uop_br_mask : _slots_23_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_668 ? _slots_26_io_out_uop_br_tag : _GEN_667 ? _slots_25_io_out_uop_br_tag : _GEN_666 ? _slots_24_io_out_uop_br_tag : _slots_23_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_668 ? _slots_26_io_out_uop_ftq_idx : _GEN_667 ? _slots_25_io_out_uop_ftq_idx : _GEN_666 ? _slots_24_io_out_uop_ftq_idx : _slots_23_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_668 ? _slots_26_io_out_uop_edge_inst : _GEN_667 ? _slots_25_io_out_uop_edge_inst : _GEN_666 ? _slots_24_io_out_uop_edge_inst : _slots_23_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_668 ? _slots_26_io_out_uop_pc_lob : _GEN_667 ? _slots_25_io_out_uop_pc_lob : _GEN_666 ? _slots_24_io_out_uop_pc_lob : _slots_23_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_668 ? _slots_26_io_out_uop_taken : _GEN_667 ? _slots_25_io_out_uop_taken : _GEN_666 ? _slots_24_io_out_uop_taken : _slots_23_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_668 ? _slots_26_io_out_uop_imm_packed : _GEN_667 ? _slots_25_io_out_uop_imm_packed : _GEN_666 ? _slots_24_io_out_uop_imm_packed : _slots_23_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_668 ? _slots_26_io_out_uop_rob_idx : _GEN_667 ? _slots_25_io_out_uop_rob_idx : _GEN_666 ? _slots_24_io_out_uop_rob_idx : _slots_23_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_668 ? _slots_26_io_out_uop_ldq_idx : _GEN_667 ? _slots_25_io_out_uop_ldq_idx : _GEN_666 ? _slots_24_io_out_uop_ldq_idx : _slots_23_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_668 ? _slots_26_io_out_uop_stq_idx : _GEN_667 ? _slots_25_io_out_uop_stq_idx : _GEN_666 ? _slots_24_io_out_uop_stq_idx : _slots_23_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_668 ? _slots_26_io_out_uop_pdst : _GEN_667 ? _slots_25_io_out_uop_pdst : _GEN_666 ? _slots_24_io_out_uop_pdst : _slots_23_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_668 ? _slots_26_io_out_uop_prs1 : _GEN_667 ? _slots_25_io_out_uop_prs1 : _GEN_666 ? _slots_24_io_out_uop_prs1 : _slots_23_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_668 ? _slots_26_io_out_uop_prs2 : _GEN_667 ? _slots_25_io_out_uop_prs2 : _GEN_666 ? _slots_24_io_out_uop_prs2 : _slots_23_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_668 ? _slots_26_io_out_uop_prs3 : _GEN_667 ? _slots_25_io_out_uop_prs3 : _GEN_666 ? _slots_24_io_out_uop_prs3 : _slots_23_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_668 ? _slots_26_io_out_uop_prs1_busy : _GEN_667 ? _slots_25_io_out_uop_prs1_busy : _GEN_666 ? _slots_24_io_out_uop_prs1_busy : _slots_23_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_668 ? _slots_26_io_out_uop_prs2_busy : _GEN_667 ? _slots_25_io_out_uop_prs2_busy : _GEN_666 ? _slots_24_io_out_uop_prs2_busy : _slots_23_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_668 ? _slots_26_io_out_uop_prs3_busy : _GEN_667 ? _slots_25_io_out_uop_prs3_busy : _GEN_666 ? _slots_24_io_out_uop_prs3_busy : _slots_23_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_668 ? _slots_26_io_out_uop_ppred_busy : _GEN_667 ? _slots_25_io_out_uop_ppred_busy : _GEN_666 ? _slots_24_io_out_uop_ppred_busy : _slots_23_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_668 ? _slots_26_io_out_uop_bypassable : _GEN_667 ? _slots_25_io_out_uop_bypassable : _GEN_666 ? _slots_24_io_out_uop_bypassable : _slots_23_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_668 ? _slots_26_io_out_uop_mem_cmd : _GEN_667 ? _slots_25_io_out_uop_mem_cmd : _GEN_666 ? _slots_24_io_out_uop_mem_cmd : _slots_23_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_668 ? _slots_26_io_out_uop_mem_size : _GEN_667 ? _slots_25_io_out_uop_mem_size : _GEN_666 ? _slots_24_io_out_uop_mem_size : _slots_23_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_668 ? _slots_26_io_out_uop_mem_signed : _GEN_667 ? _slots_25_io_out_uop_mem_signed : _GEN_666 ? _slots_24_io_out_uop_mem_signed : _slots_23_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_668 ? _slots_26_io_out_uop_is_fence : _GEN_667 ? _slots_25_io_out_uop_is_fence : _GEN_666 ? _slots_24_io_out_uop_is_fence : _slots_23_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_668 ? _slots_26_io_out_uop_is_amo : _GEN_667 ? _slots_25_io_out_uop_is_amo : _GEN_666 ? _slots_24_io_out_uop_is_amo : _slots_23_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_668 ? _slots_26_io_out_uop_uses_ldq : _GEN_667 ? _slots_25_io_out_uop_uses_ldq : _GEN_666 ? _slots_24_io_out_uop_uses_ldq : _slots_23_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_668 ? _slots_26_io_out_uop_uses_stq : _GEN_667 ? _slots_25_io_out_uop_uses_stq : _GEN_666 ? _slots_24_io_out_uop_uses_stq : _slots_23_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_668 ? _slots_26_io_out_uop_ldst_val : _GEN_667 ? _slots_25_io_out_uop_ldst_val : _GEN_666 ? _slots_24_io_out_uop_ldst_val : _slots_23_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_668 ? _slots_26_io_out_uop_dst_rtype : _GEN_667 ? _slots_25_io_out_uop_dst_rtype : _GEN_666 ? _slots_24_io_out_uop_dst_rtype : _slots_23_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_668 ? _slots_26_io_out_uop_lrs1_rtype : _GEN_667 ? _slots_25_io_out_uop_lrs1_rtype : _GEN_666 ? _slots_24_io_out_uop_lrs1_rtype : _slots_23_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_668 ? _slots_26_io_out_uop_lrs2_rtype : _GEN_667 ? _slots_25_io_out_uop_lrs2_rtype : _GEN_666 ? _slots_24_io_out_uop_lrs2_rtype : _slots_23_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_668 ? _slots_26_io_out_uop_fp_val : _GEN_667 ? _slots_25_io_out_uop_fp_val : _GEN_666 ? _slots_24_io_out_uop_fp_val : _slots_23_io_out_uop_fp_val),
    .io_valid                       (_slots_22_io_valid),
    .io_will_be_valid               (_slots_22_io_will_be_valid),
    .io_request                     (_slots_22_io_request),
    .io_out_uop_uopc                (_slots_22_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_22_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_22_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_22_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_22_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_22_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_22_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_22_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_22_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_22_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_22_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_22_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_22_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_22_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_22_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_22_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_22_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_22_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_22_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_22_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_22_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_22_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_22_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_22_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_22_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_22_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_22_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_22_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_22_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_22_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_22_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_22_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_22_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_22_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_22_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_22_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_22_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_22_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_22_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_22_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_22_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_22_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_22_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_22_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_22_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_22_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_22_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_22_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_22_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_22_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_22_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_22_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_22_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_22_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_22_io_uop_pc_lob),
    .io_uop_taken                   (_slots_22_io_uop_taken),
    .io_uop_imm_packed              (_slots_22_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_22_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_22_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_22_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_22_io_uop_pdst),
    .io_uop_prs1                    (_slots_22_io_uop_prs1),
    .io_uop_prs2                    (_slots_22_io_uop_prs2),
    .io_uop_bypassable              (_slots_22_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_22_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_22_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_22_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_22_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_22_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_22_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_22_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_22_io_uop_fp_val)
  );
  IssueSlot_32 slots_23 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_23_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_65),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_23_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_671 ? _slots_27_io_out_uop_uopc : _GEN_670 ? _slots_26_io_out_uop_uopc : _GEN_669 ? _slots_25_io_out_uop_uopc : _slots_24_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_671 ? _slots_27_io_out_uop_is_rvc : _GEN_670 ? _slots_26_io_out_uop_is_rvc : _GEN_669 ? _slots_25_io_out_uop_is_rvc : _slots_24_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_671 ? _slots_27_io_out_uop_fu_code : _GEN_670 ? _slots_26_io_out_uop_fu_code : _GEN_669 ? _slots_25_io_out_uop_fu_code : _slots_24_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_671 ? _slots_27_io_out_uop_iw_state : _GEN_670 ? _slots_26_io_out_uop_iw_state : _GEN_669 ? _slots_25_io_out_uop_iw_state : _slots_24_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_671 ? _slots_27_io_out_uop_iw_p1_poisoned : _GEN_670 ? _slots_26_io_out_uop_iw_p1_poisoned : _GEN_669 ? _slots_25_io_out_uop_iw_p1_poisoned : _slots_24_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_671 ? _slots_27_io_out_uop_iw_p2_poisoned : _GEN_670 ? _slots_26_io_out_uop_iw_p2_poisoned : _GEN_669 ? _slots_25_io_out_uop_iw_p2_poisoned : _slots_24_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_671 ? _slots_27_io_out_uop_is_br : _GEN_670 ? _slots_26_io_out_uop_is_br : _GEN_669 ? _slots_25_io_out_uop_is_br : _slots_24_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_671 ? _slots_27_io_out_uop_is_jalr : _GEN_670 ? _slots_26_io_out_uop_is_jalr : _GEN_669 ? _slots_25_io_out_uop_is_jalr : _slots_24_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_671 ? _slots_27_io_out_uop_is_jal : _GEN_670 ? _slots_26_io_out_uop_is_jal : _GEN_669 ? _slots_25_io_out_uop_is_jal : _slots_24_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_671 ? _slots_27_io_out_uop_is_sfb : _GEN_670 ? _slots_26_io_out_uop_is_sfb : _GEN_669 ? _slots_25_io_out_uop_is_sfb : _slots_24_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_671 ? _slots_27_io_out_uop_br_mask : _GEN_670 ? _slots_26_io_out_uop_br_mask : _GEN_669 ? _slots_25_io_out_uop_br_mask : _slots_24_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_671 ? _slots_27_io_out_uop_br_tag : _GEN_670 ? _slots_26_io_out_uop_br_tag : _GEN_669 ? _slots_25_io_out_uop_br_tag : _slots_24_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_671 ? _slots_27_io_out_uop_ftq_idx : _GEN_670 ? _slots_26_io_out_uop_ftq_idx : _GEN_669 ? _slots_25_io_out_uop_ftq_idx : _slots_24_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_671 ? _slots_27_io_out_uop_edge_inst : _GEN_670 ? _slots_26_io_out_uop_edge_inst : _GEN_669 ? _slots_25_io_out_uop_edge_inst : _slots_24_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_671 ? _slots_27_io_out_uop_pc_lob : _GEN_670 ? _slots_26_io_out_uop_pc_lob : _GEN_669 ? _slots_25_io_out_uop_pc_lob : _slots_24_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_671 ? _slots_27_io_out_uop_taken : _GEN_670 ? _slots_26_io_out_uop_taken : _GEN_669 ? _slots_25_io_out_uop_taken : _slots_24_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_671 ? _slots_27_io_out_uop_imm_packed : _GEN_670 ? _slots_26_io_out_uop_imm_packed : _GEN_669 ? _slots_25_io_out_uop_imm_packed : _slots_24_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_671 ? _slots_27_io_out_uop_rob_idx : _GEN_670 ? _slots_26_io_out_uop_rob_idx : _GEN_669 ? _slots_25_io_out_uop_rob_idx : _slots_24_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_671 ? _slots_27_io_out_uop_ldq_idx : _GEN_670 ? _slots_26_io_out_uop_ldq_idx : _GEN_669 ? _slots_25_io_out_uop_ldq_idx : _slots_24_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_671 ? _slots_27_io_out_uop_stq_idx : _GEN_670 ? _slots_26_io_out_uop_stq_idx : _GEN_669 ? _slots_25_io_out_uop_stq_idx : _slots_24_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_671 ? _slots_27_io_out_uop_pdst : _GEN_670 ? _slots_26_io_out_uop_pdst : _GEN_669 ? _slots_25_io_out_uop_pdst : _slots_24_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_671 ? _slots_27_io_out_uop_prs1 : _GEN_670 ? _slots_26_io_out_uop_prs1 : _GEN_669 ? _slots_25_io_out_uop_prs1 : _slots_24_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_671 ? _slots_27_io_out_uop_prs2 : _GEN_670 ? _slots_26_io_out_uop_prs2 : _GEN_669 ? _slots_25_io_out_uop_prs2 : _slots_24_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_671 ? _slots_27_io_out_uop_prs3 : _GEN_670 ? _slots_26_io_out_uop_prs3 : _GEN_669 ? _slots_25_io_out_uop_prs3 : _slots_24_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_671 ? _slots_27_io_out_uop_prs1_busy : _GEN_670 ? _slots_26_io_out_uop_prs1_busy : _GEN_669 ? _slots_25_io_out_uop_prs1_busy : _slots_24_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_671 ? _slots_27_io_out_uop_prs2_busy : _GEN_670 ? _slots_26_io_out_uop_prs2_busy : _GEN_669 ? _slots_25_io_out_uop_prs2_busy : _slots_24_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_671 ? _slots_27_io_out_uop_prs3_busy : _GEN_670 ? _slots_26_io_out_uop_prs3_busy : _GEN_669 ? _slots_25_io_out_uop_prs3_busy : _slots_24_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_671 ? _slots_27_io_out_uop_ppred_busy : _GEN_670 ? _slots_26_io_out_uop_ppred_busy : _GEN_669 ? _slots_25_io_out_uop_ppred_busy : _slots_24_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_671 ? _slots_27_io_out_uop_bypassable : _GEN_670 ? _slots_26_io_out_uop_bypassable : _GEN_669 ? _slots_25_io_out_uop_bypassable : _slots_24_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_671 ? _slots_27_io_out_uop_mem_cmd : _GEN_670 ? _slots_26_io_out_uop_mem_cmd : _GEN_669 ? _slots_25_io_out_uop_mem_cmd : _slots_24_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_671 ? _slots_27_io_out_uop_mem_size : _GEN_670 ? _slots_26_io_out_uop_mem_size : _GEN_669 ? _slots_25_io_out_uop_mem_size : _slots_24_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_671 ? _slots_27_io_out_uop_mem_signed : _GEN_670 ? _slots_26_io_out_uop_mem_signed : _GEN_669 ? _slots_25_io_out_uop_mem_signed : _slots_24_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_671 ? _slots_27_io_out_uop_is_fence : _GEN_670 ? _slots_26_io_out_uop_is_fence : _GEN_669 ? _slots_25_io_out_uop_is_fence : _slots_24_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_671 ? _slots_27_io_out_uop_is_amo : _GEN_670 ? _slots_26_io_out_uop_is_amo : _GEN_669 ? _slots_25_io_out_uop_is_amo : _slots_24_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_671 ? _slots_27_io_out_uop_uses_ldq : _GEN_670 ? _slots_26_io_out_uop_uses_ldq : _GEN_669 ? _slots_25_io_out_uop_uses_ldq : _slots_24_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_671 ? _slots_27_io_out_uop_uses_stq : _GEN_670 ? _slots_26_io_out_uop_uses_stq : _GEN_669 ? _slots_25_io_out_uop_uses_stq : _slots_24_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_671 ? _slots_27_io_out_uop_ldst_val : _GEN_670 ? _slots_26_io_out_uop_ldst_val : _GEN_669 ? _slots_25_io_out_uop_ldst_val : _slots_24_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_671 ? _slots_27_io_out_uop_dst_rtype : _GEN_670 ? _slots_26_io_out_uop_dst_rtype : _GEN_669 ? _slots_25_io_out_uop_dst_rtype : _slots_24_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_671 ? _slots_27_io_out_uop_lrs1_rtype : _GEN_670 ? _slots_26_io_out_uop_lrs1_rtype : _GEN_669 ? _slots_25_io_out_uop_lrs1_rtype : _slots_24_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_671 ? _slots_27_io_out_uop_lrs2_rtype : _GEN_670 ? _slots_26_io_out_uop_lrs2_rtype : _GEN_669 ? _slots_25_io_out_uop_lrs2_rtype : _slots_24_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_671 ? _slots_27_io_out_uop_fp_val : _GEN_670 ? _slots_26_io_out_uop_fp_val : _GEN_669 ? _slots_25_io_out_uop_fp_val : _slots_24_io_out_uop_fp_val),
    .io_valid                       (_slots_23_io_valid),
    .io_will_be_valid               (_slots_23_io_will_be_valid),
    .io_request                     (_slots_23_io_request),
    .io_out_uop_uopc                (_slots_23_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_23_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_23_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_23_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_23_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_23_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_23_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_23_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_23_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_23_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_23_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_23_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_23_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_23_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_23_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_23_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_23_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_23_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_23_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_23_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_23_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_23_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_23_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_23_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_23_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_23_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_23_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_23_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_23_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_23_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_23_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_23_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_23_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_23_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_23_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_23_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_23_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_23_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_23_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_23_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_23_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_23_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_23_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_23_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_23_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_23_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_23_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_23_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_23_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_23_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_23_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_23_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_23_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_23_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_23_io_uop_pc_lob),
    .io_uop_taken                   (_slots_23_io_uop_taken),
    .io_uop_imm_packed              (_slots_23_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_23_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_23_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_23_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_23_io_uop_pdst),
    .io_uop_prs1                    (_slots_23_io_uop_prs1),
    .io_uop_prs2                    (_slots_23_io_uop_prs2),
    .io_uop_bypassable              (_slots_23_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_23_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_23_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_23_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_23_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_23_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_23_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_23_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_23_io_uop_fp_val)
  );
  IssueSlot_32 slots_24 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_24_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_67),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_24_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_674 ? _slots_28_io_out_uop_uopc : _GEN_673 ? _slots_27_io_out_uop_uopc : _GEN_672 ? _slots_26_io_out_uop_uopc : _slots_25_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_674 ? _slots_28_io_out_uop_is_rvc : _GEN_673 ? _slots_27_io_out_uop_is_rvc : _GEN_672 ? _slots_26_io_out_uop_is_rvc : _slots_25_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_674 ? _slots_28_io_out_uop_fu_code : _GEN_673 ? _slots_27_io_out_uop_fu_code : _GEN_672 ? _slots_26_io_out_uop_fu_code : _slots_25_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_674 ? _slots_28_io_out_uop_iw_state : _GEN_673 ? _slots_27_io_out_uop_iw_state : _GEN_672 ? _slots_26_io_out_uop_iw_state : _slots_25_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_674 ? _slots_28_io_out_uop_iw_p1_poisoned : _GEN_673 ? _slots_27_io_out_uop_iw_p1_poisoned : _GEN_672 ? _slots_26_io_out_uop_iw_p1_poisoned : _slots_25_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_674 ? _slots_28_io_out_uop_iw_p2_poisoned : _GEN_673 ? _slots_27_io_out_uop_iw_p2_poisoned : _GEN_672 ? _slots_26_io_out_uop_iw_p2_poisoned : _slots_25_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_674 ? _slots_28_io_out_uop_is_br : _GEN_673 ? _slots_27_io_out_uop_is_br : _GEN_672 ? _slots_26_io_out_uop_is_br : _slots_25_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_674 ? _slots_28_io_out_uop_is_jalr : _GEN_673 ? _slots_27_io_out_uop_is_jalr : _GEN_672 ? _slots_26_io_out_uop_is_jalr : _slots_25_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_674 ? _slots_28_io_out_uop_is_jal : _GEN_673 ? _slots_27_io_out_uop_is_jal : _GEN_672 ? _slots_26_io_out_uop_is_jal : _slots_25_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_674 ? _slots_28_io_out_uop_is_sfb : _GEN_673 ? _slots_27_io_out_uop_is_sfb : _GEN_672 ? _slots_26_io_out_uop_is_sfb : _slots_25_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_674 ? _slots_28_io_out_uop_br_mask : _GEN_673 ? _slots_27_io_out_uop_br_mask : _GEN_672 ? _slots_26_io_out_uop_br_mask : _slots_25_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_674 ? _slots_28_io_out_uop_br_tag : _GEN_673 ? _slots_27_io_out_uop_br_tag : _GEN_672 ? _slots_26_io_out_uop_br_tag : _slots_25_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_674 ? _slots_28_io_out_uop_ftq_idx : _GEN_673 ? _slots_27_io_out_uop_ftq_idx : _GEN_672 ? _slots_26_io_out_uop_ftq_idx : _slots_25_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_674 ? _slots_28_io_out_uop_edge_inst : _GEN_673 ? _slots_27_io_out_uop_edge_inst : _GEN_672 ? _slots_26_io_out_uop_edge_inst : _slots_25_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_674 ? _slots_28_io_out_uop_pc_lob : _GEN_673 ? _slots_27_io_out_uop_pc_lob : _GEN_672 ? _slots_26_io_out_uop_pc_lob : _slots_25_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_674 ? _slots_28_io_out_uop_taken : _GEN_673 ? _slots_27_io_out_uop_taken : _GEN_672 ? _slots_26_io_out_uop_taken : _slots_25_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_674 ? _slots_28_io_out_uop_imm_packed : _GEN_673 ? _slots_27_io_out_uop_imm_packed : _GEN_672 ? _slots_26_io_out_uop_imm_packed : _slots_25_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_674 ? _slots_28_io_out_uop_rob_idx : _GEN_673 ? _slots_27_io_out_uop_rob_idx : _GEN_672 ? _slots_26_io_out_uop_rob_idx : _slots_25_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_674 ? _slots_28_io_out_uop_ldq_idx : _GEN_673 ? _slots_27_io_out_uop_ldq_idx : _GEN_672 ? _slots_26_io_out_uop_ldq_idx : _slots_25_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_674 ? _slots_28_io_out_uop_stq_idx : _GEN_673 ? _slots_27_io_out_uop_stq_idx : _GEN_672 ? _slots_26_io_out_uop_stq_idx : _slots_25_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_674 ? _slots_28_io_out_uop_pdst : _GEN_673 ? _slots_27_io_out_uop_pdst : _GEN_672 ? _slots_26_io_out_uop_pdst : _slots_25_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_674 ? _slots_28_io_out_uop_prs1 : _GEN_673 ? _slots_27_io_out_uop_prs1 : _GEN_672 ? _slots_26_io_out_uop_prs1 : _slots_25_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_674 ? _slots_28_io_out_uop_prs2 : _GEN_673 ? _slots_27_io_out_uop_prs2 : _GEN_672 ? _slots_26_io_out_uop_prs2 : _slots_25_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_674 ? _slots_28_io_out_uop_prs3 : _GEN_673 ? _slots_27_io_out_uop_prs3 : _GEN_672 ? _slots_26_io_out_uop_prs3 : _slots_25_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_674 ? _slots_28_io_out_uop_prs1_busy : _GEN_673 ? _slots_27_io_out_uop_prs1_busy : _GEN_672 ? _slots_26_io_out_uop_prs1_busy : _slots_25_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_674 ? _slots_28_io_out_uop_prs2_busy : _GEN_673 ? _slots_27_io_out_uop_prs2_busy : _GEN_672 ? _slots_26_io_out_uop_prs2_busy : _slots_25_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_674 ? _slots_28_io_out_uop_prs3_busy : _GEN_673 ? _slots_27_io_out_uop_prs3_busy : _GEN_672 ? _slots_26_io_out_uop_prs3_busy : _slots_25_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_674 ? _slots_28_io_out_uop_ppred_busy : _GEN_673 ? _slots_27_io_out_uop_ppred_busy : _GEN_672 ? _slots_26_io_out_uop_ppred_busy : _slots_25_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_674 ? _slots_28_io_out_uop_bypassable : _GEN_673 ? _slots_27_io_out_uop_bypassable : _GEN_672 ? _slots_26_io_out_uop_bypassable : _slots_25_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_674 ? _slots_28_io_out_uop_mem_cmd : _GEN_673 ? _slots_27_io_out_uop_mem_cmd : _GEN_672 ? _slots_26_io_out_uop_mem_cmd : _slots_25_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_674 ? _slots_28_io_out_uop_mem_size : _GEN_673 ? _slots_27_io_out_uop_mem_size : _GEN_672 ? _slots_26_io_out_uop_mem_size : _slots_25_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_674 ? _slots_28_io_out_uop_mem_signed : _GEN_673 ? _slots_27_io_out_uop_mem_signed : _GEN_672 ? _slots_26_io_out_uop_mem_signed : _slots_25_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_674 ? _slots_28_io_out_uop_is_fence : _GEN_673 ? _slots_27_io_out_uop_is_fence : _GEN_672 ? _slots_26_io_out_uop_is_fence : _slots_25_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_674 ? _slots_28_io_out_uop_is_amo : _GEN_673 ? _slots_27_io_out_uop_is_amo : _GEN_672 ? _slots_26_io_out_uop_is_amo : _slots_25_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_674 ? _slots_28_io_out_uop_uses_ldq : _GEN_673 ? _slots_27_io_out_uop_uses_ldq : _GEN_672 ? _slots_26_io_out_uop_uses_ldq : _slots_25_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_674 ? _slots_28_io_out_uop_uses_stq : _GEN_673 ? _slots_27_io_out_uop_uses_stq : _GEN_672 ? _slots_26_io_out_uop_uses_stq : _slots_25_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_674 ? _slots_28_io_out_uop_ldst_val : _GEN_673 ? _slots_27_io_out_uop_ldst_val : _GEN_672 ? _slots_26_io_out_uop_ldst_val : _slots_25_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_674 ? _slots_28_io_out_uop_dst_rtype : _GEN_673 ? _slots_27_io_out_uop_dst_rtype : _GEN_672 ? _slots_26_io_out_uop_dst_rtype : _slots_25_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_674 ? _slots_28_io_out_uop_lrs1_rtype : _GEN_673 ? _slots_27_io_out_uop_lrs1_rtype : _GEN_672 ? _slots_26_io_out_uop_lrs1_rtype : _slots_25_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_674 ? _slots_28_io_out_uop_lrs2_rtype : _GEN_673 ? _slots_27_io_out_uop_lrs2_rtype : _GEN_672 ? _slots_26_io_out_uop_lrs2_rtype : _slots_25_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_674 ? _slots_28_io_out_uop_fp_val : _GEN_673 ? _slots_27_io_out_uop_fp_val : _GEN_672 ? _slots_26_io_out_uop_fp_val : _slots_25_io_out_uop_fp_val),
    .io_valid                       (_slots_24_io_valid),
    .io_will_be_valid               (_slots_24_io_will_be_valid),
    .io_request                     (_slots_24_io_request),
    .io_out_uop_uopc                (_slots_24_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_24_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_24_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_24_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_24_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_24_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_24_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_24_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_24_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_24_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_24_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_24_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_24_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_24_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_24_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_24_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_24_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_24_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_24_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_24_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_24_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_24_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_24_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_24_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_24_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_24_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_24_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_24_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_24_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_24_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_24_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_24_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_24_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_24_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_24_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_24_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_24_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_24_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_24_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_24_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_24_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_24_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_24_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_24_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_24_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_24_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_24_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_24_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_24_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_24_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_24_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_24_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_24_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_24_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_24_io_uop_pc_lob),
    .io_uop_taken                   (_slots_24_io_uop_taken),
    .io_uop_imm_packed              (_slots_24_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_24_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_24_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_24_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_24_io_uop_pdst),
    .io_uop_prs1                    (_slots_24_io_uop_prs1),
    .io_uop_prs2                    (_slots_24_io_uop_prs2),
    .io_uop_bypassable              (_slots_24_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_24_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_24_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_24_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_24_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_24_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_24_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_24_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_24_io_uop_fp_val)
  );
  IssueSlot_32 slots_25 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_25_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_69),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_25_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_677 ? _slots_29_io_out_uop_uopc : _GEN_676 ? _slots_28_io_out_uop_uopc : _GEN_675 ? _slots_27_io_out_uop_uopc : _slots_26_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_677 ? _slots_29_io_out_uop_is_rvc : _GEN_676 ? _slots_28_io_out_uop_is_rvc : _GEN_675 ? _slots_27_io_out_uop_is_rvc : _slots_26_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_677 ? _slots_29_io_out_uop_fu_code : _GEN_676 ? _slots_28_io_out_uop_fu_code : _GEN_675 ? _slots_27_io_out_uop_fu_code : _slots_26_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_677 ? _slots_29_io_out_uop_iw_state : _GEN_676 ? _slots_28_io_out_uop_iw_state : _GEN_675 ? _slots_27_io_out_uop_iw_state : _slots_26_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_677 ? _slots_29_io_out_uop_iw_p1_poisoned : _GEN_676 ? _slots_28_io_out_uop_iw_p1_poisoned : _GEN_675 ? _slots_27_io_out_uop_iw_p1_poisoned : _slots_26_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_677 ? _slots_29_io_out_uop_iw_p2_poisoned : _GEN_676 ? _slots_28_io_out_uop_iw_p2_poisoned : _GEN_675 ? _slots_27_io_out_uop_iw_p2_poisoned : _slots_26_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_677 ? _slots_29_io_out_uop_is_br : _GEN_676 ? _slots_28_io_out_uop_is_br : _GEN_675 ? _slots_27_io_out_uop_is_br : _slots_26_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_677 ? _slots_29_io_out_uop_is_jalr : _GEN_676 ? _slots_28_io_out_uop_is_jalr : _GEN_675 ? _slots_27_io_out_uop_is_jalr : _slots_26_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_677 ? _slots_29_io_out_uop_is_jal : _GEN_676 ? _slots_28_io_out_uop_is_jal : _GEN_675 ? _slots_27_io_out_uop_is_jal : _slots_26_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_677 ? _slots_29_io_out_uop_is_sfb : _GEN_676 ? _slots_28_io_out_uop_is_sfb : _GEN_675 ? _slots_27_io_out_uop_is_sfb : _slots_26_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_677 ? _slots_29_io_out_uop_br_mask : _GEN_676 ? _slots_28_io_out_uop_br_mask : _GEN_675 ? _slots_27_io_out_uop_br_mask : _slots_26_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_677 ? _slots_29_io_out_uop_br_tag : _GEN_676 ? _slots_28_io_out_uop_br_tag : _GEN_675 ? _slots_27_io_out_uop_br_tag : _slots_26_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_677 ? _slots_29_io_out_uop_ftq_idx : _GEN_676 ? _slots_28_io_out_uop_ftq_idx : _GEN_675 ? _slots_27_io_out_uop_ftq_idx : _slots_26_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_677 ? _slots_29_io_out_uop_edge_inst : _GEN_676 ? _slots_28_io_out_uop_edge_inst : _GEN_675 ? _slots_27_io_out_uop_edge_inst : _slots_26_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_677 ? _slots_29_io_out_uop_pc_lob : _GEN_676 ? _slots_28_io_out_uop_pc_lob : _GEN_675 ? _slots_27_io_out_uop_pc_lob : _slots_26_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_677 ? _slots_29_io_out_uop_taken : _GEN_676 ? _slots_28_io_out_uop_taken : _GEN_675 ? _slots_27_io_out_uop_taken : _slots_26_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_677 ? _slots_29_io_out_uop_imm_packed : _GEN_676 ? _slots_28_io_out_uop_imm_packed : _GEN_675 ? _slots_27_io_out_uop_imm_packed : _slots_26_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_677 ? _slots_29_io_out_uop_rob_idx : _GEN_676 ? _slots_28_io_out_uop_rob_idx : _GEN_675 ? _slots_27_io_out_uop_rob_idx : _slots_26_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_677 ? _slots_29_io_out_uop_ldq_idx : _GEN_676 ? _slots_28_io_out_uop_ldq_idx : _GEN_675 ? _slots_27_io_out_uop_ldq_idx : _slots_26_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_677 ? _slots_29_io_out_uop_stq_idx : _GEN_676 ? _slots_28_io_out_uop_stq_idx : _GEN_675 ? _slots_27_io_out_uop_stq_idx : _slots_26_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_677 ? _slots_29_io_out_uop_pdst : _GEN_676 ? _slots_28_io_out_uop_pdst : _GEN_675 ? _slots_27_io_out_uop_pdst : _slots_26_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_677 ? _slots_29_io_out_uop_prs1 : _GEN_676 ? _slots_28_io_out_uop_prs1 : _GEN_675 ? _slots_27_io_out_uop_prs1 : _slots_26_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_677 ? _slots_29_io_out_uop_prs2 : _GEN_676 ? _slots_28_io_out_uop_prs2 : _GEN_675 ? _slots_27_io_out_uop_prs2 : _slots_26_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_677 ? _slots_29_io_out_uop_prs3 : _GEN_676 ? _slots_28_io_out_uop_prs3 : _GEN_675 ? _slots_27_io_out_uop_prs3 : _slots_26_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_677 ? _slots_29_io_out_uop_prs1_busy : _GEN_676 ? _slots_28_io_out_uop_prs1_busy : _GEN_675 ? _slots_27_io_out_uop_prs1_busy : _slots_26_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_677 ? _slots_29_io_out_uop_prs2_busy : _GEN_676 ? _slots_28_io_out_uop_prs2_busy : _GEN_675 ? _slots_27_io_out_uop_prs2_busy : _slots_26_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_677 ? _slots_29_io_out_uop_prs3_busy : _GEN_676 ? _slots_28_io_out_uop_prs3_busy : _GEN_675 ? _slots_27_io_out_uop_prs3_busy : _slots_26_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_677 ? _slots_29_io_out_uop_ppred_busy : _GEN_676 ? _slots_28_io_out_uop_ppred_busy : _GEN_675 ? _slots_27_io_out_uop_ppred_busy : _slots_26_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_677 ? _slots_29_io_out_uop_bypassable : _GEN_676 ? _slots_28_io_out_uop_bypassable : _GEN_675 ? _slots_27_io_out_uop_bypassable : _slots_26_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_677 ? _slots_29_io_out_uop_mem_cmd : _GEN_676 ? _slots_28_io_out_uop_mem_cmd : _GEN_675 ? _slots_27_io_out_uop_mem_cmd : _slots_26_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_677 ? _slots_29_io_out_uop_mem_size : _GEN_676 ? _slots_28_io_out_uop_mem_size : _GEN_675 ? _slots_27_io_out_uop_mem_size : _slots_26_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_677 ? _slots_29_io_out_uop_mem_signed : _GEN_676 ? _slots_28_io_out_uop_mem_signed : _GEN_675 ? _slots_27_io_out_uop_mem_signed : _slots_26_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_677 ? _slots_29_io_out_uop_is_fence : _GEN_676 ? _slots_28_io_out_uop_is_fence : _GEN_675 ? _slots_27_io_out_uop_is_fence : _slots_26_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_677 ? _slots_29_io_out_uop_is_amo : _GEN_676 ? _slots_28_io_out_uop_is_amo : _GEN_675 ? _slots_27_io_out_uop_is_amo : _slots_26_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_677 ? _slots_29_io_out_uop_uses_ldq : _GEN_676 ? _slots_28_io_out_uop_uses_ldq : _GEN_675 ? _slots_27_io_out_uop_uses_ldq : _slots_26_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_677 ? _slots_29_io_out_uop_uses_stq : _GEN_676 ? _slots_28_io_out_uop_uses_stq : _GEN_675 ? _slots_27_io_out_uop_uses_stq : _slots_26_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_677 ? _slots_29_io_out_uop_ldst_val : _GEN_676 ? _slots_28_io_out_uop_ldst_val : _GEN_675 ? _slots_27_io_out_uop_ldst_val : _slots_26_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_677 ? _slots_29_io_out_uop_dst_rtype : _GEN_676 ? _slots_28_io_out_uop_dst_rtype : _GEN_675 ? _slots_27_io_out_uop_dst_rtype : _slots_26_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_677 ? _slots_29_io_out_uop_lrs1_rtype : _GEN_676 ? _slots_28_io_out_uop_lrs1_rtype : _GEN_675 ? _slots_27_io_out_uop_lrs1_rtype : _slots_26_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_677 ? _slots_29_io_out_uop_lrs2_rtype : _GEN_676 ? _slots_28_io_out_uop_lrs2_rtype : _GEN_675 ? _slots_27_io_out_uop_lrs2_rtype : _slots_26_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_677 ? _slots_29_io_out_uop_fp_val : _GEN_676 ? _slots_28_io_out_uop_fp_val : _GEN_675 ? _slots_27_io_out_uop_fp_val : _slots_26_io_out_uop_fp_val),
    .io_valid                       (_slots_25_io_valid),
    .io_will_be_valid               (_slots_25_io_will_be_valid),
    .io_request                     (_slots_25_io_request),
    .io_out_uop_uopc                (_slots_25_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_25_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_25_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_25_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_25_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_25_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_25_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_25_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_25_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_25_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_25_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_25_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_25_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_25_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_25_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_25_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_25_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_25_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_25_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_25_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_25_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_25_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_25_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_25_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_25_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_25_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_25_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_25_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_25_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_25_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_25_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_25_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_25_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_25_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_25_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_25_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_25_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_25_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_25_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_25_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_25_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_25_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_25_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_25_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_25_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_25_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_25_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_25_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_25_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_25_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_25_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_25_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_25_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_25_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_25_io_uop_pc_lob),
    .io_uop_taken                   (_slots_25_io_uop_taken),
    .io_uop_imm_packed              (_slots_25_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_25_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_25_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_25_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_25_io_uop_pdst),
    .io_uop_prs1                    (_slots_25_io_uop_prs1),
    .io_uop_prs2                    (_slots_25_io_uop_prs2),
    .io_uop_bypassable              (_slots_25_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_25_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_25_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_25_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_25_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_25_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_25_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_25_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_25_io_uop_fp_val)
  );
  IssueSlot_32 slots_26 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_26_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_71),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_26_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_680 ? _slots_30_io_out_uop_uopc : _GEN_679 ? _slots_29_io_out_uop_uopc : _GEN_678 ? _slots_28_io_out_uop_uopc : _slots_27_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_680 ? _slots_30_io_out_uop_is_rvc : _GEN_679 ? _slots_29_io_out_uop_is_rvc : _GEN_678 ? _slots_28_io_out_uop_is_rvc : _slots_27_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_680 ? _slots_30_io_out_uop_fu_code : _GEN_679 ? _slots_29_io_out_uop_fu_code : _GEN_678 ? _slots_28_io_out_uop_fu_code : _slots_27_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_680 ? _slots_30_io_out_uop_iw_state : _GEN_679 ? _slots_29_io_out_uop_iw_state : _GEN_678 ? _slots_28_io_out_uop_iw_state : _slots_27_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_680 ? _slots_30_io_out_uop_iw_p1_poisoned : _GEN_679 ? _slots_29_io_out_uop_iw_p1_poisoned : _GEN_678 ? _slots_28_io_out_uop_iw_p1_poisoned : _slots_27_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_680 ? _slots_30_io_out_uop_iw_p2_poisoned : _GEN_679 ? _slots_29_io_out_uop_iw_p2_poisoned : _GEN_678 ? _slots_28_io_out_uop_iw_p2_poisoned : _slots_27_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_680 ? _slots_30_io_out_uop_is_br : _GEN_679 ? _slots_29_io_out_uop_is_br : _GEN_678 ? _slots_28_io_out_uop_is_br : _slots_27_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_680 ? _slots_30_io_out_uop_is_jalr : _GEN_679 ? _slots_29_io_out_uop_is_jalr : _GEN_678 ? _slots_28_io_out_uop_is_jalr : _slots_27_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_680 ? _slots_30_io_out_uop_is_jal : _GEN_679 ? _slots_29_io_out_uop_is_jal : _GEN_678 ? _slots_28_io_out_uop_is_jal : _slots_27_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_680 ? _slots_30_io_out_uop_is_sfb : _GEN_679 ? _slots_29_io_out_uop_is_sfb : _GEN_678 ? _slots_28_io_out_uop_is_sfb : _slots_27_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_680 ? _slots_30_io_out_uop_br_mask : _GEN_679 ? _slots_29_io_out_uop_br_mask : _GEN_678 ? _slots_28_io_out_uop_br_mask : _slots_27_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_680 ? _slots_30_io_out_uop_br_tag : _GEN_679 ? _slots_29_io_out_uop_br_tag : _GEN_678 ? _slots_28_io_out_uop_br_tag : _slots_27_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_680 ? _slots_30_io_out_uop_ftq_idx : _GEN_679 ? _slots_29_io_out_uop_ftq_idx : _GEN_678 ? _slots_28_io_out_uop_ftq_idx : _slots_27_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_680 ? _slots_30_io_out_uop_edge_inst : _GEN_679 ? _slots_29_io_out_uop_edge_inst : _GEN_678 ? _slots_28_io_out_uop_edge_inst : _slots_27_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_680 ? _slots_30_io_out_uop_pc_lob : _GEN_679 ? _slots_29_io_out_uop_pc_lob : _GEN_678 ? _slots_28_io_out_uop_pc_lob : _slots_27_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_680 ? _slots_30_io_out_uop_taken : _GEN_679 ? _slots_29_io_out_uop_taken : _GEN_678 ? _slots_28_io_out_uop_taken : _slots_27_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_680 ? _slots_30_io_out_uop_imm_packed : _GEN_679 ? _slots_29_io_out_uop_imm_packed : _GEN_678 ? _slots_28_io_out_uop_imm_packed : _slots_27_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_680 ? _slots_30_io_out_uop_rob_idx : _GEN_679 ? _slots_29_io_out_uop_rob_idx : _GEN_678 ? _slots_28_io_out_uop_rob_idx : _slots_27_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_680 ? _slots_30_io_out_uop_ldq_idx : _GEN_679 ? _slots_29_io_out_uop_ldq_idx : _GEN_678 ? _slots_28_io_out_uop_ldq_idx : _slots_27_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_680 ? _slots_30_io_out_uop_stq_idx : _GEN_679 ? _slots_29_io_out_uop_stq_idx : _GEN_678 ? _slots_28_io_out_uop_stq_idx : _slots_27_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_680 ? _slots_30_io_out_uop_pdst : _GEN_679 ? _slots_29_io_out_uop_pdst : _GEN_678 ? _slots_28_io_out_uop_pdst : _slots_27_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_680 ? _slots_30_io_out_uop_prs1 : _GEN_679 ? _slots_29_io_out_uop_prs1 : _GEN_678 ? _slots_28_io_out_uop_prs1 : _slots_27_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_680 ? _slots_30_io_out_uop_prs2 : _GEN_679 ? _slots_29_io_out_uop_prs2 : _GEN_678 ? _slots_28_io_out_uop_prs2 : _slots_27_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_680 ? _slots_30_io_out_uop_prs3 : _GEN_679 ? _slots_29_io_out_uop_prs3 : _GEN_678 ? _slots_28_io_out_uop_prs3 : _slots_27_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_680 ? _slots_30_io_out_uop_prs1_busy : _GEN_679 ? _slots_29_io_out_uop_prs1_busy : _GEN_678 ? _slots_28_io_out_uop_prs1_busy : _slots_27_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_680 ? _slots_30_io_out_uop_prs2_busy : _GEN_679 ? _slots_29_io_out_uop_prs2_busy : _GEN_678 ? _slots_28_io_out_uop_prs2_busy : _slots_27_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_680 ? _slots_30_io_out_uop_prs3_busy : _GEN_679 ? _slots_29_io_out_uop_prs3_busy : _GEN_678 ? _slots_28_io_out_uop_prs3_busy : _slots_27_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_680 ? _slots_30_io_out_uop_ppred_busy : _GEN_679 ? _slots_29_io_out_uop_ppred_busy : _GEN_678 ? _slots_28_io_out_uop_ppred_busy : _slots_27_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_680 ? _slots_30_io_out_uop_bypassable : _GEN_679 ? _slots_29_io_out_uop_bypassable : _GEN_678 ? _slots_28_io_out_uop_bypassable : _slots_27_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_680 ? _slots_30_io_out_uop_mem_cmd : _GEN_679 ? _slots_29_io_out_uop_mem_cmd : _GEN_678 ? _slots_28_io_out_uop_mem_cmd : _slots_27_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_680 ? _slots_30_io_out_uop_mem_size : _GEN_679 ? _slots_29_io_out_uop_mem_size : _GEN_678 ? _slots_28_io_out_uop_mem_size : _slots_27_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_680 ? _slots_30_io_out_uop_mem_signed : _GEN_679 ? _slots_29_io_out_uop_mem_signed : _GEN_678 ? _slots_28_io_out_uop_mem_signed : _slots_27_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_680 ? _slots_30_io_out_uop_is_fence : _GEN_679 ? _slots_29_io_out_uop_is_fence : _GEN_678 ? _slots_28_io_out_uop_is_fence : _slots_27_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_680 ? _slots_30_io_out_uop_is_amo : _GEN_679 ? _slots_29_io_out_uop_is_amo : _GEN_678 ? _slots_28_io_out_uop_is_amo : _slots_27_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_680 ? _slots_30_io_out_uop_uses_ldq : _GEN_679 ? _slots_29_io_out_uop_uses_ldq : _GEN_678 ? _slots_28_io_out_uop_uses_ldq : _slots_27_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_680 ? _slots_30_io_out_uop_uses_stq : _GEN_679 ? _slots_29_io_out_uop_uses_stq : _GEN_678 ? _slots_28_io_out_uop_uses_stq : _slots_27_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_680 ? _slots_30_io_out_uop_ldst_val : _GEN_679 ? _slots_29_io_out_uop_ldst_val : _GEN_678 ? _slots_28_io_out_uop_ldst_val : _slots_27_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_680 ? _slots_30_io_out_uop_dst_rtype : _GEN_679 ? _slots_29_io_out_uop_dst_rtype : _GEN_678 ? _slots_28_io_out_uop_dst_rtype : _slots_27_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_680 ? _slots_30_io_out_uop_lrs1_rtype : _GEN_679 ? _slots_29_io_out_uop_lrs1_rtype : _GEN_678 ? _slots_28_io_out_uop_lrs1_rtype : _slots_27_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_680 ? _slots_30_io_out_uop_lrs2_rtype : _GEN_679 ? _slots_29_io_out_uop_lrs2_rtype : _GEN_678 ? _slots_28_io_out_uop_lrs2_rtype : _slots_27_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_680 ? _slots_30_io_out_uop_fp_val : _GEN_679 ? _slots_29_io_out_uop_fp_val : _GEN_678 ? _slots_28_io_out_uop_fp_val : _slots_27_io_out_uop_fp_val),
    .io_valid                       (_slots_26_io_valid),
    .io_will_be_valid               (_slots_26_io_will_be_valid),
    .io_request                     (_slots_26_io_request),
    .io_out_uop_uopc                (_slots_26_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_26_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_26_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_26_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_26_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_26_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_26_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_26_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_26_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_26_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_26_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_26_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_26_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_26_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_26_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_26_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_26_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_26_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_26_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_26_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_26_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_26_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_26_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_26_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_26_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_26_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_26_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_26_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_26_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_26_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_26_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_26_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_26_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_26_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_26_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_26_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_26_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_26_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_26_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_26_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_26_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_26_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_26_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_26_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_26_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_26_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_26_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_26_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_26_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_26_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_26_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_26_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_26_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_26_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_26_io_uop_pc_lob),
    .io_uop_taken                   (_slots_26_io_uop_taken),
    .io_uop_imm_packed              (_slots_26_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_26_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_26_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_26_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_26_io_uop_pdst),
    .io_uop_prs1                    (_slots_26_io_uop_prs1),
    .io_uop_prs2                    (_slots_26_io_uop_prs2),
    .io_uop_bypassable              (_slots_26_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_26_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_26_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_26_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_26_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_26_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_26_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_26_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_26_io_uop_fp_val)
  );
  IssueSlot_32 slots_27 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_27_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_73),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_27_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_683 ? _slots_31_io_out_uop_uopc : _GEN_682 ? _slots_30_io_out_uop_uopc : _GEN_681 ? _slots_29_io_out_uop_uopc : _slots_28_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_683 ? _slots_31_io_out_uop_is_rvc : _GEN_682 ? _slots_30_io_out_uop_is_rvc : _GEN_681 ? _slots_29_io_out_uop_is_rvc : _slots_28_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_683 ? _slots_31_io_out_uop_fu_code : _GEN_682 ? _slots_30_io_out_uop_fu_code : _GEN_681 ? _slots_29_io_out_uop_fu_code : _slots_28_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_683 ? _slots_31_io_out_uop_iw_state : _GEN_682 ? _slots_30_io_out_uop_iw_state : _GEN_681 ? _slots_29_io_out_uop_iw_state : _slots_28_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_683 ? _slots_31_io_out_uop_iw_p1_poisoned : _GEN_682 ? _slots_30_io_out_uop_iw_p1_poisoned : _GEN_681 ? _slots_29_io_out_uop_iw_p1_poisoned : _slots_28_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_683 ? _slots_31_io_out_uop_iw_p2_poisoned : _GEN_682 ? _slots_30_io_out_uop_iw_p2_poisoned : _GEN_681 ? _slots_29_io_out_uop_iw_p2_poisoned : _slots_28_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_683 ? _slots_31_io_out_uop_is_br : _GEN_682 ? _slots_30_io_out_uop_is_br : _GEN_681 ? _slots_29_io_out_uop_is_br : _slots_28_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_683 ? _slots_31_io_out_uop_is_jalr : _GEN_682 ? _slots_30_io_out_uop_is_jalr : _GEN_681 ? _slots_29_io_out_uop_is_jalr : _slots_28_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_683 ? _slots_31_io_out_uop_is_jal : _GEN_682 ? _slots_30_io_out_uop_is_jal : _GEN_681 ? _slots_29_io_out_uop_is_jal : _slots_28_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_683 ? _slots_31_io_out_uop_is_sfb : _GEN_682 ? _slots_30_io_out_uop_is_sfb : _GEN_681 ? _slots_29_io_out_uop_is_sfb : _slots_28_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_683 ? _slots_31_io_out_uop_br_mask : _GEN_682 ? _slots_30_io_out_uop_br_mask : _GEN_681 ? _slots_29_io_out_uop_br_mask : _slots_28_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_683 ? _slots_31_io_out_uop_br_tag : _GEN_682 ? _slots_30_io_out_uop_br_tag : _GEN_681 ? _slots_29_io_out_uop_br_tag : _slots_28_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_683 ? _slots_31_io_out_uop_ftq_idx : _GEN_682 ? _slots_30_io_out_uop_ftq_idx : _GEN_681 ? _slots_29_io_out_uop_ftq_idx : _slots_28_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_683 ? _slots_31_io_out_uop_edge_inst : _GEN_682 ? _slots_30_io_out_uop_edge_inst : _GEN_681 ? _slots_29_io_out_uop_edge_inst : _slots_28_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_683 ? _slots_31_io_out_uop_pc_lob : _GEN_682 ? _slots_30_io_out_uop_pc_lob : _GEN_681 ? _slots_29_io_out_uop_pc_lob : _slots_28_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_683 ? _slots_31_io_out_uop_taken : _GEN_682 ? _slots_30_io_out_uop_taken : _GEN_681 ? _slots_29_io_out_uop_taken : _slots_28_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_683 ? _slots_31_io_out_uop_imm_packed : _GEN_682 ? _slots_30_io_out_uop_imm_packed : _GEN_681 ? _slots_29_io_out_uop_imm_packed : _slots_28_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_683 ? _slots_31_io_out_uop_rob_idx : _GEN_682 ? _slots_30_io_out_uop_rob_idx : _GEN_681 ? _slots_29_io_out_uop_rob_idx : _slots_28_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_683 ? _slots_31_io_out_uop_ldq_idx : _GEN_682 ? _slots_30_io_out_uop_ldq_idx : _GEN_681 ? _slots_29_io_out_uop_ldq_idx : _slots_28_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_683 ? _slots_31_io_out_uop_stq_idx : _GEN_682 ? _slots_30_io_out_uop_stq_idx : _GEN_681 ? _slots_29_io_out_uop_stq_idx : _slots_28_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_683 ? _slots_31_io_out_uop_pdst : _GEN_682 ? _slots_30_io_out_uop_pdst : _GEN_681 ? _slots_29_io_out_uop_pdst : _slots_28_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_683 ? _slots_31_io_out_uop_prs1 : _GEN_682 ? _slots_30_io_out_uop_prs1 : _GEN_681 ? _slots_29_io_out_uop_prs1 : _slots_28_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_683 ? _slots_31_io_out_uop_prs2 : _GEN_682 ? _slots_30_io_out_uop_prs2 : _GEN_681 ? _slots_29_io_out_uop_prs2 : _slots_28_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_683 ? _slots_31_io_out_uop_prs3 : _GEN_682 ? _slots_30_io_out_uop_prs3 : _GEN_681 ? _slots_29_io_out_uop_prs3 : _slots_28_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_683 ? _slots_31_io_out_uop_prs1_busy : _GEN_682 ? _slots_30_io_out_uop_prs1_busy : _GEN_681 ? _slots_29_io_out_uop_prs1_busy : _slots_28_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_683 ? _slots_31_io_out_uop_prs2_busy : _GEN_682 ? _slots_30_io_out_uop_prs2_busy : _GEN_681 ? _slots_29_io_out_uop_prs2_busy : _slots_28_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_683 ? _slots_31_io_out_uop_prs3_busy : _GEN_682 ? _slots_30_io_out_uop_prs3_busy : _GEN_681 ? _slots_29_io_out_uop_prs3_busy : _slots_28_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_683 ? _slots_31_io_out_uop_ppred_busy : _GEN_682 ? _slots_30_io_out_uop_ppred_busy : _GEN_681 ? _slots_29_io_out_uop_ppred_busy : _slots_28_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_683 ? _slots_31_io_out_uop_bypassable : _GEN_682 ? _slots_30_io_out_uop_bypassable : _GEN_681 ? _slots_29_io_out_uop_bypassable : _slots_28_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_683 ? _slots_31_io_out_uop_mem_cmd : _GEN_682 ? _slots_30_io_out_uop_mem_cmd : _GEN_681 ? _slots_29_io_out_uop_mem_cmd : _slots_28_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_683 ? _slots_31_io_out_uop_mem_size : _GEN_682 ? _slots_30_io_out_uop_mem_size : _GEN_681 ? _slots_29_io_out_uop_mem_size : _slots_28_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_683 ? _slots_31_io_out_uop_mem_signed : _GEN_682 ? _slots_30_io_out_uop_mem_signed : _GEN_681 ? _slots_29_io_out_uop_mem_signed : _slots_28_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_683 ? _slots_31_io_out_uop_is_fence : _GEN_682 ? _slots_30_io_out_uop_is_fence : _GEN_681 ? _slots_29_io_out_uop_is_fence : _slots_28_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_683 ? _slots_31_io_out_uop_is_amo : _GEN_682 ? _slots_30_io_out_uop_is_amo : _GEN_681 ? _slots_29_io_out_uop_is_amo : _slots_28_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_683 ? _slots_31_io_out_uop_uses_ldq : _GEN_682 ? _slots_30_io_out_uop_uses_ldq : _GEN_681 ? _slots_29_io_out_uop_uses_ldq : _slots_28_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_683 ? _slots_31_io_out_uop_uses_stq : _GEN_682 ? _slots_30_io_out_uop_uses_stq : _GEN_681 ? _slots_29_io_out_uop_uses_stq : _slots_28_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_683 ? _slots_31_io_out_uop_ldst_val : _GEN_682 ? _slots_30_io_out_uop_ldst_val : _GEN_681 ? _slots_29_io_out_uop_ldst_val : _slots_28_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_683 ? _slots_31_io_out_uop_dst_rtype : _GEN_682 ? _slots_30_io_out_uop_dst_rtype : _GEN_681 ? _slots_29_io_out_uop_dst_rtype : _slots_28_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_683 ? _slots_31_io_out_uop_lrs1_rtype : _GEN_682 ? _slots_30_io_out_uop_lrs1_rtype : _GEN_681 ? _slots_29_io_out_uop_lrs1_rtype : _slots_28_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_683 ? _slots_31_io_out_uop_lrs2_rtype : _GEN_682 ? _slots_30_io_out_uop_lrs2_rtype : _GEN_681 ? _slots_29_io_out_uop_lrs2_rtype : _slots_28_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_683 ? _slots_31_io_out_uop_fp_val : _GEN_682 ? _slots_30_io_out_uop_fp_val : _GEN_681 ? _slots_29_io_out_uop_fp_val : _slots_28_io_out_uop_fp_val),
    .io_valid                       (_slots_27_io_valid),
    .io_will_be_valid               (_slots_27_io_will_be_valid),
    .io_request                     (_slots_27_io_request),
    .io_out_uop_uopc                (_slots_27_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_27_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_27_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_27_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_27_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_27_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_27_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_27_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_27_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_27_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_27_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_27_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_27_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_27_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_27_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_27_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_27_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_27_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_27_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_27_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_27_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_27_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_27_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_27_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_27_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_27_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_27_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_27_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_27_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_27_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_27_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_27_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_27_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_27_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_27_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_27_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_27_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_27_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_27_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_27_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_27_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_27_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_27_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_27_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_27_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_27_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_27_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_27_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_27_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_27_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_27_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_27_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_27_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_27_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_27_io_uop_pc_lob),
    .io_uop_taken                   (_slots_27_io_uop_taken),
    .io_uop_imm_packed              (_slots_27_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_27_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_27_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_27_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_27_io_uop_pdst),
    .io_uop_prs1                    (_slots_27_io_uop_prs1),
    .io_uop_prs2                    (_slots_27_io_uop_prs2),
    .io_uop_bypassable              (_slots_27_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_27_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_27_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_27_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_27_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_27_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_27_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_27_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_27_io_uop_fp_val)
  );
  IssueSlot_32 slots_28 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_28_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_75),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_28_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_686 ? _slots_32_io_out_uop_uopc : _GEN_685 ? _slots_31_io_out_uop_uopc : _GEN_684 ? _slots_30_io_out_uop_uopc : _slots_29_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_686 ? _slots_32_io_out_uop_is_rvc : _GEN_685 ? _slots_31_io_out_uop_is_rvc : _GEN_684 ? _slots_30_io_out_uop_is_rvc : _slots_29_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_686 ? _slots_32_io_out_uop_fu_code : _GEN_685 ? _slots_31_io_out_uop_fu_code : _GEN_684 ? _slots_30_io_out_uop_fu_code : _slots_29_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_686 ? _slots_32_io_out_uop_iw_state : _GEN_685 ? _slots_31_io_out_uop_iw_state : _GEN_684 ? _slots_30_io_out_uop_iw_state : _slots_29_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_686 ? _slots_32_io_out_uop_iw_p1_poisoned : _GEN_685 ? _slots_31_io_out_uop_iw_p1_poisoned : _GEN_684 ? _slots_30_io_out_uop_iw_p1_poisoned : _slots_29_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_686 ? _slots_32_io_out_uop_iw_p2_poisoned : _GEN_685 ? _slots_31_io_out_uop_iw_p2_poisoned : _GEN_684 ? _slots_30_io_out_uop_iw_p2_poisoned : _slots_29_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_686 ? _slots_32_io_out_uop_is_br : _GEN_685 ? _slots_31_io_out_uop_is_br : _GEN_684 ? _slots_30_io_out_uop_is_br : _slots_29_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_686 ? _slots_32_io_out_uop_is_jalr : _GEN_685 ? _slots_31_io_out_uop_is_jalr : _GEN_684 ? _slots_30_io_out_uop_is_jalr : _slots_29_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_686 ? _slots_32_io_out_uop_is_jal : _GEN_685 ? _slots_31_io_out_uop_is_jal : _GEN_684 ? _slots_30_io_out_uop_is_jal : _slots_29_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_686 ? _slots_32_io_out_uop_is_sfb : _GEN_685 ? _slots_31_io_out_uop_is_sfb : _GEN_684 ? _slots_30_io_out_uop_is_sfb : _slots_29_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_686 ? _slots_32_io_out_uop_br_mask : _GEN_685 ? _slots_31_io_out_uop_br_mask : _GEN_684 ? _slots_30_io_out_uop_br_mask : _slots_29_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_686 ? _slots_32_io_out_uop_br_tag : _GEN_685 ? _slots_31_io_out_uop_br_tag : _GEN_684 ? _slots_30_io_out_uop_br_tag : _slots_29_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_686 ? _slots_32_io_out_uop_ftq_idx : _GEN_685 ? _slots_31_io_out_uop_ftq_idx : _GEN_684 ? _slots_30_io_out_uop_ftq_idx : _slots_29_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_686 ? _slots_32_io_out_uop_edge_inst : _GEN_685 ? _slots_31_io_out_uop_edge_inst : _GEN_684 ? _slots_30_io_out_uop_edge_inst : _slots_29_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_686 ? _slots_32_io_out_uop_pc_lob : _GEN_685 ? _slots_31_io_out_uop_pc_lob : _GEN_684 ? _slots_30_io_out_uop_pc_lob : _slots_29_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_686 ? _slots_32_io_out_uop_taken : _GEN_685 ? _slots_31_io_out_uop_taken : _GEN_684 ? _slots_30_io_out_uop_taken : _slots_29_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_686 ? _slots_32_io_out_uop_imm_packed : _GEN_685 ? _slots_31_io_out_uop_imm_packed : _GEN_684 ? _slots_30_io_out_uop_imm_packed : _slots_29_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_686 ? _slots_32_io_out_uop_rob_idx : _GEN_685 ? _slots_31_io_out_uop_rob_idx : _GEN_684 ? _slots_30_io_out_uop_rob_idx : _slots_29_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_686 ? _slots_32_io_out_uop_ldq_idx : _GEN_685 ? _slots_31_io_out_uop_ldq_idx : _GEN_684 ? _slots_30_io_out_uop_ldq_idx : _slots_29_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_686 ? _slots_32_io_out_uop_stq_idx : _GEN_685 ? _slots_31_io_out_uop_stq_idx : _GEN_684 ? _slots_30_io_out_uop_stq_idx : _slots_29_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_686 ? _slots_32_io_out_uop_pdst : _GEN_685 ? _slots_31_io_out_uop_pdst : _GEN_684 ? _slots_30_io_out_uop_pdst : _slots_29_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_686 ? _slots_32_io_out_uop_prs1 : _GEN_685 ? _slots_31_io_out_uop_prs1 : _GEN_684 ? _slots_30_io_out_uop_prs1 : _slots_29_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_686 ? _slots_32_io_out_uop_prs2 : _GEN_685 ? _slots_31_io_out_uop_prs2 : _GEN_684 ? _slots_30_io_out_uop_prs2 : _slots_29_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_686 ? _slots_32_io_out_uop_prs3 : _GEN_685 ? _slots_31_io_out_uop_prs3 : _GEN_684 ? _slots_30_io_out_uop_prs3 : _slots_29_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_686 ? _slots_32_io_out_uop_prs1_busy : _GEN_685 ? _slots_31_io_out_uop_prs1_busy : _GEN_684 ? _slots_30_io_out_uop_prs1_busy : _slots_29_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_686 ? _slots_32_io_out_uop_prs2_busy : _GEN_685 ? _slots_31_io_out_uop_prs2_busy : _GEN_684 ? _slots_30_io_out_uop_prs2_busy : _slots_29_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_686 ? _slots_32_io_out_uop_prs3_busy : _GEN_685 ? _slots_31_io_out_uop_prs3_busy : _GEN_684 ? _slots_30_io_out_uop_prs3_busy : _slots_29_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_686 ? _slots_32_io_out_uop_ppred_busy : _GEN_685 ? _slots_31_io_out_uop_ppred_busy : _GEN_684 ? _slots_30_io_out_uop_ppred_busy : _slots_29_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_686 ? _slots_32_io_out_uop_bypassable : _GEN_685 ? _slots_31_io_out_uop_bypassable : _GEN_684 ? _slots_30_io_out_uop_bypassable : _slots_29_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_686 ? _slots_32_io_out_uop_mem_cmd : _GEN_685 ? _slots_31_io_out_uop_mem_cmd : _GEN_684 ? _slots_30_io_out_uop_mem_cmd : _slots_29_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_686 ? _slots_32_io_out_uop_mem_size : _GEN_685 ? _slots_31_io_out_uop_mem_size : _GEN_684 ? _slots_30_io_out_uop_mem_size : _slots_29_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_686 ? _slots_32_io_out_uop_mem_signed : _GEN_685 ? _slots_31_io_out_uop_mem_signed : _GEN_684 ? _slots_30_io_out_uop_mem_signed : _slots_29_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_686 ? _slots_32_io_out_uop_is_fence : _GEN_685 ? _slots_31_io_out_uop_is_fence : _GEN_684 ? _slots_30_io_out_uop_is_fence : _slots_29_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_686 ? _slots_32_io_out_uop_is_amo : _GEN_685 ? _slots_31_io_out_uop_is_amo : _GEN_684 ? _slots_30_io_out_uop_is_amo : _slots_29_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_686 ? _slots_32_io_out_uop_uses_ldq : _GEN_685 ? _slots_31_io_out_uop_uses_ldq : _GEN_684 ? _slots_30_io_out_uop_uses_ldq : _slots_29_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_686 ? _slots_32_io_out_uop_uses_stq : _GEN_685 ? _slots_31_io_out_uop_uses_stq : _GEN_684 ? _slots_30_io_out_uop_uses_stq : _slots_29_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_686 ? _slots_32_io_out_uop_ldst_val : _GEN_685 ? _slots_31_io_out_uop_ldst_val : _GEN_684 ? _slots_30_io_out_uop_ldst_val : _slots_29_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_686 ? _slots_32_io_out_uop_dst_rtype : _GEN_685 ? _slots_31_io_out_uop_dst_rtype : _GEN_684 ? _slots_30_io_out_uop_dst_rtype : _slots_29_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_686 ? _slots_32_io_out_uop_lrs1_rtype : _GEN_685 ? _slots_31_io_out_uop_lrs1_rtype : _GEN_684 ? _slots_30_io_out_uop_lrs1_rtype : _slots_29_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_686 ? _slots_32_io_out_uop_lrs2_rtype : _GEN_685 ? _slots_31_io_out_uop_lrs2_rtype : _GEN_684 ? _slots_30_io_out_uop_lrs2_rtype : _slots_29_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_686 ? _slots_32_io_out_uop_fp_val : _GEN_685 ? _slots_31_io_out_uop_fp_val : _GEN_684 ? _slots_30_io_out_uop_fp_val : _slots_29_io_out_uop_fp_val),
    .io_valid                       (_slots_28_io_valid),
    .io_will_be_valid               (_slots_28_io_will_be_valid),
    .io_request                     (_slots_28_io_request),
    .io_out_uop_uopc                (_slots_28_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_28_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_28_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_28_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_28_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_28_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_28_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_28_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_28_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_28_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_28_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_28_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_28_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_28_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_28_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_28_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_28_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_28_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_28_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_28_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_28_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_28_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_28_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_28_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_28_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_28_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_28_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_28_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_28_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_28_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_28_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_28_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_28_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_28_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_28_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_28_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_28_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_28_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_28_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_28_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_28_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_28_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_28_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_28_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_28_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_28_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_28_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_28_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_28_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_28_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_28_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_28_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_28_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_28_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_28_io_uop_pc_lob),
    .io_uop_taken                   (_slots_28_io_uop_taken),
    .io_uop_imm_packed              (_slots_28_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_28_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_28_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_28_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_28_io_uop_pdst),
    .io_uop_prs1                    (_slots_28_io_uop_prs1),
    .io_uop_prs2                    (_slots_28_io_uop_prs2),
    .io_uop_bypassable              (_slots_28_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_28_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_28_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_28_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_28_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_28_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_28_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_28_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_28_io_uop_fp_val)
  );
  IssueSlot_32 slots_29 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_29_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_77),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_29_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_689 ? _slots_33_io_out_uop_uopc : _GEN_688 ? _slots_32_io_out_uop_uopc : _GEN_687 ? _slots_31_io_out_uop_uopc : _slots_30_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_689 ? _slots_33_io_out_uop_is_rvc : _GEN_688 ? _slots_32_io_out_uop_is_rvc : _GEN_687 ? _slots_31_io_out_uop_is_rvc : _slots_30_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_689 ? _slots_33_io_out_uop_fu_code : _GEN_688 ? _slots_32_io_out_uop_fu_code : _GEN_687 ? _slots_31_io_out_uop_fu_code : _slots_30_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_689 ? _slots_33_io_out_uop_iw_state : _GEN_688 ? _slots_32_io_out_uop_iw_state : _GEN_687 ? _slots_31_io_out_uop_iw_state : _slots_30_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_689 ? _slots_33_io_out_uop_iw_p1_poisoned : _GEN_688 ? _slots_32_io_out_uop_iw_p1_poisoned : _GEN_687 ? _slots_31_io_out_uop_iw_p1_poisoned : _slots_30_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_689 ? _slots_33_io_out_uop_iw_p2_poisoned : _GEN_688 ? _slots_32_io_out_uop_iw_p2_poisoned : _GEN_687 ? _slots_31_io_out_uop_iw_p2_poisoned : _slots_30_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_689 ? _slots_33_io_out_uop_is_br : _GEN_688 ? _slots_32_io_out_uop_is_br : _GEN_687 ? _slots_31_io_out_uop_is_br : _slots_30_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_689 ? _slots_33_io_out_uop_is_jalr : _GEN_688 ? _slots_32_io_out_uop_is_jalr : _GEN_687 ? _slots_31_io_out_uop_is_jalr : _slots_30_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_689 ? _slots_33_io_out_uop_is_jal : _GEN_688 ? _slots_32_io_out_uop_is_jal : _GEN_687 ? _slots_31_io_out_uop_is_jal : _slots_30_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_689 ? _slots_33_io_out_uop_is_sfb : _GEN_688 ? _slots_32_io_out_uop_is_sfb : _GEN_687 ? _slots_31_io_out_uop_is_sfb : _slots_30_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_689 ? _slots_33_io_out_uop_br_mask : _GEN_688 ? _slots_32_io_out_uop_br_mask : _GEN_687 ? _slots_31_io_out_uop_br_mask : _slots_30_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_689 ? _slots_33_io_out_uop_br_tag : _GEN_688 ? _slots_32_io_out_uop_br_tag : _GEN_687 ? _slots_31_io_out_uop_br_tag : _slots_30_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_689 ? _slots_33_io_out_uop_ftq_idx : _GEN_688 ? _slots_32_io_out_uop_ftq_idx : _GEN_687 ? _slots_31_io_out_uop_ftq_idx : _slots_30_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_689 ? _slots_33_io_out_uop_edge_inst : _GEN_688 ? _slots_32_io_out_uop_edge_inst : _GEN_687 ? _slots_31_io_out_uop_edge_inst : _slots_30_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_689 ? _slots_33_io_out_uop_pc_lob : _GEN_688 ? _slots_32_io_out_uop_pc_lob : _GEN_687 ? _slots_31_io_out_uop_pc_lob : _slots_30_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_689 ? _slots_33_io_out_uop_taken : _GEN_688 ? _slots_32_io_out_uop_taken : _GEN_687 ? _slots_31_io_out_uop_taken : _slots_30_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_689 ? _slots_33_io_out_uop_imm_packed : _GEN_688 ? _slots_32_io_out_uop_imm_packed : _GEN_687 ? _slots_31_io_out_uop_imm_packed : _slots_30_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_689 ? _slots_33_io_out_uop_rob_idx : _GEN_688 ? _slots_32_io_out_uop_rob_idx : _GEN_687 ? _slots_31_io_out_uop_rob_idx : _slots_30_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_689 ? _slots_33_io_out_uop_ldq_idx : _GEN_688 ? _slots_32_io_out_uop_ldq_idx : _GEN_687 ? _slots_31_io_out_uop_ldq_idx : _slots_30_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_689 ? _slots_33_io_out_uop_stq_idx : _GEN_688 ? _slots_32_io_out_uop_stq_idx : _GEN_687 ? _slots_31_io_out_uop_stq_idx : _slots_30_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_689 ? _slots_33_io_out_uop_pdst : _GEN_688 ? _slots_32_io_out_uop_pdst : _GEN_687 ? _slots_31_io_out_uop_pdst : _slots_30_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_689 ? _slots_33_io_out_uop_prs1 : _GEN_688 ? _slots_32_io_out_uop_prs1 : _GEN_687 ? _slots_31_io_out_uop_prs1 : _slots_30_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_689 ? _slots_33_io_out_uop_prs2 : _GEN_688 ? _slots_32_io_out_uop_prs2 : _GEN_687 ? _slots_31_io_out_uop_prs2 : _slots_30_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_689 ? _slots_33_io_out_uop_prs3 : _GEN_688 ? _slots_32_io_out_uop_prs3 : _GEN_687 ? _slots_31_io_out_uop_prs3 : _slots_30_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_689 ? _slots_33_io_out_uop_prs1_busy : _GEN_688 ? _slots_32_io_out_uop_prs1_busy : _GEN_687 ? _slots_31_io_out_uop_prs1_busy : _slots_30_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_689 ? _slots_33_io_out_uop_prs2_busy : _GEN_688 ? _slots_32_io_out_uop_prs2_busy : _GEN_687 ? _slots_31_io_out_uop_prs2_busy : _slots_30_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_689 ? _slots_33_io_out_uop_prs3_busy : _GEN_688 ? _slots_32_io_out_uop_prs3_busy : _GEN_687 ? _slots_31_io_out_uop_prs3_busy : _slots_30_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_689 ? _slots_33_io_out_uop_ppred_busy : _GEN_688 ? _slots_32_io_out_uop_ppred_busy : _GEN_687 ? _slots_31_io_out_uop_ppred_busy : _slots_30_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_689 ? _slots_33_io_out_uop_bypassable : _GEN_688 ? _slots_32_io_out_uop_bypassable : _GEN_687 ? _slots_31_io_out_uop_bypassable : _slots_30_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_689 ? _slots_33_io_out_uop_mem_cmd : _GEN_688 ? _slots_32_io_out_uop_mem_cmd : _GEN_687 ? _slots_31_io_out_uop_mem_cmd : _slots_30_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_689 ? _slots_33_io_out_uop_mem_size : _GEN_688 ? _slots_32_io_out_uop_mem_size : _GEN_687 ? _slots_31_io_out_uop_mem_size : _slots_30_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_689 ? _slots_33_io_out_uop_mem_signed : _GEN_688 ? _slots_32_io_out_uop_mem_signed : _GEN_687 ? _slots_31_io_out_uop_mem_signed : _slots_30_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_689 ? _slots_33_io_out_uop_is_fence : _GEN_688 ? _slots_32_io_out_uop_is_fence : _GEN_687 ? _slots_31_io_out_uop_is_fence : _slots_30_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_689 ? _slots_33_io_out_uop_is_amo : _GEN_688 ? _slots_32_io_out_uop_is_amo : _GEN_687 ? _slots_31_io_out_uop_is_amo : _slots_30_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_689 ? _slots_33_io_out_uop_uses_ldq : _GEN_688 ? _slots_32_io_out_uop_uses_ldq : _GEN_687 ? _slots_31_io_out_uop_uses_ldq : _slots_30_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_689 ? _slots_33_io_out_uop_uses_stq : _GEN_688 ? _slots_32_io_out_uop_uses_stq : _GEN_687 ? _slots_31_io_out_uop_uses_stq : _slots_30_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_689 ? _slots_33_io_out_uop_ldst_val : _GEN_688 ? _slots_32_io_out_uop_ldst_val : _GEN_687 ? _slots_31_io_out_uop_ldst_val : _slots_30_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_689 ? _slots_33_io_out_uop_dst_rtype : _GEN_688 ? _slots_32_io_out_uop_dst_rtype : _GEN_687 ? _slots_31_io_out_uop_dst_rtype : _slots_30_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_689 ? _slots_33_io_out_uop_lrs1_rtype : _GEN_688 ? _slots_32_io_out_uop_lrs1_rtype : _GEN_687 ? _slots_31_io_out_uop_lrs1_rtype : _slots_30_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_689 ? _slots_33_io_out_uop_lrs2_rtype : _GEN_688 ? _slots_32_io_out_uop_lrs2_rtype : _GEN_687 ? _slots_31_io_out_uop_lrs2_rtype : _slots_30_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_689 ? _slots_33_io_out_uop_fp_val : _GEN_688 ? _slots_32_io_out_uop_fp_val : _GEN_687 ? _slots_31_io_out_uop_fp_val : _slots_30_io_out_uop_fp_val),
    .io_valid                       (_slots_29_io_valid),
    .io_will_be_valid               (_slots_29_io_will_be_valid),
    .io_request                     (_slots_29_io_request),
    .io_out_uop_uopc                (_slots_29_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_29_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_29_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_29_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_29_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_29_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_29_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_29_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_29_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_29_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_29_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_29_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_29_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_29_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_29_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_29_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_29_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_29_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_29_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_29_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_29_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_29_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_29_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_29_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_29_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_29_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_29_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_29_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_29_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_29_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_29_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_29_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_29_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_29_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_29_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_29_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_29_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_29_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_29_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_29_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_29_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_29_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_29_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_29_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_29_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_29_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_29_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_29_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_29_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_29_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_29_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_29_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_29_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_29_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_29_io_uop_pc_lob),
    .io_uop_taken                   (_slots_29_io_uop_taken),
    .io_uop_imm_packed              (_slots_29_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_29_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_29_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_29_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_29_io_uop_pdst),
    .io_uop_prs1                    (_slots_29_io_uop_prs1),
    .io_uop_prs2                    (_slots_29_io_uop_prs2),
    .io_uop_bypassable              (_slots_29_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_29_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_29_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_29_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_29_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_29_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_29_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_29_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_29_io_uop_fp_val)
  );
  IssueSlot_32 slots_30 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_30_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_79),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_30_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_692 ? _slots_34_io_out_uop_uopc : _GEN_691 ? _slots_33_io_out_uop_uopc : _GEN_690 ? _slots_32_io_out_uop_uopc : _slots_31_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_692 ? _slots_34_io_out_uop_is_rvc : _GEN_691 ? _slots_33_io_out_uop_is_rvc : _GEN_690 ? _slots_32_io_out_uop_is_rvc : _slots_31_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_692 ? _slots_34_io_out_uop_fu_code : _GEN_691 ? _slots_33_io_out_uop_fu_code : _GEN_690 ? _slots_32_io_out_uop_fu_code : _slots_31_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_692 ? _slots_34_io_out_uop_iw_state : _GEN_691 ? _slots_33_io_out_uop_iw_state : _GEN_690 ? _slots_32_io_out_uop_iw_state : _slots_31_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_692 ? _slots_34_io_out_uop_iw_p1_poisoned : _GEN_691 ? _slots_33_io_out_uop_iw_p1_poisoned : _GEN_690 ? _slots_32_io_out_uop_iw_p1_poisoned : _slots_31_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_692 ? _slots_34_io_out_uop_iw_p2_poisoned : _GEN_691 ? _slots_33_io_out_uop_iw_p2_poisoned : _GEN_690 ? _slots_32_io_out_uop_iw_p2_poisoned : _slots_31_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_692 ? _slots_34_io_out_uop_is_br : _GEN_691 ? _slots_33_io_out_uop_is_br : _GEN_690 ? _slots_32_io_out_uop_is_br : _slots_31_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_692 ? _slots_34_io_out_uop_is_jalr : _GEN_691 ? _slots_33_io_out_uop_is_jalr : _GEN_690 ? _slots_32_io_out_uop_is_jalr : _slots_31_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_692 ? _slots_34_io_out_uop_is_jal : _GEN_691 ? _slots_33_io_out_uop_is_jal : _GEN_690 ? _slots_32_io_out_uop_is_jal : _slots_31_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_692 ? _slots_34_io_out_uop_is_sfb : _GEN_691 ? _slots_33_io_out_uop_is_sfb : _GEN_690 ? _slots_32_io_out_uop_is_sfb : _slots_31_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_692 ? _slots_34_io_out_uop_br_mask : _GEN_691 ? _slots_33_io_out_uop_br_mask : _GEN_690 ? _slots_32_io_out_uop_br_mask : _slots_31_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_692 ? _slots_34_io_out_uop_br_tag : _GEN_691 ? _slots_33_io_out_uop_br_tag : _GEN_690 ? _slots_32_io_out_uop_br_tag : _slots_31_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_692 ? _slots_34_io_out_uop_ftq_idx : _GEN_691 ? _slots_33_io_out_uop_ftq_idx : _GEN_690 ? _slots_32_io_out_uop_ftq_idx : _slots_31_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_692 ? _slots_34_io_out_uop_edge_inst : _GEN_691 ? _slots_33_io_out_uop_edge_inst : _GEN_690 ? _slots_32_io_out_uop_edge_inst : _slots_31_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_692 ? _slots_34_io_out_uop_pc_lob : _GEN_691 ? _slots_33_io_out_uop_pc_lob : _GEN_690 ? _slots_32_io_out_uop_pc_lob : _slots_31_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_692 ? _slots_34_io_out_uop_taken : _GEN_691 ? _slots_33_io_out_uop_taken : _GEN_690 ? _slots_32_io_out_uop_taken : _slots_31_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_692 ? _slots_34_io_out_uop_imm_packed : _GEN_691 ? _slots_33_io_out_uop_imm_packed : _GEN_690 ? _slots_32_io_out_uop_imm_packed : _slots_31_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_692 ? _slots_34_io_out_uop_rob_idx : _GEN_691 ? _slots_33_io_out_uop_rob_idx : _GEN_690 ? _slots_32_io_out_uop_rob_idx : _slots_31_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_692 ? _slots_34_io_out_uop_ldq_idx : _GEN_691 ? _slots_33_io_out_uop_ldq_idx : _GEN_690 ? _slots_32_io_out_uop_ldq_idx : _slots_31_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_692 ? _slots_34_io_out_uop_stq_idx : _GEN_691 ? _slots_33_io_out_uop_stq_idx : _GEN_690 ? _slots_32_io_out_uop_stq_idx : _slots_31_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_692 ? _slots_34_io_out_uop_pdst : _GEN_691 ? _slots_33_io_out_uop_pdst : _GEN_690 ? _slots_32_io_out_uop_pdst : _slots_31_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_692 ? _slots_34_io_out_uop_prs1 : _GEN_691 ? _slots_33_io_out_uop_prs1 : _GEN_690 ? _slots_32_io_out_uop_prs1 : _slots_31_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_692 ? _slots_34_io_out_uop_prs2 : _GEN_691 ? _slots_33_io_out_uop_prs2 : _GEN_690 ? _slots_32_io_out_uop_prs2 : _slots_31_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_692 ? _slots_34_io_out_uop_prs3 : _GEN_691 ? _slots_33_io_out_uop_prs3 : _GEN_690 ? _slots_32_io_out_uop_prs3 : _slots_31_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_692 ? _slots_34_io_out_uop_prs1_busy : _GEN_691 ? _slots_33_io_out_uop_prs1_busy : _GEN_690 ? _slots_32_io_out_uop_prs1_busy : _slots_31_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_692 ? _slots_34_io_out_uop_prs2_busy : _GEN_691 ? _slots_33_io_out_uop_prs2_busy : _GEN_690 ? _slots_32_io_out_uop_prs2_busy : _slots_31_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_692 ? _slots_34_io_out_uop_prs3_busy : _GEN_691 ? _slots_33_io_out_uop_prs3_busy : _GEN_690 ? _slots_32_io_out_uop_prs3_busy : _slots_31_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_692 ? _slots_34_io_out_uop_ppred_busy : _GEN_691 ? _slots_33_io_out_uop_ppred_busy : _GEN_690 ? _slots_32_io_out_uop_ppred_busy : _slots_31_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_692 ? _slots_34_io_out_uop_bypassable : _GEN_691 ? _slots_33_io_out_uop_bypassable : _GEN_690 ? _slots_32_io_out_uop_bypassable : _slots_31_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_692 ? _slots_34_io_out_uop_mem_cmd : _GEN_691 ? _slots_33_io_out_uop_mem_cmd : _GEN_690 ? _slots_32_io_out_uop_mem_cmd : _slots_31_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_692 ? _slots_34_io_out_uop_mem_size : _GEN_691 ? _slots_33_io_out_uop_mem_size : _GEN_690 ? _slots_32_io_out_uop_mem_size : _slots_31_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_692 ? _slots_34_io_out_uop_mem_signed : _GEN_691 ? _slots_33_io_out_uop_mem_signed : _GEN_690 ? _slots_32_io_out_uop_mem_signed : _slots_31_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_692 ? _slots_34_io_out_uop_is_fence : _GEN_691 ? _slots_33_io_out_uop_is_fence : _GEN_690 ? _slots_32_io_out_uop_is_fence : _slots_31_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_692 ? _slots_34_io_out_uop_is_amo : _GEN_691 ? _slots_33_io_out_uop_is_amo : _GEN_690 ? _slots_32_io_out_uop_is_amo : _slots_31_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_692 ? _slots_34_io_out_uop_uses_ldq : _GEN_691 ? _slots_33_io_out_uop_uses_ldq : _GEN_690 ? _slots_32_io_out_uop_uses_ldq : _slots_31_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_692 ? _slots_34_io_out_uop_uses_stq : _GEN_691 ? _slots_33_io_out_uop_uses_stq : _GEN_690 ? _slots_32_io_out_uop_uses_stq : _slots_31_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_692 ? _slots_34_io_out_uop_ldst_val : _GEN_691 ? _slots_33_io_out_uop_ldst_val : _GEN_690 ? _slots_32_io_out_uop_ldst_val : _slots_31_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_692 ? _slots_34_io_out_uop_dst_rtype : _GEN_691 ? _slots_33_io_out_uop_dst_rtype : _GEN_690 ? _slots_32_io_out_uop_dst_rtype : _slots_31_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_692 ? _slots_34_io_out_uop_lrs1_rtype : _GEN_691 ? _slots_33_io_out_uop_lrs1_rtype : _GEN_690 ? _slots_32_io_out_uop_lrs1_rtype : _slots_31_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_692 ? _slots_34_io_out_uop_lrs2_rtype : _GEN_691 ? _slots_33_io_out_uop_lrs2_rtype : _GEN_690 ? _slots_32_io_out_uop_lrs2_rtype : _slots_31_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_692 ? _slots_34_io_out_uop_fp_val : _GEN_691 ? _slots_33_io_out_uop_fp_val : _GEN_690 ? _slots_32_io_out_uop_fp_val : _slots_31_io_out_uop_fp_val),
    .io_valid                       (_slots_30_io_valid),
    .io_will_be_valid               (_slots_30_io_will_be_valid),
    .io_request                     (_slots_30_io_request),
    .io_out_uop_uopc                (_slots_30_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_30_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_30_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_30_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_30_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_30_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_30_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_30_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_30_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_30_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_30_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_30_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_30_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_30_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_30_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_30_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_30_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_30_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_30_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_30_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_30_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_30_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_30_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_30_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_30_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_30_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_30_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_30_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_30_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_30_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_30_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_30_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_30_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_30_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_30_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_30_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_30_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_30_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_30_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_30_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_30_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_30_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_30_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_30_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_30_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_30_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_30_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_30_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_30_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_30_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_30_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_30_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_30_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_30_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_30_io_uop_pc_lob),
    .io_uop_taken                   (_slots_30_io_uop_taken),
    .io_uop_imm_packed              (_slots_30_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_30_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_30_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_30_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_30_io_uop_pdst),
    .io_uop_prs1                    (_slots_30_io_uop_prs1),
    .io_uop_prs2                    (_slots_30_io_uop_prs2),
    .io_uop_bypassable              (_slots_30_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_30_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_30_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_30_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_30_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_30_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_30_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_30_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_30_io_uop_fp_val)
  );
  IssueSlot_32 slots_31 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_31_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_81),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_31_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_695 ? _slots_35_io_out_uop_uopc : _GEN_694 ? _slots_34_io_out_uop_uopc : _GEN_693 ? _slots_33_io_out_uop_uopc : _slots_32_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_695 ? _slots_35_io_out_uop_is_rvc : _GEN_694 ? _slots_34_io_out_uop_is_rvc : _GEN_693 ? _slots_33_io_out_uop_is_rvc : _slots_32_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_695 ? _slots_35_io_out_uop_fu_code : _GEN_694 ? _slots_34_io_out_uop_fu_code : _GEN_693 ? _slots_33_io_out_uop_fu_code : _slots_32_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_695 ? _slots_35_io_out_uop_iw_state : _GEN_694 ? _slots_34_io_out_uop_iw_state : _GEN_693 ? _slots_33_io_out_uop_iw_state : _slots_32_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_695 ? _slots_35_io_out_uop_iw_p1_poisoned : _GEN_694 ? _slots_34_io_out_uop_iw_p1_poisoned : _GEN_693 ? _slots_33_io_out_uop_iw_p1_poisoned : _slots_32_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_695 ? _slots_35_io_out_uop_iw_p2_poisoned : _GEN_694 ? _slots_34_io_out_uop_iw_p2_poisoned : _GEN_693 ? _slots_33_io_out_uop_iw_p2_poisoned : _slots_32_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_695 ? _slots_35_io_out_uop_is_br : _GEN_694 ? _slots_34_io_out_uop_is_br : _GEN_693 ? _slots_33_io_out_uop_is_br : _slots_32_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_695 ? _slots_35_io_out_uop_is_jalr : _GEN_694 ? _slots_34_io_out_uop_is_jalr : _GEN_693 ? _slots_33_io_out_uop_is_jalr : _slots_32_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_695 ? _slots_35_io_out_uop_is_jal : _GEN_694 ? _slots_34_io_out_uop_is_jal : _GEN_693 ? _slots_33_io_out_uop_is_jal : _slots_32_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_695 ? _slots_35_io_out_uop_is_sfb : _GEN_694 ? _slots_34_io_out_uop_is_sfb : _GEN_693 ? _slots_33_io_out_uop_is_sfb : _slots_32_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_695 ? _slots_35_io_out_uop_br_mask : _GEN_694 ? _slots_34_io_out_uop_br_mask : _GEN_693 ? _slots_33_io_out_uop_br_mask : _slots_32_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_695 ? _slots_35_io_out_uop_br_tag : _GEN_694 ? _slots_34_io_out_uop_br_tag : _GEN_693 ? _slots_33_io_out_uop_br_tag : _slots_32_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_695 ? _slots_35_io_out_uop_ftq_idx : _GEN_694 ? _slots_34_io_out_uop_ftq_idx : _GEN_693 ? _slots_33_io_out_uop_ftq_idx : _slots_32_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_695 ? _slots_35_io_out_uop_edge_inst : _GEN_694 ? _slots_34_io_out_uop_edge_inst : _GEN_693 ? _slots_33_io_out_uop_edge_inst : _slots_32_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_695 ? _slots_35_io_out_uop_pc_lob : _GEN_694 ? _slots_34_io_out_uop_pc_lob : _GEN_693 ? _slots_33_io_out_uop_pc_lob : _slots_32_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_695 ? _slots_35_io_out_uop_taken : _GEN_694 ? _slots_34_io_out_uop_taken : _GEN_693 ? _slots_33_io_out_uop_taken : _slots_32_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_695 ? _slots_35_io_out_uop_imm_packed : _GEN_694 ? _slots_34_io_out_uop_imm_packed : _GEN_693 ? _slots_33_io_out_uop_imm_packed : _slots_32_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_695 ? _slots_35_io_out_uop_rob_idx : _GEN_694 ? _slots_34_io_out_uop_rob_idx : _GEN_693 ? _slots_33_io_out_uop_rob_idx : _slots_32_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_695 ? _slots_35_io_out_uop_ldq_idx : _GEN_694 ? _slots_34_io_out_uop_ldq_idx : _GEN_693 ? _slots_33_io_out_uop_ldq_idx : _slots_32_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_695 ? _slots_35_io_out_uop_stq_idx : _GEN_694 ? _slots_34_io_out_uop_stq_idx : _GEN_693 ? _slots_33_io_out_uop_stq_idx : _slots_32_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_695 ? _slots_35_io_out_uop_pdst : _GEN_694 ? _slots_34_io_out_uop_pdst : _GEN_693 ? _slots_33_io_out_uop_pdst : _slots_32_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_695 ? _slots_35_io_out_uop_prs1 : _GEN_694 ? _slots_34_io_out_uop_prs1 : _GEN_693 ? _slots_33_io_out_uop_prs1 : _slots_32_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_695 ? _slots_35_io_out_uop_prs2 : _GEN_694 ? _slots_34_io_out_uop_prs2 : _GEN_693 ? _slots_33_io_out_uop_prs2 : _slots_32_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_695 ? _slots_35_io_out_uop_prs3 : _GEN_694 ? _slots_34_io_out_uop_prs3 : _GEN_693 ? _slots_33_io_out_uop_prs3 : _slots_32_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_695 ? _slots_35_io_out_uop_prs1_busy : _GEN_694 ? _slots_34_io_out_uop_prs1_busy : _GEN_693 ? _slots_33_io_out_uop_prs1_busy : _slots_32_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_695 ? _slots_35_io_out_uop_prs2_busy : _GEN_694 ? _slots_34_io_out_uop_prs2_busy : _GEN_693 ? _slots_33_io_out_uop_prs2_busy : _slots_32_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_695 ? _slots_35_io_out_uop_prs3_busy : _GEN_694 ? _slots_34_io_out_uop_prs3_busy : _GEN_693 ? _slots_33_io_out_uop_prs3_busy : _slots_32_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_695 ? _slots_35_io_out_uop_ppred_busy : _GEN_694 ? _slots_34_io_out_uop_ppred_busy : _GEN_693 ? _slots_33_io_out_uop_ppred_busy : _slots_32_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_695 ? _slots_35_io_out_uop_bypassable : _GEN_694 ? _slots_34_io_out_uop_bypassable : _GEN_693 ? _slots_33_io_out_uop_bypassable : _slots_32_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_695 ? _slots_35_io_out_uop_mem_cmd : _GEN_694 ? _slots_34_io_out_uop_mem_cmd : _GEN_693 ? _slots_33_io_out_uop_mem_cmd : _slots_32_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_695 ? _slots_35_io_out_uop_mem_size : _GEN_694 ? _slots_34_io_out_uop_mem_size : _GEN_693 ? _slots_33_io_out_uop_mem_size : _slots_32_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_695 ? _slots_35_io_out_uop_mem_signed : _GEN_694 ? _slots_34_io_out_uop_mem_signed : _GEN_693 ? _slots_33_io_out_uop_mem_signed : _slots_32_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_695 ? _slots_35_io_out_uop_is_fence : _GEN_694 ? _slots_34_io_out_uop_is_fence : _GEN_693 ? _slots_33_io_out_uop_is_fence : _slots_32_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_695 ? _slots_35_io_out_uop_is_amo : _GEN_694 ? _slots_34_io_out_uop_is_amo : _GEN_693 ? _slots_33_io_out_uop_is_amo : _slots_32_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_695 ? _slots_35_io_out_uop_uses_ldq : _GEN_694 ? _slots_34_io_out_uop_uses_ldq : _GEN_693 ? _slots_33_io_out_uop_uses_ldq : _slots_32_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_695 ? _slots_35_io_out_uop_uses_stq : _GEN_694 ? _slots_34_io_out_uop_uses_stq : _GEN_693 ? _slots_33_io_out_uop_uses_stq : _slots_32_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_695 ? _slots_35_io_out_uop_ldst_val : _GEN_694 ? _slots_34_io_out_uop_ldst_val : _GEN_693 ? _slots_33_io_out_uop_ldst_val : _slots_32_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_695 ? _slots_35_io_out_uop_dst_rtype : _GEN_694 ? _slots_34_io_out_uop_dst_rtype : _GEN_693 ? _slots_33_io_out_uop_dst_rtype : _slots_32_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_695 ? _slots_35_io_out_uop_lrs1_rtype : _GEN_694 ? _slots_34_io_out_uop_lrs1_rtype : _GEN_693 ? _slots_33_io_out_uop_lrs1_rtype : _slots_32_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_695 ? _slots_35_io_out_uop_lrs2_rtype : _GEN_694 ? _slots_34_io_out_uop_lrs2_rtype : _GEN_693 ? _slots_33_io_out_uop_lrs2_rtype : _slots_32_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_695 ? _slots_35_io_out_uop_fp_val : _GEN_694 ? _slots_34_io_out_uop_fp_val : _GEN_693 ? _slots_33_io_out_uop_fp_val : _slots_32_io_out_uop_fp_val),
    .io_valid                       (_slots_31_io_valid),
    .io_will_be_valid               (_slots_31_io_will_be_valid),
    .io_request                     (_slots_31_io_request),
    .io_out_uop_uopc                (_slots_31_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_31_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_31_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_31_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_31_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_31_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_31_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_31_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_31_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_31_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_31_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_31_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_31_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_31_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_31_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_31_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_31_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_31_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_31_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_31_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_31_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_31_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_31_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_31_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_31_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_31_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_31_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_31_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_31_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_31_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_31_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_31_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_31_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_31_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_31_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_31_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_31_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_31_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_31_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_31_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_31_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_31_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_31_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_31_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_31_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_31_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_31_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_31_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_31_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_31_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_31_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_31_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_31_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_31_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_31_io_uop_pc_lob),
    .io_uop_taken                   (_slots_31_io_uop_taken),
    .io_uop_imm_packed              (_slots_31_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_31_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_31_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_31_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_31_io_uop_pdst),
    .io_uop_prs1                    (_slots_31_io_uop_prs1),
    .io_uop_prs2                    (_slots_31_io_uop_prs2),
    .io_uop_bypassable              (_slots_31_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_31_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_31_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_31_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_31_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_31_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_31_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_31_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_31_io_uop_fp_val)
  );
  IssueSlot_32 slots_32 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_32_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_83),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_32_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_698 ? _slots_36_io_out_uop_uopc : _GEN_697 ? _slots_35_io_out_uop_uopc : _GEN_696 ? _slots_34_io_out_uop_uopc : _slots_33_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_698 ? _slots_36_io_out_uop_is_rvc : _GEN_697 ? _slots_35_io_out_uop_is_rvc : _GEN_696 ? _slots_34_io_out_uop_is_rvc : _slots_33_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_698 ? _slots_36_io_out_uop_fu_code : _GEN_697 ? _slots_35_io_out_uop_fu_code : _GEN_696 ? _slots_34_io_out_uop_fu_code : _slots_33_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_698 ? _slots_36_io_out_uop_iw_state : _GEN_697 ? _slots_35_io_out_uop_iw_state : _GEN_696 ? _slots_34_io_out_uop_iw_state : _slots_33_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_698 ? _slots_36_io_out_uop_iw_p1_poisoned : _GEN_697 ? _slots_35_io_out_uop_iw_p1_poisoned : _GEN_696 ? _slots_34_io_out_uop_iw_p1_poisoned : _slots_33_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_698 ? _slots_36_io_out_uop_iw_p2_poisoned : _GEN_697 ? _slots_35_io_out_uop_iw_p2_poisoned : _GEN_696 ? _slots_34_io_out_uop_iw_p2_poisoned : _slots_33_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_698 ? _slots_36_io_out_uop_is_br : _GEN_697 ? _slots_35_io_out_uop_is_br : _GEN_696 ? _slots_34_io_out_uop_is_br : _slots_33_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_698 ? _slots_36_io_out_uop_is_jalr : _GEN_697 ? _slots_35_io_out_uop_is_jalr : _GEN_696 ? _slots_34_io_out_uop_is_jalr : _slots_33_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_698 ? _slots_36_io_out_uop_is_jal : _GEN_697 ? _slots_35_io_out_uop_is_jal : _GEN_696 ? _slots_34_io_out_uop_is_jal : _slots_33_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_698 ? _slots_36_io_out_uop_is_sfb : _GEN_697 ? _slots_35_io_out_uop_is_sfb : _GEN_696 ? _slots_34_io_out_uop_is_sfb : _slots_33_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_698 ? _slots_36_io_out_uop_br_mask : _GEN_697 ? _slots_35_io_out_uop_br_mask : _GEN_696 ? _slots_34_io_out_uop_br_mask : _slots_33_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_698 ? _slots_36_io_out_uop_br_tag : _GEN_697 ? _slots_35_io_out_uop_br_tag : _GEN_696 ? _slots_34_io_out_uop_br_tag : _slots_33_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_698 ? _slots_36_io_out_uop_ftq_idx : _GEN_697 ? _slots_35_io_out_uop_ftq_idx : _GEN_696 ? _slots_34_io_out_uop_ftq_idx : _slots_33_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_698 ? _slots_36_io_out_uop_edge_inst : _GEN_697 ? _slots_35_io_out_uop_edge_inst : _GEN_696 ? _slots_34_io_out_uop_edge_inst : _slots_33_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_698 ? _slots_36_io_out_uop_pc_lob : _GEN_697 ? _slots_35_io_out_uop_pc_lob : _GEN_696 ? _slots_34_io_out_uop_pc_lob : _slots_33_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_698 ? _slots_36_io_out_uop_taken : _GEN_697 ? _slots_35_io_out_uop_taken : _GEN_696 ? _slots_34_io_out_uop_taken : _slots_33_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_698 ? _slots_36_io_out_uop_imm_packed : _GEN_697 ? _slots_35_io_out_uop_imm_packed : _GEN_696 ? _slots_34_io_out_uop_imm_packed : _slots_33_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_698 ? _slots_36_io_out_uop_rob_idx : _GEN_697 ? _slots_35_io_out_uop_rob_idx : _GEN_696 ? _slots_34_io_out_uop_rob_idx : _slots_33_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_698 ? _slots_36_io_out_uop_ldq_idx : _GEN_697 ? _slots_35_io_out_uop_ldq_idx : _GEN_696 ? _slots_34_io_out_uop_ldq_idx : _slots_33_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_698 ? _slots_36_io_out_uop_stq_idx : _GEN_697 ? _slots_35_io_out_uop_stq_idx : _GEN_696 ? _slots_34_io_out_uop_stq_idx : _slots_33_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_698 ? _slots_36_io_out_uop_pdst : _GEN_697 ? _slots_35_io_out_uop_pdst : _GEN_696 ? _slots_34_io_out_uop_pdst : _slots_33_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_698 ? _slots_36_io_out_uop_prs1 : _GEN_697 ? _slots_35_io_out_uop_prs1 : _GEN_696 ? _slots_34_io_out_uop_prs1 : _slots_33_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_698 ? _slots_36_io_out_uop_prs2 : _GEN_697 ? _slots_35_io_out_uop_prs2 : _GEN_696 ? _slots_34_io_out_uop_prs2 : _slots_33_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_698 ? _slots_36_io_out_uop_prs3 : _GEN_697 ? _slots_35_io_out_uop_prs3 : _GEN_696 ? _slots_34_io_out_uop_prs3 : _slots_33_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_698 ? _slots_36_io_out_uop_prs1_busy : _GEN_697 ? _slots_35_io_out_uop_prs1_busy : _GEN_696 ? _slots_34_io_out_uop_prs1_busy : _slots_33_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_698 ? _slots_36_io_out_uop_prs2_busy : _GEN_697 ? _slots_35_io_out_uop_prs2_busy : _GEN_696 ? _slots_34_io_out_uop_prs2_busy : _slots_33_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_698 ? _slots_36_io_out_uop_prs3_busy : _GEN_697 ? _slots_35_io_out_uop_prs3_busy : _GEN_696 ? _slots_34_io_out_uop_prs3_busy : _slots_33_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_698 ? _slots_36_io_out_uop_ppred_busy : _GEN_697 ? _slots_35_io_out_uop_ppred_busy : _GEN_696 ? _slots_34_io_out_uop_ppred_busy : _slots_33_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_698 ? _slots_36_io_out_uop_bypassable : _GEN_697 ? _slots_35_io_out_uop_bypassable : _GEN_696 ? _slots_34_io_out_uop_bypassable : _slots_33_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_698 ? _slots_36_io_out_uop_mem_cmd : _GEN_697 ? _slots_35_io_out_uop_mem_cmd : _GEN_696 ? _slots_34_io_out_uop_mem_cmd : _slots_33_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_698 ? _slots_36_io_out_uop_mem_size : _GEN_697 ? _slots_35_io_out_uop_mem_size : _GEN_696 ? _slots_34_io_out_uop_mem_size : _slots_33_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_698 ? _slots_36_io_out_uop_mem_signed : _GEN_697 ? _slots_35_io_out_uop_mem_signed : _GEN_696 ? _slots_34_io_out_uop_mem_signed : _slots_33_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_698 ? _slots_36_io_out_uop_is_fence : _GEN_697 ? _slots_35_io_out_uop_is_fence : _GEN_696 ? _slots_34_io_out_uop_is_fence : _slots_33_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_698 ? _slots_36_io_out_uop_is_amo : _GEN_697 ? _slots_35_io_out_uop_is_amo : _GEN_696 ? _slots_34_io_out_uop_is_amo : _slots_33_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_698 ? _slots_36_io_out_uop_uses_ldq : _GEN_697 ? _slots_35_io_out_uop_uses_ldq : _GEN_696 ? _slots_34_io_out_uop_uses_ldq : _slots_33_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_698 ? _slots_36_io_out_uop_uses_stq : _GEN_697 ? _slots_35_io_out_uop_uses_stq : _GEN_696 ? _slots_34_io_out_uop_uses_stq : _slots_33_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_698 ? _slots_36_io_out_uop_ldst_val : _GEN_697 ? _slots_35_io_out_uop_ldst_val : _GEN_696 ? _slots_34_io_out_uop_ldst_val : _slots_33_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_698 ? _slots_36_io_out_uop_dst_rtype : _GEN_697 ? _slots_35_io_out_uop_dst_rtype : _GEN_696 ? _slots_34_io_out_uop_dst_rtype : _slots_33_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_698 ? _slots_36_io_out_uop_lrs1_rtype : _GEN_697 ? _slots_35_io_out_uop_lrs1_rtype : _GEN_696 ? _slots_34_io_out_uop_lrs1_rtype : _slots_33_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_698 ? _slots_36_io_out_uop_lrs2_rtype : _GEN_697 ? _slots_35_io_out_uop_lrs2_rtype : _GEN_696 ? _slots_34_io_out_uop_lrs2_rtype : _slots_33_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_698 ? _slots_36_io_out_uop_fp_val : _GEN_697 ? _slots_35_io_out_uop_fp_val : _GEN_696 ? _slots_34_io_out_uop_fp_val : _slots_33_io_out_uop_fp_val),
    .io_valid                       (_slots_32_io_valid),
    .io_will_be_valid               (_slots_32_io_will_be_valid),
    .io_request                     (_slots_32_io_request),
    .io_out_uop_uopc                (_slots_32_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_32_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_32_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_32_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_32_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_32_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_32_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_32_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_32_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_32_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_32_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_32_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_32_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_32_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_32_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_32_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_32_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_32_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_32_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_32_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_32_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_32_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_32_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_32_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_32_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_32_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_32_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_32_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_32_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_32_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_32_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_32_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_32_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_32_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_32_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_32_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_32_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_32_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_32_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_32_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_32_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_32_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_32_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_32_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_32_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_32_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_32_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_32_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_32_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_32_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_32_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_32_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_32_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_32_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_32_io_uop_pc_lob),
    .io_uop_taken                   (_slots_32_io_uop_taken),
    .io_uop_imm_packed              (_slots_32_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_32_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_32_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_32_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_32_io_uop_pdst),
    .io_uop_prs1                    (_slots_32_io_uop_prs1),
    .io_uop_prs2                    (_slots_32_io_uop_prs2),
    .io_uop_bypassable              (_slots_32_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_32_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_32_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_32_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_32_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_32_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_32_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_32_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_32_io_uop_fp_val)
  );
  IssueSlot_32 slots_33 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_33_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_85),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_33_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_701 ? _slots_37_io_out_uop_uopc : _GEN_700 ? _slots_36_io_out_uop_uopc : _GEN_699 ? _slots_35_io_out_uop_uopc : _slots_34_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_701 ? _slots_37_io_out_uop_is_rvc : _GEN_700 ? _slots_36_io_out_uop_is_rvc : _GEN_699 ? _slots_35_io_out_uop_is_rvc : _slots_34_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_701 ? _slots_37_io_out_uop_fu_code : _GEN_700 ? _slots_36_io_out_uop_fu_code : _GEN_699 ? _slots_35_io_out_uop_fu_code : _slots_34_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_701 ? _slots_37_io_out_uop_iw_state : _GEN_700 ? _slots_36_io_out_uop_iw_state : _GEN_699 ? _slots_35_io_out_uop_iw_state : _slots_34_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_701 ? _slots_37_io_out_uop_iw_p1_poisoned : _GEN_700 ? _slots_36_io_out_uop_iw_p1_poisoned : _GEN_699 ? _slots_35_io_out_uop_iw_p1_poisoned : _slots_34_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_701 ? _slots_37_io_out_uop_iw_p2_poisoned : _GEN_700 ? _slots_36_io_out_uop_iw_p2_poisoned : _GEN_699 ? _slots_35_io_out_uop_iw_p2_poisoned : _slots_34_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_701 ? _slots_37_io_out_uop_is_br : _GEN_700 ? _slots_36_io_out_uop_is_br : _GEN_699 ? _slots_35_io_out_uop_is_br : _slots_34_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_701 ? _slots_37_io_out_uop_is_jalr : _GEN_700 ? _slots_36_io_out_uop_is_jalr : _GEN_699 ? _slots_35_io_out_uop_is_jalr : _slots_34_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_701 ? _slots_37_io_out_uop_is_jal : _GEN_700 ? _slots_36_io_out_uop_is_jal : _GEN_699 ? _slots_35_io_out_uop_is_jal : _slots_34_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_701 ? _slots_37_io_out_uop_is_sfb : _GEN_700 ? _slots_36_io_out_uop_is_sfb : _GEN_699 ? _slots_35_io_out_uop_is_sfb : _slots_34_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_701 ? _slots_37_io_out_uop_br_mask : _GEN_700 ? _slots_36_io_out_uop_br_mask : _GEN_699 ? _slots_35_io_out_uop_br_mask : _slots_34_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_701 ? _slots_37_io_out_uop_br_tag : _GEN_700 ? _slots_36_io_out_uop_br_tag : _GEN_699 ? _slots_35_io_out_uop_br_tag : _slots_34_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_701 ? _slots_37_io_out_uop_ftq_idx : _GEN_700 ? _slots_36_io_out_uop_ftq_idx : _GEN_699 ? _slots_35_io_out_uop_ftq_idx : _slots_34_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_701 ? _slots_37_io_out_uop_edge_inst : _GEN_700 ? _slots_36_io_out_uop_edge_inst : _GEN_699 ? _slots_35_io_out_uop_edge_inst : _slots_34_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_701 ? _slots_37_io_out_uop_pc_lob : _GEN_700 ? _slots_36_io_out_uop_pc_lob : _GEN_699 ? _slots_35_io_out_uop_pc_lob : _slots_34_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_701 ? _slots_37_io_out_uop_taken : _GEN_700 ? _slots_36_io_out_uop_taken : _GEN_699 ? _slots_35_io_out_uop_taken : _slots_34_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_701 ? _slots_37_io_out_uop_imm_packed : _GEN_700 ? _slots_36_io_out_uop_imm_packed : _GEN_699 ? _slots_35_io_out_uop_imm_packed : _slots_34_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_701 ? _slots_37_io_out_uop_rob_idx : _GEN_700 ? _slots_36_io_out_uop_rob_idx : _GEN_699 ? _slots_35_io_out_uop_rob_idx : _slots_34_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_701 ? _slots_37_io_out_uop_ldq_idx : _GEN_700 ? _slots_36_io_out_uop_ldq_idx : _GEN_699 ? _slots_35_io_out_uop_ldq_idx : _slots_34_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_701 ? _slots_37_io_out_uop_stq_idx : _GEN_700 ? _slots_36_io_out_uop_stq_idx : _GEN_699 ? _slots_35_io_out_uop_stq_idx : _slots_34_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_701 ? _slots_37_io_out_uop_pdst : _GEN_700 ? _slots_36_io_out_uop_pdst : _GEN_699 ? _slots_35_io_out_uop_pdst : _slots_34_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_701 ? _slots_37_io_out_uop_prs1 : _GEN_700 ? _slots_36_io_out_uop_prs1 : _GEN_699 ? _slots_35_io_out_uop_prs1 : _slots_34_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_701 ? _slots_37_io_out_uop_prs2 : _GEN_700 ? _slots_36_io_out_uop_prs2 : _GEN_699 ? _slots_35_io_out_uop_prs2 : _slots_34_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_701 ? _slots_37_io_out_uop_prs3 : _GEN_700 ? _slots_36_io_out_uop_prs3 : _GEN_699 ? _slots_35_io_out_uop_prs3 : _slots_34_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_701 ? _slots_37_io_out_uop_prs1_busy : _GEN_700 ? _slots_36_io_out_uop_prs1_busy : _GEN_699 ? _slots_35_io_out_uop_prs1_busy : _slots_34_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_701 ? _slots_37_io_out_uop_prs2_busy : _GEN_700 ? _slots_36_io_out_uop_prs2_busy : _GEN_699 ? _slots_35_io_out_uop_prs2_busy : _slots_34_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_701 ? _slots_37_io_out_uop_prs3_busy : _GEN_700 ? _slots_36_io_out_uop_prs3_busy : _GEN_699 ? _slots_35_io_out_uop_prs3_busy : _slots_34_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_701 ? _slots_37_io_out_uop_ppred_busy : _GEN_700 ? _slots_36_io_out_uop_ppred_busy : _GEN_699 ? _slots_35_io_out_uop_ppred_busy : _slots_34_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_701 ? _slots_37_io_out_uop_bypassable : _GEN_700 ? _slots_36_io_out_uop_bypassable : _GEN_699 ? _slots_35_io_out_uop_bypassable : _slots_34_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_701 ? _slots_37_io_out_uop_mem_cmd : _GEN_700 ? _slots_36_io_out_uop_mem_cmd : _GEN_699 ? _slots_35_io_out_uop_mem_cmd : _slots_34_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_701 ? _slots_37_io_out_uop_mem_size : _GEN_700 ? _slots_36_io_out_uop_mem_size : _GEN_699 ? _slots_35_io_out_uop_mem_size : _slots_34_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_701 ? _slots_37_io_out_uop_mem_signed : _GEN_700 ? _slots_36_io_out_uop_mem_signed : _GEN_699 ? _slots_35_io_out_uop_mem_signed : _slots_34_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_701 ? _slots_37_io_out_uop_is_fence : _GEN_700 ? _slots_36_io_out_uop_is_fence : _GEN_699 ? _slots_35_io_out_uop_is_fence : _slots_34_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_701 ? _slots_37_io_out_uop_is_amo : _GEN_700 ? _slots_36_io_out_uop_is_amo : _GEN_699 ? _slots_35_io_out_uop_is_amo : _slots_34_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_701 ? _slots_37_io_out_uop_uses_ldq : _GEN_700 ? _slots_36_io_out_uop_uses_ldq : _GEN_699 ? _slots_35_io_out_uop_uses_ldq : _slots_34_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_701 ? _slots_37_io_out_uop_uses_stq : _GEN_700 ? _slots_36_io_out_uop_uses_stq : _GEN_699 ? _slots_35_io_out_uop_uses_stq : _slots_34_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_701 ? _slots_37_io_out_uop_ldst_val : _GEN_700 ? _slots_36_io_out_uop_ldst_val : _GEN_699 ? _slots_35_io_out_uop_ldst_val : _slots_34_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_701 ? _slots_37_io_out_uop_dst_rtype : _GEN_700 ? _slots_36_io_out_uop_dst_rtype : _GEN_699 ? _slots_35_io_out_uop_dst_rtype : _slots_34_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_701 ? _slots_37_io_out_uop_lrs1_rtype : _GEN_700 ? _slots_36_io_out_uop_lrs1_rtype : _GEN_699 ? _slots_35_io_out_uop_lrs1_rtype : _slots_34_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_701 ? _slots_37_io_out_uop_lrs2_rtype : _GEN_700 ? _slots_36_io_out_uop_lrs2_rtype : _GEN_699 ? _slots_35_io_out_uop_lrs2_rtype : _slots_34_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_701 ? _slots_37_io_out_uop_fp_val : _GEN_700 ? _slots_36_io_out_uop_fp_val : _GEN_699 ? _slots_35_io_out_uop_fp_val : _slots_34_io_out_uop_fp_val),
    .io_valid                       (_slots_33_io_valid),
    .io_will_be_valid               (_slots_33_io_will_be_valid),
    .io_request                     (_slots_33_io_request),
    .io_out_uop_uopc                (_slots_33_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_33_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_33_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_33_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_33_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_33_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_33_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_33_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_33_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_33_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_33_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_33_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_33_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_33_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_33_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_33_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_33_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_33_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_33_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_33_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_33_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_33_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_33_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_33_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_33_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_33_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_33_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_33_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_33_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_33_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_33_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_33_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_33_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_33_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_33_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_33_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_33_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_33_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_33_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_33_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_33_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_33_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_33_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_33_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_33_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_33_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_33_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_33_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_33_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_33_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_33_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_33_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_33_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_33_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_33_io_uop_pc_lob),
    .io_uop_taken                   (_slots_33_io_uop_taken),
    .io_uop_imm_packed              (_slots_33_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_33_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_33_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_33_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_33_io_uop_pdst),
    .io_uop_prs1                    (_slots_33_io_uop_prs1),
    .io_uop_prs2                    (_slots_33_io_uop_prs2),
    .io_uop_bypassable              (_slots_33_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_33_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_33_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_33_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_33_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_33_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_33_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_33_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_33_io_uop_fp_val)
  );
  IssueSlot_32 slots_34 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_34_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_87),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_34_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_704 ? _slots_38_io_out_uop_uopc : _GEN_703 ? _slots_37_io_out_uop_uopc : _GEN_702 ? _slots_36_io_out_uop_uopc : _slots_35_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_704 ? _slots_38_io_out_uop_is_rvc : _GEN_703 ? _slots_37_io_out_uop_is_rvc : _GEN_702 ? _slots_36_io_out_uop_is_rvc : _slots_35_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_704 ? _slots_38_io_out_uop_fu_code : _GEN_703 ? _slots_37_io_out_uop_fu_code : _GEN_702 ? _slots_36_io_out_uop_fu_code : _slots_35_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_704 ? _slots_38_io_out_uop_iw_state : _GEN_703 ? _slots_37_io_out_uop_iw_state : _GEN_702 ? _slots_36_io_out_uop_iw_state : _slots_35_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_704 ? _slots_38_io_out_uop_iw_p1_poisoned : _GEN_703 ? _slots_37_io_out_uop_iw_p1_poisoned : _GEN_702 ? _slots_36_io_out_uop_iw_p1_poisoned : _slots_35_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_704 ? _slots_38_io_out_uop_iw_p2_poisoned : _GEN_703 ? _slots_37_io_out_uop_iw_p2_poisoned : _GEN_702 ? _slots_36_io_out_uop_iw_p2_poisoned : _slots_35_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_704 ? _slots_38_io_out_uop_is_br : _GEN_703 ? _slots_37_io_out_uop_is_br : _GEN_702 ? _slots_36_io_out_uop_is_br : _slots_35_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_704 ? _slots_38_io_out_uop_is_jalr : _GEN_703 ? _slots_37_io_out_uop_is_jalr : _GEN_702 ? _slots_36_io_out_uop_is_jalr : _slots_35_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_704 ? _slots_38_io_out_uop_is_jal : _GEN_703 ? _slots_37_io_out_uop_is_jal : _GEN_702 ? _slots_36_io_out_uop_is_jal : _slots_35_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_704 ? _slots_38_io_out_uop_is_sfb : _GEN_703 ? _slots_37_io_out_uop_is_sfb : _GEN_702 ? _slots_36_io_out_uop_is_sfb : _slots_35_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_704 ? _slots_38_io_out_uop_br_mask : _GEN_703 ? _slots_37_io_out_uop_br_mask : _GEN_702 ? _slots_36_io_out_uop_br_mask : _slots_35_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_704 ? _slots_38_io_out_uop_br_tag : _GEN_703 ? _slots_37_io_out_uop_br_tag : _GEN_702 ? _slots_36_io_out_uop_br_tag : _slots_35_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_704 ? _slots_38_io_out_uop_ftq_idx : _GEN_703 ? _slots_37_io_out_uop_ftq_idx : _GEN_702 ? _slots_36_io_out_uop_ftq_idx : _slots_35_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_704 ? _slots_38_io_out_uop_edge_inst : _GEN_703 ? _slots_37_io_out_uop_edge_inst : _GEN_702 ? _slots_36_io_out_uop_edge_inst : _slots_35_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_704 ? _slots_38_io_out_uop_pc_lob : _GEN_703 ? _slots_37_io_out_uop_pc_lob : _GEN_702 ? _slots_36_io_out_uop_pc_lob : _slots_35_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_704 ? _slots_38_io_out_uop_taken : _GEN_703 ? _slots_37_io_out_uop_taken : _GEN_702 ? _slots_36_io_out_uop_taken : _slots_35_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_704 ? _slots_38_io_out_uop_imm_packed : _GEN_703 ? _slots_37_io_out_uop_imm_packed : _GEN_702 ? _slots_36_io_out_uop_imm_packed : _slots_35_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_704 ? _slots_38_io_out_uop_rob_idx : _GEN_703 ? _slots_37_io_out_uop_rob_idx : _GEN_702 ? _slots_36_io_out_uop_rob_idx : _slots_35_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_704 ? _slots_38_io_out_uop_ldq_idx : _GEN_703 ? _slots_37_io_out_uop_ldq_idx : _GEN_702 ? _slots_36_io_out_uop_ldq_idx : _slots_35_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_704 ? _slots_38_io_out_uop_stq_idx : _GEN_703 ? _slots_37_io_out_uop_stq_idx : _GEN_702 ? _slots_36_io_out_uop_stq_idx : _slots_35_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_704 ? _slots_38_io_out_uop_pdst : _GEN_703 ? _slots_37_io_out_uop_pdst : _GEN_702 ? _slots_36_io_out_uop_pdst : _slots_35_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_704 ? _slots_38_io_out_uop_prs1 : _GEN_703 ? _slots_37_io_out_uop_prs1 : _GEN_702 ? _slots_36_io_out_uop_prs1 : _slots_35_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_704 ? _slots_38_io_out_uop_prs2 : _GEN_703 ? _slots_37_io_out_uop_prs2 : _GEN_702 ? _slots_36_io_out_uop_prs2 : _slots_35_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_704 ? _slots_38_io_out_uop_prs3 : _GEN_703 ? _slots_37_io_out_uop_prs3 : _GEN_702 ? _slots_36_io_out_uop_prs3 : _slots_35_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_704 ? _slots_38_io_out_uop_prs1_busy : _GEN_703 ? _slots_37_io_out_uop_prs1_busy : _GEN_702 ? _slots_36_io_out_uop_prs1_busy : _slots_35_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_704 ? _slots_38_io_out_uop_prs2_busy : _GEN_703 ? _slots_37_io_out_uop_prs2_busy : _GEN_702 ? _slots_36_io_out_uop_prs2_busy : _slots_35_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_704 ? _slots_38_io_out_uop_prs3_busy : _GEN_703 ? _slots_37_io_out_uop_prs3_busy : _GEN_702 ? _slots_36_io_out_uop_prs3_busy : _slots_35_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_704 ? _slots_38_io_out_uop_ppred_busy : _GEN_703 ? _slots_37_io_out_uop_ppred_busy : _GEN_702 ? _slots_36_io_out_uop_ppred_busy : _slots_35_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_704 ? _slots_38_io_out_uop_bypassable : _GEN_703 ? _slots_37_io_out_uop_bypassable : _GEN_702 ? _slots_36_io_out_uop_bypassable : _slots_35_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_704 ? _slots_38_io_out_uop_mem_cmd : _GEN_703 ? _slots_37_io_out_uop_mem_cmd : _GEN_702 ? _slots_36_io_out_uop_mem_cmd : _slots_35_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_704 ? _slots_38_io_out_uop_mem_size : _GEN_703 ? _slots_37_io_out_uop_mem_size : _GEN_702 ? _slots_36_io_out_uop_mem_size : _slots_35_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_704 ? _slots_38_io_out_uop_mem_signed : _GEN_703 ? _slots_37_io_out_uop_mem_signed : _GEN_702 ? _slots_36_io_out_uop_mem_signed : _slots_35_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_704 ? _slots_38_io_out_uop_is_fence : _GEN_703 ? _slots_37_io_out_uop_is_fence : _GEN_702 ? _slots_36_io_out_uop_is_fence : _slots_35_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_704 ? _slots_38_io_out_uop_is_amo : _GEN_703 ? _slots_37_io_out_uop_is_amo : _GEN_702 ? _slots_36_io_out_uop_is_amo : _slots_35_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_704 ? _slots_38_io_out_uop_uses_ldq : _GEN_703 ? _slots_37_io_out_uop_uses_ldq : _GEN_702 ? _slots_36_io_out_uop_uses_ldq : _slots_35_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_704 ? _slots_38_io_out_uop_uses_stq : _GEN_703 ? _slots_37_io_out_uop_uses_stq : _GEN_702 ? _slots_36_io_out_uop_uses_stq : _slots_35_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_704 ? _slots_38_io_out_uop_ldst_val : _GEN_703 ? _slots_37_io_out_uop_ldst_val : _GEN_702 ? _slots_36_io_out_uop_ldst_val : _slots_35_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_704 ? _slots_38_io_out_uop_dst_rtype : _GEN_703 ? _slots_37_io_out_uop_dst_rtype : _GEN_702 ? _slots_36_io_out_uop_dst_rtype : _slots_35_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_704 ? _slots_38_io_out_uop_lrs1_rtype : _GEN_703 ? _slots_37_io_out_uop_lrs1_rtype : _GEN_702 ? _slots_36_io_out_uop_lrs1_rtype : _slots_35_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_704 ? _slots_38_io_out_uop_lrs2_rtype : _GEN_703 ? _slots_37_io_out_uop_lrs2_rtype : _GEN_702 ? _slots_36_io_out_uop_lrs2_rtype : _slots_35_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_704 ? _slots_38_io_out_uop_fp_val : _GEN_703 ? _slots_37_io_out_uop_fp_val : _GEN_702 ? _slots_36_io_out_uop_fp_val : _slots_35_io_out_uop_fp_val),
    .io_valid                       (_slots_34_io_valid),
    .io_will_be_valid               (_slots_34_io_will_be_valid),
    .io_request                     (_slots_34_io_request),
    .io_out_uop_uopc                (_slots_34_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_34_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_34_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_34_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_34_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_34_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_34_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_34_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_34_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_34_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_34_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_34_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_34_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_34_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_34_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_34_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_34_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_34_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_34_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_34_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_34_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_34_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_34_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_34_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_34_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_34_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_34_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_34_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_34_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_34_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_34_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_34_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_34_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_34_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_34_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_34_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_34_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_34_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_34_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_34_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_34_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_34_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_34_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_34_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_34_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_34_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_34_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_34_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_34_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_34_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_34_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_34_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_34_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_34_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_34_io_uop_pc_lob),
    .io_uop_taken                   (_slots_34_io_uop_taken),
    .io_uop_imm_packed              (_slots_34_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_34_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_34_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_34_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_34_io_uop_pdst),
    .io_uop_prs1                    (_slots_34_io_uop_prs1),
    .io_uop_prs2                    (_slots_34_io_uop_prs2),
    .io_uop_bypassable              (_slots_34_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_34_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_34_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_34_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_34_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_34_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_34_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_34_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_34_io_uop_fp_val)
  );
  IssueSlot_32 slots_35 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_35_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_89),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_35_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_707 ? _slots_39_io_out_uop_uopc : _GEN_706 ? _slots_38_io_out_uop_uopc : _GEN_705 ? _slots_37_io_out_uop_uopc : _slots_36_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_707 ? _slots_39_io_out_uop_is_rvc : _GEN_706 ? _slots_38_io_out_uop_is_rvc : _GEN_705 ? _slots_37_io_out_uop_is_rvc : _slots_36_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_707 ? _slots_39_io_out_uop_fu_code : _GEN_706 ? _slots_38_io_out_uop_fu_code : _GEN_705 ? _slots_37_io_out_uop_fu_code : _slots_36_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_707 ? _slots_39_io_out_uop_iw_state : _GEN_706 ? _slots_38_io_out_uop_iw_state : _GEN_705 ? _slots_37_io_out_uop_iw_state : _slots_36_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (_GEN_707 ? _slots_39_io_out_uop_iw_p1_poisoned : _GEN_706 ? _slots_38_io_out_uop_iw_p1_poisoned : _GEN_705 ? _slots_37_io_out_uop_iw_p1_poisoned : _slots_36_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (_GEN_707 ? _slots_39_io_out_uop_iw_p2_poisoned : _GEN_706 ? _slots_38_io_out_uop_iw_p2_poisoned : _GEN_705 ? _slots_37_io_out_uop_iw_p2_poisoned : _slots_36_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_707 ? _slots_39_io_out_uop_is_br : _GEN_706 ? _slots_38_io_out_uop_is_br : _GEN_705 ? _slots_37_io_out_uop_is_br : _slots_36_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_707 ? _slots_39_io_out_uop_is_jalr : _GEN_706 ? _slots_38_io_out_uop_is_jalr : _GEN_705 ? _slots_37_io_out_uop_is_jalr : _slots_36_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_707 ? _slots_39_io_out_uop_is_jal : _GEN_706 ? _slots_38_io_out_uop_is_jal : _GEN_705 ? _slots_37_io_out_uop_is_jal : _slots_36_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_707 ? _slots_39_io_out_uop_is_sfb : _GEN_706 ? _slots_38_io_out_uop_is_sfb : _GEN_705 ? _slots_37_io_out_uop_is_sfb : _slots_36_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_707 ? _slots_39_io_out_uop_br_mask : _GEN_706 ? _slots_38_io_out_uop_br_mask : _GEN_705 ? _slots_37_io_out_uop_br_mask : _slots_36_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_707 ? _slots_39_io_out_uop_br_tag : _GEN_706 ? _slots_38_io_out_uop_br_tag : _GEN_705 ? _slots_37_io_out_uop_br_tag : _slots_36_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_707 ? _slots_39_io_out_uop_ftq_idx : _GEN_706 ? _slots_38_io_out_uop_ftq_idx : _GEN_705 ? _slots_37_io_out_uop_ftq_idx : _slots_36_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_707 ? _slots_39_io_out_uop_edge_inst : _GEN_706 ? _slots_38_io_out_uop_edge_inst : _GEN_705 ? _slots_37_io_out_uop_edge_inst : _slots_36_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_707 ? _slots_39_io_out_uop_pc_lob : _GEN_706 ? _slots_38_io_out_uop_pc_lob : _GEN_705 ? _slots_37_io_out_uop_pc_lob : _slots_36_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_707 ? _slots_39_io_out_uop_taken : _GEN_706 ? _slots_38_io_out_uop_taken : _GEN_705 ? _slots_37_io_out_uop_taken : _slots_36_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_707 ? _slots_39_io_out_uop_imm_packed : _GEN_706 ? _slots_38_io_out_uop_imm_packed : _GEN_705 ? _slots_37_io_out_uop_imm_packed : _slots_36_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_707 ? _slots_39_io_out_uop_rob_idx : _GEN_706 ? _slots_38_io_out_uop_rob_idx : _GEN_705 ? _slots_37_io_out_uop_rob_idx : _slots_36_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_707 ? _slots_39_io_out_uop_ldq_idx : _GEN_706 ? _slots_38_io_out_uop_ldq_idx : _GEN_705 ? _slots_37_io_out_uop_ldq_idx : _slots_36_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_707 ? _slots_39_io_out_uop_stq_idx : _GEN_706 ? _slots_38_io_out_uop_stq_idx : _GEN_705 ? _slots_37_io_out_uop_stq_idx : _slots_36_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_707 ? _slots_39_io_out_uop_pdst : _GEN_706 ? _slots_38_io_out_uop_pdst : _GEN_705 ? _slots_37_io_out_uop_pdst : _slots_36_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_707 ? _slots_39_io_out_uop_prs1 : _GEN_706 ? _slots_38_io_out_uop_prs1 : _GEN_705 ? _slots_37_io_out_uop_prs1 : _slots_36_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_707 ? _slots_39_io_out_uop_prs2 : _GEN_706 ? _slots_38_io_out_uop_prs2 : _GEN_705 ? _slots_37_io_out_uop_prs2 : _slots_36_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_707 ? _slots_39_io_out_uop_prs3 : _GEN_706 ? _slots_38_io_out_uop_prs3 : _GEN_705 ? _slots_37_io_out_uop_prs3 : _slots_36_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_707 ? _slots_39_io_out_uop_prs1_busy : _GEN_706 ? _slots_38_io_out_uop_prs1_busy : _GEN_705 ? _slots_37_io_out_uop_prs1_busy : _slots_36_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_707 ? _slots_39_io_out_uop_prs2_busy : _GEN_706 ? _slots_38_io_out_uop_prs2_busy : _GEN_705 ? _slots_37_io_out_uop_prs2_busy : _slots_36_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (_GEN_707 ? _slots_39_io_out_uop_prs3_busy : _GEN_706 ? _slots_38_io_out_uop_prs3_busy : _GEN_705 ? _slots_37_io_out_uop_prs3_busy : _slots_36_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (_GEN_707 ? _slots_39_io_out_uop_ppred_busy : _GEN_706 ? _slots_38_io_out_uop_ppred_busy : _GEN_705 ? _slots_37_io_out_uop_ppred_busy : _slots_36_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_707 ? _slots_39_io_out_uop_bypassable : _GEN_706 ? _slots_38_io_out_uop_bypassable : _GEN_705 ? _slots_37_io_out_uop_bypassable : _slots_36_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_707 ? _slots_39_io_out_uop_mem_cmd : _GEN_706 ? _slots_38_io_out_uop_mem_cmd : _GEN_705 ? _slots_37_io_out_uop_mem_cmd : _slots_36_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_707 ? _slots_39_io_out_uop_mem_size : _GEN_706 ? _slots_38_io_out_uop_mem_size : _GEN_705 ? _slots_37_io_out_uop_mem_size : _slots_36_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_707 ? _slots_39_io_out_uop_mem_signed : _GEN_706 ? _slots_38_io_out_uop_mem_signed : _GEN_705 ? _slots_37_io_out_uop_mem_signed : _slots_36_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_707 ? _slots_39_io_out_uop_is_fence : _GEN_706 ? _slots_38_io_out_uop_is_fence : _GEN_705 ? _slots_37_io_out_uop_is_fence : _slots_36_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_707 ? _slots_39_io_out_uop_is_amo : _GEN_706 ? _slots_38_io_out_uop_is_amo : _GEN_705 ? _slots_37_io_out_uop_is_amo : _slots_36_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_707 ? _slots_39_io_out_uop_uses_ldq : _GEN_706 ? _slots_38_io_out_uop_uses_ldq : _GEN_705 ? _slots_37_io_out_uop_uses_ldq : _slots_36_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_707 ? _slots_39_io_out_uop_uses_stq : _GEN_706 ? _slots_38_io_out_uop_uses_stq : _GEN_705 ? _slots_37_io_out_uop_uses_stq : _slots_36_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_707 ? _slots_39_io_out_uop_ldst_val : _GEN_706 ? _slots_38_io_out_uop_ldst_val : _GEN_705 ? _slots_37_io_out_uop_ldst_val : _slots_36_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_707 ? _slots_39_io_out_uop_dst_rtype : _GEN_706 ? _slots_38_io_out_uop_dst_rtype : _GEN_705 ? _slots_37_io_out_uop_dst_rtype : _slots_36_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_707 ? _slots_39_io_out_uop_lrs1_rtype : _GEN_706 ? _slots_38_io_out_uop_lrs1_rtype : _GEN_705 ? _slots_37_io_out_uop_lrs1_rtype : _slots_36_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_707 ? _slots_39_io_out_uop_lrs2_rtype : _GEN_706 ? _slots_38_io_out_uop_lrs2_rtype : _GEN_705 ? _slots_37_io_out_uop_lrs2_rtype : _slots_36_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_707 ? _slots_39_io_out_uop_fp_val : _GEN_706 ? _slots_38_io_out_uop_fp_val : _GEN_705 ? _slots_37_io_out_uop_fp_val : _slots_36_io_out_uop_fp_val),
    .io_valid                       (_slots_35_io_valid),
    .io_will_be_valid               (_slots_35_io_will_be_valid),
    .io_request                     (_slots_35_io_request),
    .io_out_uop_uopc                (_slots_35_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_35_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_35_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_35_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_35_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_35_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_35_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_35_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_35_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_35_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_35_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_35_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_35_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_35_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_35_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_35_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_35_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_35_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_35_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_35_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_35_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_35_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_35_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_35_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_35_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_35_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_35_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_35_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_35_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_35_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_35_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_35_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_35_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_35_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_35_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_35_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_35_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_35_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_35_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_35_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_35_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_35_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_35_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_35_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_35_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_35_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_35_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_35_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_35_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_35_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_35_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_35_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_35_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_35_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_35_io_uop_pc_lob),
    .io_uop_taken                   (_slots_35_io_uop_taken),
    .io_uop_imm_packed              (_slots_35_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_35_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_35_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_35_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_35_io_uop_pdst),
    .io_uop_prs1                    (_slots_35_io_uop_prs1),
    .io_uop_prs2                    (_slots_35_io_uop_prs2),
    .io_uop_bypassable              (_slots_35_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_35_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_35_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_35_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_35_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_35_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_35_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_35_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_35_io_uop_fp_val)
  );
  IssueSlot_32 slots_36 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_36_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_91),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_36_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_710 ? io_dis_uops_0_bits_uopc : _GEN_709 ? _slots_39_io_out_uop_uopc : _GEN_708 ? _slots_38_io_out_uop_uopc : _slots_37_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_710 ? io_dis_uops_0_bits_is_rvc : _GEN_709 ? _slots_39_io_out_uop_is_rvc : _GEN_708 ? _slots_38_io_out_uop_is_rvc : _slots_37_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_710 ? io_dis_uops_0_bits_fu_code : _GEN_709 ? _slots_39_io_out_uop_fu_code : _GEN_708 ? _slots_38_io_out_uop_fu_code : _slots_37_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_710 ? _GEN_12648 : _GEN_709 ? _slots_39_io_out_uop_iw_state : _GEN_708 ? _slots_38_io_out_uop_iw_state : _slots_37_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_710 & (_GEN_709 ? _slots_39_io_out_uop_iw_p1_poisoned : _GEN_708 ? _slots_38_io_out_uop_iw_p1_poisoned : _slots_37_io_out_uop_iw_p1_poisoned)),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_710 & (_GEN_709 ? _slots_39_io_out_uop_iw_p2_poisoned : _GEN_708 ? _slots_38_io_out_uop_iw_p2_poisoned : _slots_37_io_out_uop_iw_p2_poisoned)),
    .io_in_uop_bits_is_br           (_GEN_710 ? io_dis_uops_0_bits_is_br : _GEN_709 ? _slots_39_io_out_uop_is_br : _GEN_708 ? _slots_38_io_out_uop_is_br : _slots_37_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_710 ? io_dis_uops_0_bits_is_jalr : _GEN_709 ? _slots_39_io_out_uop_is_jalr : _GEN_708 ? _slots_38_io_out_uop_is_jalr : _slots_37_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_710 ? io_dis_uops_0_bits_is_jal : _GEN_709 ? _slots_39_io_out_uop_is_jal : _GEN_708 ? _slots_38_io_out_uop_is_jal : _slots_37_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_710 ? io_dis_uops_0_bits_is_sfb : _GEN_709 ? _slots_39_io_out_uop_is_sfb : _GEN_708 ? _slots_38_io_out_uop_is_sfb : _slots_37_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_710 ? io_dis_uops_0_bits_br_mask : _GEN_709 ? _slots_39_io_out_uop_br_mask : _GEN_708 ? _slots_38_io_out_uop_br_mask : _slots_37_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_710 ? io_dis_uops_0_bits_br_tag : _GEN_709 ? _slots_39_io_out_uop_br_tag : _GEN_708 ? _slots_38_io_out_uop_br_tag : _slots_37_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_710 ? io_dis_uops_0_bits_ftq_idx : _GEN_709 ? _slots_39_io_out_uop_ftq_idx : _GEN_708 ? _slots_38_io_out_uop_ftq_idx : _slots_37_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_710 ? io_dis_uops_0_bits_edge_inst : _GEN_709 ? _slots_39_io_out_uop_edge_inst : _GEN_708 ? _slots_38_io_out_uop_edge_inst : _slots_37_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_710 ? io_dis_uops_0_bits_pc_lob : _GEN_709 ? _slots_39_io_out_uop_pc_lob : _GEN_708 ? _slots_38_io_out_uop_pc_lob : _slots_37_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_710 ? io_dis_uops_0_bits_taken : _GEN_709 ? _slots_39_io_out_uop_taken : _GEN_708 ? _slots_38_io_out_uop_taken : _slots_37_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_710 ? io_dis_uops_0_bits_imm_packed : _GEN_709 ? _slots_39_io_out_uop_imm_packed : _GEN_708 ? _slots_38_io_out_uop_imm_packed : _slots_37_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_710 ? io_dis_uops_0_bits_rob_idx : _GEN_709 ? _slots_39_io_out_uop_rob_idx : _GEN_708 ? _slots_38_io_out_uop_rob_idx : _slots_37_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_710 ? io_dis_uops_0_bits_ldq_idx : _GEN_709 ? _slots_39_io_out_uop_ldq_idx : _GEN_708 ? _slots_38_io_out_uop_ldq_idx : _slots_37_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_710 ? io_dis_uops_0_bits_stq_idx : _GEN_709 ? _slots_39_io_out_uop_stq_idx : _GEN_708 ? _slots_38_io_out_uop_stq_idx : _slots_37_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_710 ? io_dis_uops_0_bits_pdst : _GEN_709 ? _slots_39_io_out_uop_pdst : _GEN_708 ? _slots_38_io_out_uop_pdst : _slots_37_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_710 ? io_dis_uops_0_bits_prs1 : _GEN_709 ? _slots_39_io_out_uop_prs1 : _GEN_708 ? _slots_38_io_out_uop_prs1 : _slots_37_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_710 ? io_dis_uops_0_bits_prs2 : _GEN_709 ? _slots_39_io_out_uop_prs2 : _GEN_708 ? _slots_38_io_out_uop_prs2 : _slots_37_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_710 ? io_dis_uops_0_bits_prs3 : _GEN_709 ? _slots_39_io_out_uop_prs3 : _GEN_708 ? _slots_38_io_out_uop_prs3 : _slots_37_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_710 ? io_dis_uops_0_bits_prs1_busy : _GEN_709 ? _slots_39_io_out_uop_prs1_busy : _GEN_708 ? _slots_38_io_out_uop_prs1_busy : _slots_37_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_710 ? _GEN_12623 : _GEN_709 ? _slots_39_io_out_uop_prs2_busy : _GEN_708 ? _slots_38_io_out_uop_prs2_busy : _slots_37_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_710 & (_GEN_709 ? _slots_39_io_out_uop_prs3_busy : _GEN_708 ? _slots_38_io_out_uop_prs3_busy : _slots_37_io_out_uop_prs3_busy)),
    .io_in_uop_bits_ppred_busy      (~_GEN_710 & (_GEN_709 ? _slots_39_io_out_uop_ppred_busy : _GEN_708 ? _slots_38_io_out_uop_ppred_busy : _slots_37_io_out_uop_ppred_busy)),
    .io_in_uop_bits_bypassable      (_GEN_710 ? io_dis_uops_0_bits_bypassable : _GEN_709 ? _slots_39_io_out_uop_bypassable : _GEN_708 ? _slots_38_io_out_uop_bypassable : _slots_37_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_710 ? io_dis_uops_0_bits_mem_cmd : _GEN_709 ? _slots_39_io_out_uop_mem_cmd : _GEN_708 ? _slots_38_io_out_uop_mem_cmd : _slots_37_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_710 ? io_dis_uops_0_bits_mem_size : _GEN_709 ? _slots_39_io_out_uop_mem_size : _GEN_708 ? _slots_38_io_out_uop_mem_size : _slots_37_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_710 ? io_dis_uops_0_bits_mem_signed : _GEN_709 ? _slots_39_io_out_uop_mem_signed : _GEN_708 ? _slots_38_io_out_uop_mem_signed : _slots_37_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_710 ? io_dis_uops_0_bits_is_fence : _GEN_709 ? _slots_39_io_out_uop_is_fence : _GEN_708 ? _slots_38_io_out_uop_is_fence : _slots_37_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_710 ? io_dis_uops_0_bits_is_amo : _GEN_709 ? _slots_39_io_out_uop_is_amo : _GEN_708 ? _slots_38_io_out_uop_is_amo : _slots_37_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_710 ? io_dis_uops_0_bits_uses_ldq : _GEN_709 ? _slots_39_io_out_uop_uses_ldq : _GEN_708 ? _slots_38_io_out_uop_uses_ldq : _slots_37_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_710 ? io_dis_uops_0_bits_uses_stq : _GEN_709 ? _slots_39_io_out_uop_uses_stq : _GEN_708 ? _slots_38_io_out_uop_uses_stq : _slots_37_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_710 ? io_dis_uops_0_bits_ldst_val : _GEN_709 ? _slots_39_io_out_uop_ldst_val : _GEN_708 ? _slots_38_io_out_uop_ldst_val : _slots_37_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_710 ? io_dis_uops_0_bits_dst_rtype : _GEN_709 ? _slots_39_io_out_uop_dst_rtype : _GEN_708 ? _slots_38_io_out_uop_dst_rtype : _slots_37_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_710 ? io_dis_uops_0_bits_lrs1_rtype : _GEN_709 ? _slots_39_io_out_uop_lrs1_rtype : _GEN_708 ? _slots_38_io_out_uop_lrs1_rtype : _slots_37_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_710 ? _GEN_12597 : _GEN_709 ? _slots_39_io_out_uop_lrs2_rtype : _GEN_708 ? _slots_38_io_out_uop_lrs2_rtype : _slots_37_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_710 ? io_dis_uops_0_bits_fp_val : _GEN_709 ? _slots_39_io_out_uop_fp_val : _GEN_708 ? _slots_38_io_out_uop_fp_val : _slots_37_io_out_uop_fp_val),
    .io_valid                       (_slots_36_io_valid),
    .io_will_be_valid               (_slots_36_io_will_be_valid),
    .io_request                     (_slots_36_io_request),
    .io_out_uop_uopc                (_slots_36_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_36_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_36_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_36_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_36_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_36_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_36_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_36_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_36_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_36_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_36_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_36_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_36_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_36_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_36_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_36_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_36_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_36_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_36_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_36_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_36_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_36_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_36_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_36_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_36_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_36_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_36_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_36_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_36_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_36_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_36_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_36_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_36_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_36_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_36_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_36_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_36_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_36_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_36_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_36_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_36_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_36_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_36_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_36_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_36_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_36_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_36_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_36_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_36_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_36_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_36_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_36_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_36_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_36_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_36_io_uop_pc_lob),
    .io_uop_taken                   (_slots_36_io_uop_taken),
    .io_uop_imm_packed              (_slots_36_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_36_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_36_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_36_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_36_io_uop_pdst),
    .io_uop_prs1                    (_slots_36_io_uop_prs1),
    .io_uop_prs2                    (_slots_36_io_uop_prs2),
    .io_uop_bypassable              (_slots_36_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_36_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_36_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_36_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_36_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_36_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_36_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_36_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_36_io_uop_fp_val)
  );
  IssueSlot_32 slots_37 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_37_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_93),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_37_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_713 ? io_dis_uops_1_bits_uopc : _GEN_712 ? io_dis_uops_0_bits_uopc : _GEN_711 ? _slots_39_io_out_uop_uopc : _slots_38_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_713 ? io_dis_uops_1_bits_is_rvc : _GEN_712 ? io_dis_uops_0_bits_is_rvc : _GEN_711 ? _slots_39_io_out_uop_is_rvc : _slots_38_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_713 ? io_dis_uops_1_bits_fu_code : _GEN_712 ? io_dis_uops_0_bits_fu_code : _GEN_711 ? _slots_39_io_out_uop_fu_code : _slots_38_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_713 ? _GEN_7 : _GEN_712 ? _GEN_12648 : _GEN_711 ? _slots_39_io_out_uop_iw_state : _slots_38_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_714 & (_GEN_711 ? _slots_39_io_out_uop_iw_p1_poisoned : _slots_38_io_out_uop_iw_p1_poisoned)),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_714 & (_GEN_711 ? _slots_39_io_out_uop_iw_p2_poisoned : _slots_38_io_out_uop_iw_p2_poisoned)),
    .io_in_uop_bits_is_br           (_GEN_713 ? io_dis_uops_1_bits_is_br : _GEN_712 ? io_dis_uops_0_bits_is_br : _GEN_711 ? _slots_39_io_out_uop_is_br : _slots_38_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_713 ? io_dis_uops_1_bits_is_jalr : _GEN_712 ? io_dis_uops_0_bits_is_jalr : _GEN_711 ? _slots_39_io_out_uop_is_jalr : _slots_38_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_713 ? io_dis_uops_1_bits_is_jal : _GEN_712 ? io_dis_uops_0_bits_is_jal : _GEN_711 ? _slots_39_io_out_uop_is_jal : _slots_38_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_713 ? io_dis_uops_1_bits_is_sfb : _GEN_712 ? io_dis_uops_0_bits_is_sfb : _GEN_711 ? _slots_39_io_out_uop_is_sfb : _slots_38_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_713 ? io_dis_uops_1_bits_br_mask : _GEN_712 ? io_dis_uops_0_bits_br_mask : _GEN_711 ? _slots_39_io_out_uop_br_mask : _slots_38_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_713 ? io_dis_uops_1_bits_br_tag : _GEN_712 ? io_dis_uops_0_bits_br_tag : _GEN_711 ? _slots_39_io_out_uop_br_tag : _slots_38_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_713 ? io_dis_uops_1_bits_ftq_idx : _GEN_712 ? io_dis_uops_0_bits_ftq_idx : _GEN_711 ? _slots_39_io_out_uop_ftq_idx : _slots_38_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_713 ? io_dis_uops_1_bits_edge_inst : _GEN_712 ? io_dis_uops_0_bits_edge_inst : _GEN_711 ? _slots_39_io_out_uop_edge_inst : _slots_38_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_713 ? io_dis_uops_1_bits_pc_lob : _GEN_712 ? io_dis_uops_0_bits_pc_lob : _GEN_711 ? _slots_39_io_out_uop_pc_lob : _slots_38_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_713 ? io_dis_uops_1_bits_taken : _GEN_712 ? io_dis_uops_0_bits_taken : _GEN_711 ? _slots_39_io_out_uop_taken : _slots_38_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_713 ? io_dis_uops_1_bits_imm_packed : _GEN_712 ? io_dis_uops_0_bits_imm_packed : _GEN_711 ? _slots_39_io_out_uop_imm_packed : _slots_38_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_713 ? io_dis_uops_1_bits_rob_idx : _GEN_712 ? io_dis_uops_0_bits_rob_idx : _GEN_711 ? _slots_39_io_out_uop_rob_idx : _slots_38_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_713 ? io_dis_uops_1_bits_ldq_idx : _GEN_712 ? io_dis_uops_0_bits_ldq_idx : _GEN_711 ? _slots_39_io_out_uop_ldq_idx : _slots_38_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_713 ? io_dis_uops_1_bits_stq_idx : _GEN_712 ? io_dis_uops_0_bits_stq_idx : _GEN_711 ? _slots_39_io_out_uop_stq_idx : _slots_38_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_713 ? io_dis_uops_1_bits_pdst : _GEN_712 ? io_dis_uops_0_bits_pdst : _GEN_711 ? _slots_39_io_out_uop_pdst : _slots_38_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_713 ? io_dis_uops_1_bits_prs1 : _GEN_712 ? io_dis_uops_0_bits_prs1 : _GEN_711 ? _slots_39_io_out_uop_prs1 : _slots_38_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_713 ? io_dis_uops_1_bits_prs2 : _GEN_712 ? io_dis_uops_0_bits_prs2 : _GEN_711 ? _slots_39_io_out_uop_prs2 : _slots_38_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_713 ? io_dis_uops_1_bits_prs3 : _GEN_712 ? io_dis_uops_0_bits_prs3 : _GEN_711 ? _slots_39_io_out_uop_prs3 : _slots_38_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_713 ? io_dis_uops_1_bits_prs1_busy : _GEN_712 ? io_dis_uops_0_bits_prs1_busy : _GEN_711 ? _slots_39_io_out_uop_prs1_busy : _slots_38_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_713 ? _GEN_9 : _GEN_712 ? _GEN_12623 : _GEN_711 ? _slots_39_io_out_uop_prs2_busy : _slots_38_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_714 & (_GEN_711 ? _slots_39_io_out_uop_prs3_busy : _slots_38_io_out_uop_prs3_busy)),
    .io_in_uop_bits_ppred_busy      (~_GEN_714 & (_GEN_711 ? _slots_39_io_out_uop_ppred_busy : _slots_38_io_out_uop_ppred_busy)),
    .io_in_uop_bits_bypassable      (_GEN_713 ? io_dis_uops_1_bits_bypassable : _GEN_712 ? io_dis_uops_0_bits_bypassable : _GEN_711 ? _slots_39_io_out_uop_bypassable : _slots_38_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_713 ? io_dis_uops_1_bits_mem_cmd : _GEN_712 ? io_dis_uops_0_bits_mem_cmd : _GEN_711 ? _slots_39_io_out_uop_mem_cmd : _slots_38_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_713 ? io_dis_uops_1_bits_mem_size : _GEN_712 ? io_dis_uops_0_bits_mem_size : _GEN_711 ? _slots_39_io_out_uop_mem_size : _slots_38_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_713 ? io_dis_uops_1_bits_mem_signed : _GEN_712 ? io_dis_uops_0_bits_mem_signed : _GEN_711 ? _slots_39_io_out_uop_mem_signed : _slots_38_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_713 ? io_dis_uops_1_bits_is_fence : _GEN_712 ? io_dis_uops_0_bits_is_fence : _GEN_711 ? _slots_39_io_out_uop_is_fence : _slots_38_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_713 ? io_dis_uops_1_bits_is_amo : _GEN_712 ? io_dis_uops_0_bits_is_amo : _GEN_711 ? _slots_39_io_out_uop_is_amo : _slots_38_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_713 ? io_dis_uops_1_bits_uses_ldq : _GEN_712 ? io_dis_uops_0_bits_uses_ldq : _GEN_711 ? _slots_39_io_out_uop_uses_ldq : _slots_38_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_713 ? io_dis_uops_1_bits_uses_stq : _GEN_712 ? io_dis_uops_0_bits_uses_stq : _GEN_711 ? _slots_39_io_out_uop_uses_stq : _slots_38_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_713 ? io_dis_uops_1_bits_ldst_val : _GEN_712 ? io_dis_uops_0_bits_ldst_val : _GEN_711 ? _slots_39_io_out_uop_ldst_val : _slots_38_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_713 ? io_dis_uops_1_bits_dst_rtype : _GEN_712 ? io_dis_uops_0_bits_dst_rtype : _GEN_711 ? _slots_39_io_out_uop_dst_rtype : _slots_38_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_713 ? io_dis_uops_1_bits_lrs1_rtype : _GEN_712 ? io_dis_uops_0_bits_lrs1_rtype : _GEN_711 ? _slots_39_io_out_uop_lrs1_rtype : _slots_38_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_713 ? _GEN_8 : _GEN_712 ? _GEN_12597 : _GEN_711 ? _slots_39_io_out_uop_lrs2_rtype : _slots_38_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_713 ? io_dis_uops_1_bits_fp_val : _GEN_712 ? io_dis_uops_0_bits_fp_val : _GEN_711 ? _slots_39_io_out_uop_fp_val : _slots_38_io_out_uop_fp_val),
    .io_valid                       (_slots_37_io_valid),
    .io_will_be_valid               (_slots_37_io_will_be_valid),
    .io_request                     (_slots_37_io_request),
    .io_out_uop_uopc                (_slots_37_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_37_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_37_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_37_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_37_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_37_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_37_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_37_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_37_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_37_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_37_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_37_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_37_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_37_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_37_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_37_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_37_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_37_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_37_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_37_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_37_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_37_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_37_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_37_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_37_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_37_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_37_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_37_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_37_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_37_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_37_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_37_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_37_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_37_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_37_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_37_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_37_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_37_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_37_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_37_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_37_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_37_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_37_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_37_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_37_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_37_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_37_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_37_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_37_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_37_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_37_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_37_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_37_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_37_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_37_io_uop_pc_lob),
    .io_uop_taken                   (_slots_37_io_uop_taken),
    .io_uop_imm_packed              (_slots_37_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_37_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_37_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_37_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_37_io_uop_pdst),
    .io_uop_prs1                    (_slots_37_io_uop_prs1),
    .io_uop_prs2                    (_slots_37_io_uop_prs2),
    .io_uop_bypassable              (_slots_37_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_37_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_37_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_37_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_37_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_37_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_37_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_37_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_37_io_uop_fp_val)
  );
  IssueSlot_32 slots_38 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_38_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_95),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_38_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_717 ? io_dis_uops_2_bits_uopc : _GEN_716 ? io_dis_uops_1_bits_uopc : _GEN_715 ? io_dis_uops_0_bits_uopc : _slots_39_io_out_uop_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_717 ? io_dis_uops_2_bits_is_rvc : _GEN_716 ? io_dis_uops_1_bits_is_rvc : _GEN_715 ? io_dis_uops_0_bits_is_rvc : _slots_39_io_out_uop_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_717 ? io_dis_uops_2_bits_fu_code : _GEN_716 ? io_dis_uops_1_bits_fu_code : _GEN_715 ? io_dis_uops_0_bits_fu_code : _slots_39_io_out_uop_fu_code),
    .io_in_uop_bits_iw_state        (_GEN_717 ? (_GEN_6 ? 2'h2 : 2'h1) : _GEN_716 ? _GEN_7 : _GEN_715 ? _GEN_12648 : _slots_39_io_out_uop_iw_state),
    .io_in_uop_bits_iw_p1_poisoned  (~_GEN_718 & _slots_39_io_out_uop_iw_p1_poisoned),
    .io_in_uop_bits_iw_p2_poisoned  (~_GEN_718 & _slots_39_io_out_uop_iw_p2_poisoned),
    .io_in_uop_bits_is_br           (_GEN_717 ? io_dis_uops_2_bits_is_br : _GEN_716 ? io_dis_uops_1_bits_is_br : _GEN_715 ? io_dis_uops_0_bits_is_br : _slots_39_io_out_uop_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_717 ? io_dis_uops_2_bits_is_jalr : _GEN_716 ? io_dis_uops_1_bits_is_jalr : _GEN_715 ? io_dis_uops_0_bits_is_jalr : _slots_39_io_out_uop_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_717 ? io_dis_uops_2_bits_is_jal : _GEN_716 ? io_dis_uops_1_bits_is_jal : _GEN_715 ? io_dis_uops_0_bits_is_jal : _slots_39_io_out_uop_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_717 ? io_dis_uops_2_bits_is_sfb : _GEN_716 ? io_dis_uops_1_bits_is_sfb : _GEN_715 ? io_dis_uops_0_bits_is_sfb : _slots_39_io_out_uop_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_717 ? io_dis_uops_2_bits_br_mask : _GEN_716 ? io_dis_uops_1_bits_br_mask : _GEN_715 ? io_dis_uops_0_bits_br_mask : _slots_39_io_out_uop_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_717 ? io_dis_uops_2_bits_br_tag : _GEN_716 ? io_dis_uops_1_bits_br_tag : _GEN_715 ? io_dis_uops_0_bits_br_tag : _slots_39_io_out_uop_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_717 ? io_dis_uops_2_bits_ftq_idx : _GEN_716 ? io_dis_uops_1_bits_ftq_idx : _GEN_715 ? io_dis_uops_0_bits_ftq_idx : _slots_39_io_out_uop_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_717 ? io_dis_uops_2_bits_edge_inst : _GEN_716 ? io_dis_uops_1_bits_edge_inst : _GEN_715 ? io_dis_uops_0_bits_edge_inst : _slots_39_io_out_uop_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_717 ? io_dis_uops_2_bits_pc_lob : _GEN_716 ? io_dis_uops_1_bits_pc_lob : _GEN_715 ? io_dis_uops_0_bits_pc_lob : _slots_39_io_out_uop_pc_lob),
    .io_in_uop_bits_taken           (_GEN_717 ? io_dis_uops_2_bits_taken : _GEN_716 ? io_dis_uops_1_bits_taken : _GEN_715 ? io_dis_uops_0_bits_taken : _slots_39_io_out_uop_taken),
    .io_in_uop_bits_imm_packed      (_GEN_717 ? io_dis_uops_2_bits_imm_packed : _GEN_716 ? io_dis_uops_1_bits_imm_packed : _GEN_715 ? io_dis_uops_0_bits_imm_packed : _slots_39_io_out_uop_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_717 ? io_dis_uops_2_bits_rob_idx : _GEN_716 ? io_dis_uops_1_bits_rob_idx : _GEN_715 ? io_dis_uops_0_bits_rob_idx : _slots_39_io_out_uop_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_717 ? io_dis_uops_2_bits_ldq_idx : _GEN_716 ? io_dis_uops_1_bits_ldq_idx : _GEN_715 ? io_dis_uops_0_bits_ldq_idx : _slots_39_io_out_uop_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_717 ? io_dis_uops_2_bits_stq_idx : _GEN_716 ? io_dis_uops_1_bits_stq_idx : _GEN_715 ? io_dis_uops_0_bits_stq_idx : _slots_39_io_out_uop_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_717 ? io_dis_uops_2_bits_pdst : _GEN_716 ? io_dis_uops_1_bits_pdst : _GEN_715 ? io_dis_uops_0_bits_pdst : _slots_39_io_out_uop_pdst),
    .io_in_uop_bits_prs1            (_GEN_717 ? io_dis_uops_2_bits_prs1 : _GEN_716 ? io_dis_uops_1_bits_prs1 : _GEN_715 ? io_dis_uops_0_bits_prs1 : _slots_39_io_out_uop_prs1),
    .io_in_uop_bits_prs2            (_GEN_717 ? io_dis_uops_2_bits_prs2 : _GEN_716 ? io_dis_uops_1_bits_prs2 : _GEN_715 ? io_dis_uops_0_bits_prs2 : _slots_39_io_out_uop_prs2),
    .io_in_uop_bits_prs3            (_GEN_717 ? io_dis_uops_2_bits_prs3 : _GEN_716 ? io_dis_uops_1_bits_prs3 : _GEN_715 ? io_dis_uops_0_bits_prs3 : _slots_39_io_out_uop_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_717 ? io_dis_uops_2_bits_prs1_busy : _GEN_716 ? io_dis_uops_1_bits_prs1_busy : _GEN_715 ? io_dis_uops_0_bits_prs1_busy : _slots_39_io_out_uop_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_717 ? _GEN_14 : _GEN_716 ? _GEN_9 : _GEN_715 ? _GEN_12623 : _slots_39_io_out_uop_prs2_busy),
    .io_in_uop_bits_prs3_busy       (~_GEN_718 & _slots_39_io_out_uop_prs3_busy),
    .io_in_uop_bits_ppred_busy      (~_GEN_718 & _slots_39_io_out_uop_ppred_busy),
    .io_in_uop_bits_bypassable      (_GEN_717 ? io_dis_uops_2_bits_bypassable : _GEN_716 ? io_dis_uops_1_bits_bypassable : _GEN_715 ? io_dis_uops_0_bits_bypassable : _slots_39_io_out_uop_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_717 ? io_dis_uops_2_bits_mem_cmd : _GEN_716 ? io_dis_uops_1_bits_mem_cmd : _GEN_715 ? io_dis_uops_0_bits_mem_cmd : _slots_39_io_out_uop_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_717 ? io_dis_uops_2_bits_mem_size : _GEN_716 ? io_dis_uops_1_bits_mem_size : _GEN_715 ? io_dis_uops_0_bits_mem_size : _slots_39_io_out_uop_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_717 ? io_dis_uops_2_bits_mem_signed : _GEN_716 ? io_dis_uops_1_bits_mem_signed : _GEN_715 ? io_dis_uops_0_bits_mem_signed : _slots_39_io_out_uop_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_717 ? io_dis_uops_2_bits_is_fence : _GEN_716 ? io_dis_uops_1_bits_is_fence : _GEN_715 ? io_dis_uops_0_bits_is_fence : _slots_39_io_out_uop_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_717 ? io_dis_uops_2_bits_is_amo : _GEN_716 ? io_dis_uops_1_bits_is_amo : _GEN_715 ? io_dis_uops_0_bits_is_amo : _slots_39_io_out_uop_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_717 ? io_dis_uops_2_bits_uses_ldq : _GEN_716 ? io_dis_uops_1_bits_uses_ldq : _GEN_715 ? io_dis_uops_0_bits_uses_ldq : _slots_39_io_out_uop_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_717 ? io_dis_uops_2_bits_uses_stq : _GEN_716 ? io_dis_uops_1_bits_uses_stq : _GEN_715 ? io_dis_uops_0_bits_uses_stq : _slots_39_io_out_uop_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_717 ? io_dis_uops_2_bits_ldst_val : _GEN_716 ? io_dis_uops_1_bits_ldst_val : _GEN_715 ? io_dis_uops_0_bits_ldst_val : _slots_39_io_out_uop_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_717 ? io_dis_uops_2_bits_dst_rtype : _GEN_716 ? io_dis_uops_1_bits_dst_rtype : _GEN_715 ? io_dis_uops_0_bits_dst_rtype : _slots_39_io_out_uop_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_717 ? io_dis_uops_2_bits_lrs1_rtype : _GEN_716 ? io_dis_uops_1_bits_lrs1_rtype : _GEN_715 ? io_dis_uops_0_bits_lrs1_rtype : _slots_39_io_out_uop_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_717 ? _GEN_13 : _GEN_716 ? _GEN_8 : _GEN_715 ? _GEN_12597 : _slots_39_io_out_uop_lrs2_rtype),
    .io_in_uop_bits_fp_val          (_GEN_717 ? io_dis_uops_2_bits_fp_val : _GEN_716 ? io_dis_uops_1_bits_fp_val : _GEN_715 ? io_dis_uops_0_bits_fp_val : _slots_39_io_out_uop_fp_val),
    .io_valid                       (_slots_38_io_valid),
    .io_will_be_valid               (_slots_38_io_will_be_valid),
    .io_request                     (_slots_38_io_request),
    .io_out_uop_uopc                (_slots_38_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_38_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_38_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_38_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_38_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_38_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_38_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_38_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_38_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_38_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_38_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_38_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_38_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_38_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_38_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_38_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_38_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_38_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_38_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_38_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_38_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_38_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_38_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_38_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_38_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_38_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_38_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_38_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_38_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_38_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_38_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_38_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_38_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_38_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_38_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_38_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_38_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_38_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_38_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_38_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_38_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_38_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_38_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_38_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_38_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_38_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_38_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_38_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_38_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_38_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_38_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_38_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_38_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_38_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_38_io_uop_pc_lob),
    .io_uop_taken                   (_slots_38_io_uop_taken),
    .io_uop_imm_packed              (_slots_38_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_38_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_38_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_38_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_38_io_uop_pdst),
    .io_uop_prs1                    (_slots_38_io_uop_prs1),
    .io_uop_prs2                    (_slots_38_io_uop_prs2),
    .io_uop_bypassable              (_slots_38_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_38_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_38_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_38_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_38_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_38_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_38_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_38_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_38_io_uop_fp_val)
  );
  IssueSlot_32 slots_39 (
    .clock                          (clock),
    .reset                          (reset),
    .io_grant                       (issue_slots_39_grant),
    .io_brupdate_b1_resolve_mask    (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask (io_brupdate_b1_mispredict_mask),
    .io_kill                        (io_flush_pipeline),
    .io_clear                       (|_GEN_97),
    .io_ldspec_miss                 (io_ld_miss),
    .io_wakeup_ports_0_valid        (io_wakeup_ports_0_valid),
    .io_wakeup_ports_0_bits_pdst    (io_wakeup_ports_0_bits_pdst),
    .io_wakeup_ports_1_valid        (io_wakeup_ports_1_valid),
    .io_wakeup_ports_1_bits_pdst    (io_wakeup_ports_1_bits_pdst),
    .io_wakeup_ports_2_valid        (io_wakeup_ports_2_valid),
    .io_wakeup_ports_2_bits_pdst    (io_wakeup_ports_2_bits_pdst),
    .io_wakeup_ports_3_valid        (io_wakeup_ports_3_valid),
    .io_wakeup_ports_3_bits_pdst    (io_wakeup_ports_3_bits_pdst),
    .io_wakeup_ports_4_valid        (io_wakeup_ports_4_valid),
    .io_wakeup_ports_4_bits_pdst    (io_wakeup_ports_4_bits_pdst),
    .io_wakeup_ports_5_valid        (io_wakeup_ports_5_valid),
    .io_wakeup_ports_5_bits_pdst    (io_wakeup_ports_5_bits_pdst),
    .io_wakeup_ports_6_valid        (io_wakeup_ports_6_valid),
    .io_wakeup_ports_6_bits_pdst    (io_wakeup_ports_6_bits_pdst),
    .io_wakeup_ports_7_valid        (io_wakeup_ports_7_valid),
    .io_wakeup_ports_7_bits_pdst    (io_wakeup_ports_7_bits_pdst),
    .io_wakeup_ports_8_valid        (io_wakeup_ports_8_valid),
    .io_wakeup_ports_8_bits_pdst    (io_wakeup_ports_8_bits_pdst),
    .io_wakeup_ports_9_valid        (io_wakeup_ports_9_valid),
    .io_wakeup_ports_9_bits_pdst    (io_wakeup_ports_9_bits_pdst),
    .io_spec_ld_wakeup_0_valid      (io_spec_ld_wakeup_0_valid),
    .io_spec_ld_wakeup_0_bits       (io_spec_ld_wakeup_0_bits),
    .io_spec_ld_wakeup_1_valid      (io_spec_ld_wakeup_1_valid),
    .io_spec_ld_wakeup_1_bits       (io_spec_ld_wakeup_1_bits),
    .io_in_uop_valid                (issue_slots_39_in_uop_valid),
    .io_in_uop_bits_uopc            (_GEN_721 ? io_dis_uops_3_bits_uopc : _GEN_720 ? io_dis_uops_2_bits_uopc : _GEN_719 ? io_dis_uops_1_bits_uopc : io_dis_uops_0_bits_uopc),
    .io_in_uop_bits_is_rvc          (_GEN_721 ? io_dis_uops_3_bits_is_rvc : _GEN_720 ? io_dis_uops_2_bits_is_rvc : _GEN_719 ? io_dis_uops_1_bits_is_rvc : io_dis_uops_0_bits_is_rvc),
    .io_in_uop_bits_fu_code         (_GEN_721 ? io_dis_uops_3_bits_fu_code : _GEN_720 ? io_dis_uops_2_bits_fu_code : _GEN_719 ? io_dis_uops_1_bits_fu_code : io_dis_uops_0_bits_fu_code),
    .io_in_uop_bits_iw_state        ((_GEN_721 ? _GEN_12 : _GEN_720 ? _GEN_6 : _GEN_719 ? _GEN_3 : _GEN_0) ? 2'h2 : 2'h1),
    .io_in_uop_bits_iw_p1_poisoned  (1'h0),
    .io_in_uop_bits_iw_p2_poisoned  (1'h0),
    .io_in_uop_bits_is_br           (_GEN_721 ? io_dis_uops_3_bits_is_br : _GEN_720 ? io_dis_uops_2_bits_is_br : _GEN_719 ? io_dis_uops_1_bits_is_br : io_dis_uops_0_bits_is_br),
    .io_in_uop_bits_is_jalr         (_GEN_721 ? io_dis_uops_3_bits_is_jalr : _GEN_720 ? io_dis_uops_2_bits_is_jalr : _GEN_719 ? io_dis_uops_1_bits_is_jalr : io_dis_uops_0_bits_is_jalr),
    .io_in_uop_bits_is_jal          (_GEN_721 ? io_dis_uops_3_bits_is_jal : _GEN_720 ? io_dis_uops_2_bits_is_jal : _GEN_719 ? io_dis_uops_1_bits_is_jal : io_dis_uops_0_bits_is_jal),
    .io_in_uop_bits_is_sfb          (_GEN_721 ? io_dis_uops_3_bits_is_sfb : _GEN_720 ? io_dis_uops_2_bits_is_sfb : _GEN_719 ? io_dis_uops_1_bits_is_sfb : io_dis_uops_0_bits_is_sfb),
    .io_in_uop_bits_br_mask         (_GEN_721 ? io_dis_uops_3_bits_br_mask : _GEN_720 ? io_dis_uops_2_bits_br_mask : _GEN_719 ? io_dis_uops_1_bits_br_mask : io_dis_uops_0_bits_br_mask),
    .io_in_uop_bits_br_tag          (_GEN_721 ? io_dis_uops_3_bits_br_tag : _GEN_720 ? io_dis_uops_2_bits_br_tag : _GEN_719 ? io_dis_uops_1_bits_br_tag : io_dis_uops_0_bits_br_tag),
    .io_in_uop_bits_ftq_idx         (_GEN_721 ? io_dis_uops_3_bits_ftq_idx : _GEN_720 ? io_dis_uops_2_bits_ftq_idx : _GEN_719 ? io_dis_uops_1_bits_ftq_idx : io_dis_uops_0_bits_ftq_idx),
    .io_in_uop_bits_edge_inst       (_GEN_721 ? io_dis_uops_3_bits_edge_inst : _GEN_720 ? io_dis_uops_2_bits_edge_inst : _GEN_719 ? io_dis_uops_1_bits_edge_inst : io_dis_uops_0_bits_edge_inst),
    .io_in_uop_bits_pc_lob          (_GEN_721 ? io_dis_uops_3_bits_pc_lob : _GEN_720 ? io_dis_uops_2_bits_pc_lob : _GEN_719 ? io_dis_uops_1_bits_pc_lob : io_dis_uops_0_bits_pc_lob),
    .io_in_uop_bits_taken           (_GEN_721 ? io_dis_uops_3_bits_taken : _GEN_720 ? io_dis_uops_2_bits_taken : _GEN_719 ? io_dis_uops_1_bits_taken : io_dis_uops_0_bits_taken),
    .io_in_uop_bits_imm_packed      (_GEN_721 ? io_dis_uops_3_bits_imm_packed : _GEN_720 ? io_dis_uops_2_bits_imm_packed : _GEN_719 ? io_dis_uops_1_bits_imm_packed : io_dis_uops_0_bits_imm_packed),
    .io_in_uop_bits_rob_idx         (_GEN_721 ? io_dis_uops_3_bits_rob_idx : _GEN_720 ? io_dis_uops_2_bits_rob_idx : _GEN_719 ? io_dis_uops_1_bits_rob_idx : io_dis_uops_0_bits_rob_idx),
    .io_in_uop_bits_ldq_idx         (_GEN_721 ? io_dis_uops_3_bits_ldq_idx : _GEN_720 ? io_dis_uops_2_bits_ldq_idx : _GEN_719 ? io_dis_uops_1_bits_ldq_idx : io_dis_uops_0_bits_ldq_idx),
    .io_in_uop_bits_stq_idx         (_GEN_721 ? io_dis_uops_3_bits_stq_idx : _GEN_720 ? io_dis_uops_2_bits_stq_idx : _GEN_719 ? io_dis_uops_1_bits_stq_idx : io_dis_uops_0_bits_stq_idx),
    .io_in_uop_bits_pdst            (_GEN_721 ? io_dis_uops_3_bits_pdst : _GEN_720 ? io_dis_uops_2_bits_pdst : _GEN_719 ? io_dis_uops_1_bits_pdst : io_dis_uops_0_bits_pdst),
    .io_in_uop_bits_prs1            (_GEN_721 ? io_dis_uops_3_bits_prs1 : _GEN_720 ? io_dis_uops_2_bits_prs1 : _GEN_719 ? io_dis_uops_1_bits_prs1 : io_dis_uops_0_bits_prs1),
    .io_in_uop_bits_prs2            (_GEN_721 ? io_dis_uops_3_bits_prs2 : _GEN_720 ? io_dis_uops_2_bits_prs2 : _GEN_719 ? io_dis_uops_1_bits_prs2 : io_dis_uops_0_bits_prs2),
    .io_in_uop_bits_prs3            (_GEN_721 ? io_dis_uops_3_bits_prs3 : _GEN_720 ? io_dis_uops_2_bits_prs3 : _GEN_719 ? io_dis_uops_1_bits_prs3 : io_dis_uops_0_bits_prs3),
    .io_in_uop_bits_prs1_busy       (_GEN_721 ? io_dis_uops_3_bits_prs1_busy : _GEN_720 ? io_dis_uops_2_bits_prs1_busy : _GEN_719 ? io_dis_uops_1_bits_prs1_busy : io_dis_uops_0_bits_prs1_busy),
    .io_in_uop_bits_prs2_busy       (_GEN_721 ? _GEN_15 & io_dis_uops_3_bits_prs2_busy : _GEN_720 ? _GEN_14 : _GEN_719 ? _GEN_9 : _GEN_12623),
    .io_in_uop_bits_prs3_busy       (1'h0),
    .io_in_uop_bits_ppred_busy      (1'h0),
    .io_in_uop_bits_bypassable      (_GEN_721 ? io_dis_uops_3_bits_bypassable : _GEN_720 ? io_dis_uops_2_bits_bypassable : _GEN_719 ? io_dis_uops_1_bits_bypassable : io_dis_uops_0_bits_bypassable),
    .io_in_uop_bits_mem_cmd         (_GEN_721 ? io_dis_uops_3_bits_mem_cmd : _GEN_720 ? io_dis_uops_2_bits_mem_cmd : _GEN_719 ? io_dis_uops_1_bits_mem_cmd : io_dis_uops_0_bits_mem_cmd),
    .io_in_uop_bits_mem_size        (_GEN_721 ? io_dis_uops_3_bits_mem_size : _GEN_720 ? io_dis_uops_2_bits_mem_size : _GEN_719 ? io_dis_uops_1_bits_mem_size : io_dis_uops_0_bits_mem_size),
    .io_in_uop_bits_mem_signed      (_GEN_721 ? io_dis_uops_3_bits_mem_signed : _GEN_720 ? io_dis_uops_2_bits_mem_signed : _GEN_719 ? io_dis_uops_1_bits_mem_signed : io_dis_uops_0_bits_mem_signed),
    .io_in_uop_bits_is_fence        (_GEN_721 ? io_dis_uops_3_bits_is_fence : _GEN_720 ? io_dis_uops_2_bits_is_fence : _GEN_719 ? io_dis_uops_1_bits_is_fence : io_dis_uops_0_bits_is_fence),
    .io_in_uop_bits_is_amo          (_GEN_721 ? io_dis_uops_3_bits_is_amo : _GEN_720 ? io_dis_uops_2_bits_is_amo : _GEN_719 ? io_dis_uops_1_bits_is_amo : io_dis_uops_0_bits_is_amo),
    .io_in_uop_bits_uses_ldq        (_GEN_721 ? io_dis_uops_3_bits_uses_ldq : _GEN_720 ? io_dis_uops_2_bits_uses_ldq : _GEN_719 ? io_dis_uops_1_bits_uses_ldq : io_dis_uops_0_bits_uses_ldq),
    .io_in_uop_bits_uses_stq        (_GEN_721 ? io_dis_uops_3_bits_uses_stq : _GEN_720 ? io_dis_uops_2_bits_uses_stq : _GEN_719 ? io_dis_uops_1_bits_uses_stq : io_dis_uops_0_bits_uses_stq),
    .io_in_uop_bits_ldst_val        (_GEN_721 ? io_dis_uops_3_bits_ldst_val : _GEN_720 ? io_dis_uops_2_bits_ldst_val : _GEN_719 ? io_dis_uops_1_bits_ldst_val : io_dis_uops_0_bits_ldst_val),
    .io_in_uop_bits_dst_rtype       (_GEN_721 ? io_dis_uops_3_bits_dst_rtype : _GEN_720 ? io_dis_uops_2_bits_dst_rtype : _GEN_719 ? io_dis_uops_1_bits_dst_rtype : io_dis_uops_0_bits_dst_rtype),
    .io_in_uop_bits_lrs1_rtype      (_GEN_721 ? io_dis_uops_3_bits_lrs1_rtype : _GEN_720 ? io_dis_uops_2_bits_lrs1_rtype : _GEN_719 ? io_dis_uops_1_bits_lrs1_rtype : io_dis_uops_0_bits_lrs1_rtype),
    .io_in_uop_bits_lrs2_rtype      (_GEN_721 ? (_GEN_15 ? io_dis_uops_3_bits_lrs2_rtype : 2'h2) : _GEN_720 ? _GEN_13 : _GEN_719 ? _GEN_8 : _GEN_12597),
    .io_in_uop_bits_fp_val          (_GEN_721 ? io_dis_uops_3_bits_fp_val : _GEN_720 ? io_dis_uops_2_bits_fp_val : _GEN_719 ? io_dis_uops_1_bits_fp_val : io_dis_uops_0_bits_fp_val),
    .io_valid                       (_slots_39_io_valid),
    .io_will_be_valid               (_slots_39_io_will_be_valid),
    .io_request                     (_slots_39_io_request),
    .io_out_uop_uopc                (_slots_39_io_out_uop_uopc),
    .io_out_uop_is_rvc              (_slots_39_io_out_uop_is_rvc),
    .io_out_uop_fu_code             (_slots_39_io_out_uop_fu_code),
    .io_out_uop_iw_state            (_slots_39_io_out_uop_iw_state),
    .io_out_uop_iw_p1_poisoned      (_slots_39_io_out_uop_iw_p1_poisoned),
    .io_out_uop_iw_p2_poisoned      (_slots_39_io_out_uop_iw_p2_poisoned),
    .io_out_uop_is_br               (_slots_39_io_out_uop_is_br),
    .io_out_uop_is_jalr             (_slots_39_io_out_uop_is_jalr),
    .io_out_uop_is_jal              (_slots_39_io_out_uop_is_jal),
    .io_out_uop_is_sfb              (_slots_39_io_out_uop_is_sfb),
    .io_out_uop_br_mask             (_slots_39_io_out_uop_br_mask),
    .io_out_uop_br_tag              (_slots_39_io_out_uop_br_tag),
    .io_out_uop_ftq_idx             (_slots_39_io_out_uop_ftq_idx),
    .io_out_uop_edge_inst           (_slots_39_io_out_uop_edge_inst),
    .io_out_uop_pc_lob              (_slots_39_io_out_uop_pc_lob),
    .io_out_uop_taken               (_slots_39_io_out_uop_taken),
    .io_out_uop_imm_packed          (_slots_39_io_out_uop_imm_packed),
    .io_out_uop_rob_idx             (_slots_39_io_out_uop_rob_idx),
    .io_out_uop_ldq_idx             (_slots_39_io_out_uop_ldq_idx),
    .io_out_uop_stq_idx             (_slots_39_io_out_uop_stq_idx),
    .io_out_uop_pdst                (_slots_39_io_out_uop_pdst),
    .io_out_uop_prs1                (_slots_39_io_out_uop_prs1),
    .io_out_uop_prs2                (_slots_39_io_out_uop_prs2),
    .io_out_uop_prs3                (_slots_39_io_out_uop_prs3),
    .io_out_uop_prs1_busy           (_slots_39_io_out_uop_prs1_busy),
    .io_out_uop_prs2_busy           (_slots_39_io_out_uop_prs2_busy),
    .io_out_uop_prs3_busy           (_slots_39_io_out_uop_prs3_busy),
    .io_out_uop_ppred_busy          (_slots_39_io_out_uop_ppred_busy),
    .io_out_uop_bypassable          (_slots_39_io_out_uop_bypassable),
    .io_out_uop_mem_cmd             (_slots_39_io_out_uop_mem_cmd),
    .io_out_uop_mem_size            (_slots_39_io_out_uop_mem_size),
    .io_out_uop_mem_signed          (_slots_39_io_out_uop_mem_signed),
    .io_out_uop_is_fence            (_slots_39_io_out_uop_is_fence),
    .io_out_uop_is_amo              (_slots_39_io_out_uop_is_amo),
    .io_out_uop_uses_ldq            (_slots_39_io_out_uop_uses_ldq),
    .io_out_uop_uses_stq            (_slots_39_io_out_uop_uses_stq),
    .io_out_uop_ldst_val            (_slots_39_io_out_uop_ldst_val),
    .io_out_uop_dst_rtype           (_slots_39_io_out_uop_dst_rtype),
    .io_out_uop_lrs1_rtype          (_slots_39_io_out_uop_lrs1_rtype),
    .io_out_uop_lrs2_rtype          (_slots_39_io_out_uop_lrs2_rtype),
    .io_out_uop_fp_val              (_slots_39_io_out_uop_fp_val),
    .io_uop_uopc                    (_slots_39_io_uop_uopc),
    .io_uop_is_rvc                  (_slots_39_io_uop_is_rvc),
    .io_uop_fu_code                 (_slots_39_io_uop_fu_code),
    .io_uop_iw_p1_poisoned          (_slots_39_io_uop_iw_p1_poisoned),
    .io_uop_iw_p2_poisoned          (_slots_39_io_uop_iw_p2_poisoned),
    .io_uop_is_br                   (_slots_39_io_uop_is_br),
    .io_uop_is_jalr                 (_slots_39_io_uop_is_jalr),
    .io_uop_is_jal                  (_slots_39_io_uop_is_jal),
    .io_uop_is_sfb                  (_slots_39_io_uop_is_sfb),
    .io_uop_br_mask                 (_slots_39_io_uop_br_mask),
    .io_uop_br_tag                  (_slots_39_io_uop_br_tag),
    .io_uop_ftq_idx                 (_slots_39_io_uop_ftq_idx),
    .io_uop_edge_inst               (_slots_39_io_uop_edge_inst),
    .io_uop_pc_lob                  (_slots_39_io_uop_pc_lob),
    .io_uop_taken                   (_slots_39_io_uop_taken),
    .io_uop_imm_packed              (_slots_39_io_uop_imm_packed),
    .io_uop_rob_idx                 (_slots_39_io_uop_rob_idx),
    .io_uop_ldq_idx                 (_slots_39_io_uop_ldq_idx),
    .io_uop_stq_idx                 (_slots_39_io_uop_stq_idx),
    .io_uop_pdst                    (_slots_39_io_uop_pdst),
    .io_uop_prs1                    (_slots_39_io_uop_prs1),
    .io_uop_prs2                    (_slots_39_io_uop_prs2),
    .io_uop_bypassable              (_slots_39_io_uop_bypassable),
    .io_uop_mem_cmd                 (_slots_39_io_uop_mem_cmd),
    .io_uop_mem_size                (/* unused */),
    .io_uop_mem_signed              (/* unused */),
    .io_uop_is_fence                (/* unused */),
    .io_uop_is_amo                  (_slots_39_io_uop_is_amo),
    .io_uop_uses_ldq                (/* unused */),
    .io_uop_uses_stq                (_slots_39_io_uop_uses_stq),
    .io_uop_ldst_val                (_slots_39_io_uop_ldst_val),
    .io_uop_dst_rtype               (_slots_39_io_uop_dst_rtype),
    .io_uop_lrs1_rtype              (_slots_39_io_uop_lrs1_rtype),
    .io_uop_lrs2_rtype              (_slots_39_io_uop_lrs2_rtype),
    .io_uop_fp_val                  (_slots_39_io_uop_fp_val)
  );
  assign io_dis_uops_0_ready = io_dis_uops_0_ready_REG;
  assign io_dis_uops_1_ready = io_dis_uops_1_ready_REG;
  assign io_dis_uops_2_ready = io_dis_uops_2_ready_REG;
  assign io_dis_uops_3_ready = io_dis_uops_3_ready_REG;
  assign io_iss_valids_0 = _GEN_25541 | _GEN_25217 | _GEN_24893 | _GEN_24569 | _GEN_24245 | _GEN_23921 | _GEN_23597 | _GEN_23273 | _GEN_22949 | _GEN_22625 | _GEN_22301 | _GEN_21977 | _GEN_21653 | _GEN_21329 | _GEN_21005 | _GEN_20681 | _GEN_20357 | _GEN_20033 | _GEN_19709 | _GEN_19385 | _GEN_19061 | _GEN_18737 | _GEN_18413 | _GEN_18089 | _GEN_17765 | _GEN_17441 | _GEN_17117 | _GEN_16793 | _GEN_16469 | _GEN_16145 | _GEN_15821 | _GEN_15497 | _GEN_15173 | _GEN_14849 | _GEN_14525 | _GEN_14201 | _GEN_13877 | _GEN_13553 | _GEN_13229 | _GEN_12906;
  assign io_iss_valids_1 = _GEN_596 | _GEN_586 | _GEN_599 | _GEN_561 | _GEN_547 | _GEN_530 | _GEN_516 | _GEN_533 | _GEN_491 | _GEN_477 | _GEN_460 | _GEN_446 | _GEN_463 | _GEN_421 | _GEN_407 | _GEN_390 | _GEN_376 | _GEN_393 | _GEN_351 | _GEN_337 | _GEN_320 | _GEN_306 | _GEN_323 | _GEN_281 | _GEN_267 | _GEN_250 | _GEN_236 | _GEN_253 | _GEN_211 | _GEN_197 | _GEN_180 | _GEN_166 | _GEN_183 | _GEN_141 | _GEN_127 | _GEN_110 | _GEN_94 | _GEN_113 | _GEN_44 | _GEN_12987;
  assign io_iss_valids_2 = _GEN_595 | _GEN_584 | _GEN_598 | _GEN_559 | _GEN_545 | _GEN_528 | _GEN_514 | _GEN_532 | _GEN_489 | _GEN_475 | _GEN_458 | _GEN_444 | _GEN_462 | _GEN_419 | _GEN_405 | _GEN_388 | _GEN_374 | _GEN_392 | _GEN_349 | _GEN_335 | _GEN_318 | _GEN_304 | _GEN_322 | _GEN_279 | _GEN_265 | _GEN_248 | _GEN_234 | _GEN_252 | _GEN_209 | _GEN_195 | _GEN_178 | _GEN_164 | _GEN_182 | _GEN_139 | _GEN_125 | _GEN_108 | _GEN_90 | _GEN_112 | _GEN_40 | _GEN_13068;
  assign io_iss_valids_3 = _GEN_594 | _GEN_582 | _GEN_597 | _GEN_557 | _GEN_543 | _GEN_526 | _GEN_512 | _GEN_531 | _GEN_487 | _GEN_473 | _GEN_456 | _GEN_442 | _GEN_461 | _GEN_417 | _GEN_403 | _GEN_386 | _GEN_372 | _GEN_391 | _GEN_347 | _GEN_333 | _GEN_316 | _GEN_302 | _GEN_321 | _GEN_277 | _GEN_263 | _GEN_246 | _GEN_232 | _GEN_251 | _GEN_207 | _GEN_193 | _GEN_176 | _GEN_162 | _GEN_181 | _GEN_137 | _GEN_123 | _GEN_106 | _GEN_86 | _GEN_111 | _GEN_36 | _GEN_13149;
  assign io_iss_uops_0_uopc = _GEN_25541 ? _slots_39_io_uop_uopc : _GEN_25217 ? _slots_38_io_uop_uopc : _GEN_24893 ? _slots_37_io_uop_uopc : _GEN_24569 ? _slots_36_io_uop_uopc : _GEN_24245 ? _slots_35_io_uop_uopc : _GEN_23921 ? _slots_34_io_uop_uopc : _GEN_23597 ? _slots_33_io_uop_uopc : _GEN_23273 ? _slots_32_io_uop_uopc : _GEN_22949 ? _slots_31_io_uop_uopc : _GEN_22625 ? _slots_30_io_uop_uopc : _GEN_22301 ? _slots_29_io_uop_uopc : _GEN_21977 ? _slots_28_io_uop_uopc : _GEN_21653 ? _slots_27_io_uop_uopc : _GEN_21329 ? _slots_26_io_uop_uopc : _GEN_21005 ? _slots_25_io_uop_uopc : _GEN_20681 ? _slots_24_io_uop_uopc : _GEN_20357 ? _slots_23_io_uop_uopc : _GEN_20033 ? _slots_22_io_uop_uopc : _GEN_19709 ? _slots_21_io_uop_uopc : _GEN_19385 ? _slots_20_io_uop_uopc : _GEN_19061 ? _slots_19_io_uop_uopc : _GEN_18737 ? _slots_18_io_uop_uopc : _GEN_18413 ? _slots_17_io_uop_uopc : _GEN_18089 ? _slots_16_io_uop_uopc : _GEN_17765 ? _slots_15_io_uop_uopc : _GEN_17441 ? _slots_14_io_uop_uopc : _GEN_17117 ? _slots_13_io_uop_uopc : _GEN_16793 ? _slots_12_io_uop_uopc : _GEN_16469 ? _slots_11_io_uop_uopc : _GEN_16145 ? _slots_10_io_uop_uopc : _GEN_15821 ? _slots_9_io_uop_uopc : _GEN_15497 ? _slots_8_io_uop_uopc : _GEN_15173 ? _slots_7_io_uop_uopc : _GEN_14849 ? _slots_6_io_uop_uopc : _GEN_14525 ? _slots_5_io_uop_uopc : _GEN_14201 ? _slots_4_io_uop_uopc : _GEN_13877 ? _slots_3_io_uop_uopc : _GEN_13553 ? _slots_2_io_uop_uopc : _GEN_13229 ? _slots_1_io_uop_uopc : _GEN_12906 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_0_is_rvc = _GEN_25541 ? _slots_39_io_uop_is_rvc : _GEN_25217 ? _slots_38_io_uop_is_rvc : _GEN_24893 ? _slots_37_io_uop_is_rvc : _GEN_24569 ? _slots_36_io_uop_is_rvc : _GEN_24245 ? _slots_35_io_uop_is_rvc : _GEN_23921 ? _slots_34_io_uop_is_rvc : _GEN_23597 ? _slots_33_io_uop_is_rvc : _GEN_23273 ? _slots_32_io_uop_is_rvc : _GEN_22949 ? _slots_31_io_uop_is_rvc : _GEN_22625 ? _slots_30_io_uop_is_rvc : _GEN_22301 ? _slots_29_io_uop_is_rvc : _GEN_21977 ? _slots_28_io_uop_is_rvc : _GEN_21653 ? _slots_27_io_uop_is_rvc : _GEN_21329 ? _slots_26_io_uop_is_rvc : _GEN_21005 ? _slots_25_io_uop_is_rvc : _GEN_20681 ? _slots_24_io_uop_is_rvc : _GEN_20357 ? _slots_23_io_uop_is_rvc : _GEN_20033 ? _slots_22_io_uop_is_rvc : _GEN_19709 ? _slots_21_io_uop_is_rvc : _GEN_19385 ? _slots_20_io_uop_is_rvc : _GEN_19061 ? _slots_19_io_uop_is_rvc : _GEN_18737 ? _slots_18_io_uop_is_rvc : _GEN_18413 ? _slots_17_io_uop_is_rvc : _GEN_18089 ? _slots_16_io_uop_is_rvc : _GEN_17765 ? _slots_15_io_uop_is_rvc : _GEN_17441 ? _slots_14_io_uop_is_rvc : _GEN_17117 ? _slots_13_io_uop_is_rvc : _GEN_16793 ? _slots_12_io_uop_is_rvc : _GEN_16469 ? _slots_11_io_uop_is_rvc : _GEN_16145 ? _slots_10_io_uop_is_rvc : _GEN_15821 ? _slots_9_io_uop_is_rvc : _GEN_15497 ? _slots_8_io_uop_is_rvc : _GEN_15173 ? _slots_7_io_uop_is_rvc : _GEN_14849 ? _slots_6_io_uop_is_rvc : _GEN_14525 ? _slots_5_io_uop_is_rvc : _GEN_14201 ? _slots_4_io_uop_is_rvc : _GEN_13877 ? _slots_3_io_uop_is_rvc : _GEN_13553 ? _slots_2_io_uop_is_rvc : _GEN_13229 ? _slots_1_io_uop_is_rvc : _GEN_12906 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_0_fu_code = _GEN_25541 ? _slots_39_io_uop_fu_code : _GEN_25217 ? _slots_38_io_uop_fu_code : _GEN_24893 ? _slots_37_io_uop_fu_code : _GEN_24569 ? _slots_36_io_uop_fu_code : _GEN_24245 ? _slots_35_io_uop_fu_code : _GEN_23921 ? _slots_34_io_uop_fu_code : _GEN_23597 ? _slots_33_io_uop_fu_code : _GEN_23273 ? _slots_32_io_uop_fu_code : _GEN_22949 ? _slots_31_io_uop_fu_code : _GEN_22625 ? _slots_30_io_uop_fu_code : _GEN_22301 ? _slots_29_io_uop_fu_code : _GEN_21977 ? _slots_28_io_uop_fu_code : _GEN_21653 ? _slots_27_io_uop_fu_code : _GEN_21329 ? _slots_26_io_uop_fu_code : _GEN_21005 ? _slots_25_io_uop_fu_code : _GEN_20681 ? _slots_24_io_uop_fu_code : _GEN_20357 ? _slots_23_io_uop_fu_code : _GEN_20033 ? _slots_22_io_uop_fu_code : _GEN_19709 ? _slots_21_io_uop_fu_code : _GEN_19385 ? _slots_20_io_uop_fu_code : _GEN_19061 ? _slots_19_io_uop_fu_code : _GEN_18737 ? _slots_18_io_uop_fu_code : _GEN_18413 ? _slots_17_io_uop_fu_code : _GEN_18089 ? _slots_16_io_uop_fu_code : _GEN_17765 ? _slots_15_io_uop_fu_code : _GEN_17441 ? _slots_14_io_uop_fu_code : _GEN_17117 ? _slots_13_io_uop_fu_code : _GEN_16793 ? _slots_12_io_uop_fu_code : _GEN_16469 ? _slots_11_io_uop_fu_code : _GEN_16145 ? _slots_10_io_uop_fu_code : _GEN_15821 ? _slots_9_io_uop_fu_code : _GEN_15497 ? _slots_8_io_uop_fu_code : _GEN_15173 ? _slots_7_io_uop_fu_code : _GEN_14849 ? _slots_6_io_uop_fu_code : _GEN_14525 ? _slots_5_io_uop_fu_code : _GEN_14201 ? _slots_4_io_uop_fu_code : _GEN_13877 ? _slots_3_io_uop_fu_code : _GEN_13553 ? _slots_2_io_uop_fu_code : _GEN_13229 ? _slots_1_io_uop_fu_code : _GEN_12906 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_0_iw_p1_poisoned = _GEN_25541 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_25217 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_24893 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_24569 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_24245 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_23921 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_23597 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_23273 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_22949 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_22625 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_22301 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_21977 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_21653 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_21329 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_21005 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_20681 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_20357 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_20033 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_19709 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_19385 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_19061 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_18737 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_18413 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_18089 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_17765 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_17441 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_17117 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_16793 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_16469 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_16145 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_15821 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_15497 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_15173 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_14849 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_14525 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_14201 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_13877 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_13553 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_13229 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_12906 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_0_iw_p2_poisoned = _GEN_25541 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_25217 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_24893 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_24569 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_24245 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_23921 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_23597 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_23273 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_22949 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_22625 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_22301 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_21977 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_21653 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_21329 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_21005 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_20681 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_20357 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_20033 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_19709 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_19385 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_19061 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_18737 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_18413 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_18089 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_17765 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_17441 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_17117 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_16793 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_16469 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_16145 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_15821 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_15497 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_15173 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_14849 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_14525 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_14201 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_13877 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_13553 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_13229 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_12906 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_0_is_br = _GEN_25541 ? _slots_39_io_uop_is_br : _GEN_25217 ? _slots_38_io_uop_is_br : _GEN_24893 ? _slots_37_io_uop_is_br : _GEN_24569 ? _slots_36_io_uop_is_br : _GEN_24245 ? _slots_35_io_uop_is_br : _GEN_23921 ? _slots_34_io_uop_is_br : _GEN_23597 ? _slots_33_io_uop_is_br : _GEN_23273 ? _slots_32_io_uop_is_br : _GEN_22949 ? _slots_31_io_uop_is_br : _GEN_22625 ? _slots_30_io_uop_is_br : _GEN_22301 ? _slots_29_io_uop_is_br : _GEN_21977 ? _slots_28_io_uop_is_br : _GEN_21653 ? _slots_27_io_uop_is_br : _GEN_21329 ? _slots_26_io_uop_is_br : _GEN_21005 ? _slots_25_io_uop_is_br : _GEN_20681 ? _slots_24_io_uop_is_br : _GEN_20357 ? _slots_23_io_uop_is_br : _GEN_20033 ? _slots_22_io_uop_is_br : _GEN_19709 ? _slots_21_io_uop_is_br : _GEN_19385 ? _slots_20_io_uop_is_br : _GEN_19061 ? _slots_19_io_uop_is_br : _GEN_18737 ? _slots_18_io_uop_is_br : _GEN_18413 ? _slots_17_io_uop_is_br : _GEN_18089 ? _slots_16_io_uop_is_br : _GEN_17765 ? _slots_15_io_uop_is_br : _GEN_17441 ? _slots_14_io_uop_is_br : _GEN_17117 ? _slots_13_io_uop_is_br : _GEN_16793 ? _slots_12_io_uop_is_br : _GEN_16469 ? _slots_11_io_uop_is_br : _GEN_16145 ? _slots_10_io_uop_is_br : _GEN_15821 ? _slots_9_io_uop_is_br : _GEN_15497 ? _slots_8_io_uop_is_br : _GEN_15173 ? _slots_7_io_uop_is_br : _GEN_14849 ? _slots_6_io_uop_is_br : _GEN_14525 ? _slots_5_io_uop_is_br : _GEN_14201 ? _slots_4_io_uop_is_br : _GEN_13877 ? _slots_3_io_uop_is_br : _GEN_13553 ? _slots_2_io_uop_is_br : _GEN_13229 ? _slots_1_io_uop_is_br : _GEN_12906 & _slots_0_io_uop_is_br;
  assign io_iss_uops_0_is_jalr = _GEN_25541 ? _slots_39_io_uop_is_jalr : _GEN_25217 ? _slots_38_io_uop_is_jalr : _GEN_24893 ? _slots_37_io_uop_is_jalr : _GEN_24569 ? _slots_36_io_uop_is_jalr : _GEN_24245 ? _slots_35_io_uop_is_jalr : _GEN_23921 ? _slots_34_io_uop_is_jalr : _GEN_23597 ? _slots_33_io_uop_is_jalr : _GEN_23273 ? _slots_32_io_uop_is_jalr : _GEN_22949 ? _slots_31_io_uop_is_jalr : _GEN_22625 ? _slots_30_io_uop_is_jalr : _GEN_22301 ? _slots_29_io_uop_is_jalr : _GEN_21977 ? _slots_28_io_uop_is_jalr : _GEN_21653 ? _slots_27_io_uop_is_jalr : _GEN_21329 ? _slots_26_io_uop_is_jalr : _GEN_21005 ? _slots_25_io_uop_is_jalr : _GEN_20681 ? _slots_24_io_uop_is_jalr : _GEN_20357 ? _slots_23_io_uop_is_jalr : _GEN_20033 ? _slots_22_io_uop_is_jalr : _GEN_19709 ? _slots_21_io_uop_is_jalr : _GEN_19385 ? _slots_20_io_uop_is_jalr : _GEN_19061 ? _slots_19_io_uop_is_jalr : _GEN_18737 ? _slots_18_io_uop_is_jalr : _GEN_18413 ? _slots_17_io_uop_is_jalr : _GEN_18089 ? _slots_16_io_uop_is_jalr : _GEN_17765 ? _slots_15_io_uop_is_jalr : _GEN_17441 ? _slots_14_io_uop_is_jalr : _GEN_17117 ? _slots_13_io_uop_is_jalr : _GEN_16793 ? _slots_12_io_uop_is_jalr : _GEN_16469 ? _slots_11_io_uop_is_jalr : _GEN_16145 ? _slots_10_io_uop_is_jalr : _GEN_15821 ? _slots_9_io_uop_is_jalr : _GEN_15497 ? _slots_8_io_uop_is_jalr : _GEN_15173 ? _slots_7_io_uop_is_jalr : _GEN_14849 ? _slots_6_io_uop_is_jalr : _GEN_14525 ? _slots_5_io_uop_is_jalr : _GEN_14201 ? _slots_4_io_uop_is_jalr : _GEN_13877 ? _slots_3_io_uop_is_jalr : _GEN_13553 ? _slots_2_io_uop_is_jalr : _GEN_13229 ? _slots_1_io_uop_is_jalr : _GEN_12906 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_0_is_jal = _GEN_25541 ? _slots_39_io_uop_is_jal : _GEN_25217 ? _slots_38_io_uop_is_jal : _GEN_24893 ? _slots_37_io_uop_is_jal : _GEN_24569 ? _slots_36_io_uop_is_jal : _GEN_24245 ? _slots_35_io_uop_is_jal : _GEN_23921 ? _slots_34_io_uop_is_jal : _GEN_23597 ? _slots_33_io_uop_is_jal : _GEN_23273 ? _slots_32_io_uop_is_jal : _GEN_22949 ? _slots_31_io_uop_is_jal : _GEN_22625 ? _slots_30_io_uop_is_jal : _GEN_22301 ? _slots_29_io_uop_is_jal : _GEN_21977 ? _slots_28_io_uop_is_jal : _GEN_21653 ? _slots_27_io_uop_is_jal : _GEN_21329 ? _slots_26_io_uop_is_jal : _GEN_21005 ? _slots_25_io_uop_is_jal : _GEN_20681 ? _slots_24_io_uop_is_jal : _GEN_20357 ? _slots_23_io_uop_is_jal : _GEN_20033 ? _slots_22_io_uop_is_jal : _GEN_19709 ? _slots_21_io_uop_is_jal : _GEN_19385 ? _slots_20_io_uop_is_jal : _GEN_19061 ? _slots_19_io_uop_is_jal : _GEN_18737 ? _slots_18_io_uop_is_jal : _GEN_18413 ? _slots_17_io_uop_is_jal : _GEN_18089 ? _slots_16_io_uop_is_jal : _GEN_17765 ? _slots_15_io_uop_is_jal : _GEN_17441 ? _slots_14_io_uop_is_jal : _GEN_17117 ? _slots_13_io_uop_is_jal : _GEN_16793 ? _slots_12_io_uop_is_jal : _GEN_16469 ? _slots_11_io_uop_is_jal : _GEN_16145 ? _slots_10_io_uop_is_jal : _GEN_15821 ? _slots_9_io_uop_is_jal : _GEN_15497 ? _slots_8_io_uop_is_jal : _GEN_15173 ? _slots_7_io_uop_is_jal : _GEN_14849 ? _slots_6_io_uop_is_jal : _GEN_14525 ? _slots_5_io_uop_is_jal : _GEN_14201 ? _slots_4_io_uop_is_jal : _GEN_13877 ? _slots_3_io_uop_is_jal : _GEN_13553 ? _slots_2_io_uop_is_jal : _GEN_13229 ? _slots_1_io_uop_is_jal : _GEN_12906 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_0_is_sfb = _GEN_25541 ? _slots_39_io_uop_is_sfb : _GEN_25217 ? _slots_38_io_uop_is_sfb : _GEN_24893 ? _slots_37_io_uop_is_sfb : _GEN_24569 ? _slots_36_io_uop_is_sfb : _GEN_24245 ? _slots_35_io_uop_is_sfb : _GEN_23921 ? _slots_34_io_uop_is_sfb : _GEN_23597 ? _slots_33_io_uop_is_sfb : _GEN_23273 ? _slots_32_io_uop_is_sfb : _GEN_22949 ? _slots_31_io_uop_is_sfb : _GEN_22625 ? _slots_30_io_uop_is_sfb : _GEN_22301 ? _slots_29_io_uop_is_sfb : _GEN_21977 ? _slots_28_io_uop_is_sfb : _GEN_21653 ? _slots_27_io_uop_is_sfb : _GEN_21329 ? _slots_26_io_uop_is_sfb : _GEN_21005 ? _slots_25_io_uop_is_sfb : _GEN_20681 ? _slots_24_io_uop_is_sfb : _GEN_20357 ? _slots_23_io_uop_is_sfb : _GEN_20033 ? _slots_22_io_uop_is_sfb : _GEN_19709 ? _slots_21_io_uop_is_sfb : _GEN_19385 ? _slots_20_io_uop_is_sfb : _GEN_19061 ? _slots_19_io_uop_is_sfb : _GEN_18737 ? _slots_18_io_uop_is_sfb : _GEN_18413 ? _slots_17_io_uop_is_sfb : _GEN_18089 ? _slots_16_io_uop_is_sfb : _GEN_17765 ? _slots_15_io_uop_is_sfb : _GEN_17441 ? _slots_14_io_uop_is_sfb : _GEN_17117 ? _slots_13_io_uop_is_sfb : _GEN_16793 ? _slots_12_io_uop_is_sfb : _GEN_16469 ? _slots_11_io_uop_is_sfb : _GEN_16145 ? _slots_10_io_uop_is_sfb : _GEN_15821 ? _slots_9_io_uop_is_sfb : _GEN_15497 ? _slots_8_io_uop_is_sfb : _GEN_15173 ? _slots_7_io_uop_is_sfb : _GEN_14849 ? _slots_6_io_uop_is_sfb : _GEN_14525 ? _slots_5_io_uop_is_sfb : _GEN_14201 ? _slots_4_io_uop_is_sfb : _GEN_13877 ? _slots_3_io_uop_is_sfb : _GEN_13553 ? _slots_2_io_uop_is_sfb : _GEN_13229 ? _slots_1_io_uop_is_sfb : _GEN_12906 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_0_br_mask = _GEN_25541 ? _slots_39_io_uop_br_mask : _GEN_25217 ? _slots_38_io_uop_br_mask : _GEN_24893 ? _slots_37_io_uop_br_mask : _GEN_24569 ? _slots_36_io_uop_br_mask : _GEN_24245 ? _slots_35_io_uop_br_mask : _GEN_23921 ? _slots_34_io_uop_br_mask : _GEN_23597 ? _slots_33_io_uop_br_mask : _GEN_23273 ? _slots_32_io_uop_br_mask : _GEN_22949 ? _slots_31_io_uop_br_mask : _GEN_22625 ? _slots_30_io_uop_br_mask : _GEN_22301 ? _slots_29_io_uop_br_mask : _GEN_21977 ? _slots_28_io_uop_br_mask : _GEN_21653 ? _slots_27_io_uop_br_mask : _GEN_21329 ? _slots_26_io_uop_br_mask : _GEN_21005 ? _slots_25_io_uop_br_mask : _GEN_20681 ? _slots_24_io_uop_br_mask : _GEN_20357 ? _slots_23_io_uop_br_mask : _GEN_20033 ? _slots_22_io_uop_br_mask : _GEN_19709 ? _slots_21_io_uop_br_mask : _GEN_19385 ? _slots_20_io_uop_br_mask : _GEN_19061 ? _slots_19_io_uop_br_mask : _GEN_18737 ? _slots_18_io_uop_br_mask : _GEN_18413 ? _slots_17_io_uop_br_mask : _GEN_18089 ? _slots_16_io_uop_br_mask : _GEN_17765 ? _slots_15_io_uop_br_mask : _GEN_17441 ? _slots_14_io_uop_br_mask : _GEN_17117 ? _slots_13_io_uop_br_mask : _GEN_16793 ? _slots_12_io_uop_br_mask : _GEN_16469 ? _slots_11_io_uop_br_mask : _GEN_16145 ? _slots_10_io_uop_br_mask : _GEN_15821 ? _slots_9_io_uop_br_mask : _GEN_15497 ? _slots_8_io_uop_br_mask : _GEN_15173 ? _slots_7_io_uop_br_mask : _GEN_14849 ? _slots_6_io_uop_br_mask : _GEN_14525 ? _slots_5_io_uop_br_mask : _GEN_14201 ? _slots_4_io_uop_br_mask : _GEN_13877 ? _slots_3_io_uop_br_mask : _GEN_13553 ? _slots_2_io_uop_br_mask : _GEN_13229 ? _slots_1_io_uop_br_mask : _GEN_12906 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_0_br_tag = _GEN_25541 ? _slots_39_io_uop_br_tag : _GEN_25217 ? _slots_38_io_uop_br_tag : _GEN_24893 ? _slots_37_io_uop_br_tag : _GEN_24569 ? _slots_36_io_uop_br_tag : _GEN_24245 ? _slots_35_io_uop_br_tag : _GEN_23921 ? _slots_34_io_uop_br_tag : _GEN_23597 ? _slots_33_io_uop_br_tag : _GEN_23273 ? _slots_32_io_uop_br_tag : _GEN_22949 ? _slots_31_io_uop_br_tag : _GEN_22625 ? _slots_30_io_uop_br_tag : _GEN_22301 ? _slots_29_io_uop_br_tag : _GEN_21977 ? _slots_28_io_uop_br_tag : _GEN_21653 ? _slots_27_io_uop_br_tag : _GEN_21329 ? _slots_26_io_uop_br_tag : _GEN_21005 ? _slots_25_io_uop_br_tag : _GEN_20681 ? _slots_24_io_uop_br_tag : _GEN_20357 ? _slots_23_io_uop_br_tag : _GEN_20033 ? _slots_22_io_uop_br_tag : _GEN_19709 ? _slots_21_io_uop_br_tag : _GEN_19385 ? _slots_20_io_uop_br_tag : _GEN_19061 ? _slots_19_io_uop_br_tag : _GEN_18737 ? _slots_18_io_uop_br_tag : _GEN_18413 ? _slots_17_io_uop_br_tag : _GEN_18089 ? _slots_16_io_uop_br_tag : _GEN_17765 ? _slots_15_io_uop_br_tag : _GEN_17441 ? _slots_14_io_uop_br_tag : _GEN_17117 ? _slots_13_io_uop_br_tag : _GEN_16793 ? _slots_12_io_uop_br_tag : _GEN_16469 ? _slots_11_io_uop_br_tag : _GEN_16145 ? _slots_10_io_uop_br_tag : _GEN_15821 ? _slots_9_io_uop_br_tag : _GEN_15497 ? _slots_8_io_uop_br_tag : _GEN_15173 ? _slots_7_io_uop_br_tag : _GEN_14849 ? _slots_6_io_uop_br_tag : _GEN_14525 ? _slots_5_io_uop_br_tag : _GEN_14201 ? _slots_4_io_uop_br_tag : _GEN_13877 ? _slots_3_io_uop_br_tag : _GEN_13553 ? _slots_2_io_uop_br_tag : _GEN_13229 ? _slots_1_io_uop_br_tag : _GEN_12906 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_0_ftq_idx = _GEN_25541 ? _slots_39_io_uop_ftq_idx : _GEN_25217 ? _slots_38_io_uop_ftq_idx : _GEN_24893 ? _slots_37_io_uop_ftq_idx : _GEN_24569 ? _slots_36_io_uop_ftq_idx : _GEN_24245 ? _slots_35_io_uop_ftq_idx : _GEN_23921 ? _slots_34_io_uop_ftq_idx : _GEN_23597 ? _slots_33_io_uop_ftq_idx : _GEN_23273 ? _slots_32_io_uop_ftq_idx : _GEN_22949 ? _slots_31_io_uop_ftq_idx : _GEN_22625 ? _slots_30_io_uop_ftq_idx : _GEN_22301 ? _slots_29_io_uop_ftq_idx : _GEN_21977 ? _slots_28_io_uop_ftq_idx : _GEN_21653 ? _slots_27_io_uop_ftq_idx : _GEN_21329 ? _slots_26_io_uop_ftq_idx : _GEN_21005 ? _slots_25_io_uop_ftq_idx : _GEN_20681 ? _slots_24_io_uop_ftq_idx : _GEN_20357 ? _slots_23_io_uop_ftq_idx : _GEN_20033 ? _slots_22_io_uop_ftq_idx : _GEN_19709 ? _slots_21_io_uop_ftq_idx : _GEN_19385 ? _slots_20_io_uop_ftq_idx : _GEN_19061 ? _slots_19_io_uop_ftq_idx : _GEN_18737 ? _slots_18_io_uop_ftq_idx : _GEN_18413 ? _slots_17_io_uop_ftq_idx : _GEN_18089 ? _slots_16_io_uop_ftq_idx : _GEN_17765 ? _slots_15_io_uop_ftq_idx : _GEN_17441 ? _slots_14_io_uop_ftq_idx : _GEN_17117 ? _slots_13_io_uop_ftq_idx : _GEN_16793 ? _slots_12_io_uop_ftq_idx : _GEN_16469 ? _slots_11_io_uop_ftq_idx : _GEN_16145 ? _slots_10_io_uop_ftq_idx : _GEN_15821 ? _slots_9_io_uop_ftq_idx : _GEN_15497 ? _slots_8_io_uop_ftq_idx : _GEN_15173 ? _slots_7_io_uop_ftq_idx : _GEN_14849 ? _slots_6_io_uop_ftq_idx : _GEN_14525 ? _slots_5_io_uop_ftq_idx : _GEN_14201 ? _slots_4_io_uop_ftq_idx : _GEN_13877 ? _slots_3_io_uop_ftq_idx : _GEN_13553 ? _slots_2_io_uop_ftq_idx : _GEN_13229 ? _slots_1_io_uop_ftq_idx : _GEN_12906 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_0_edge_inst = _GEN_25541 ? _slots_39_io_uop_edge_inst : _GEN_25217 ? _slots_38_io_uop_edge_inst : _GEN_24893 ? _slots_37_io_uop_edge_inst : _GEN_24569 ? _slots_36_io_uop_edge_inst : _GEN_24245 ? _slots_35_io_uop_edge_inst : _GEN_23921 ? _slots_34_io_uop_edge_inst : _GEN_23597 ? _slots_33_io_uop_edge_inst : _GEN_23273 ? _slots_32_io_uop_edge_inst : _GEN_22949 ? _slots_31_io_uop_edge_inst : _GEN_22625 ? _slots_30_io_uop_edge_inst : _GEN_22301 ? _slots_29_io_uop_edge_inst : _GEN_21977 ? _slots_28_io_uop_edge_inst : _GEN_21653 ? _slots_27_io_uop_edge_inst : _GEN_21329 ? _slots_26_io_uop_edge_inst : _GEN_21005 ? _slots_25_io_uop_edge_inst : _GEN_20681 ? _slots_24_io_uop_edge_inst : _GEN_20357 ? _slots_23_io_uop_edge_inst : _GEN_20033 ? _slots_22_io_uop_edge_inst : _GEN_19709 ? _slots_21_io_uop_edge_inst : _GEN_19385 ? _slots_20_io_uop_edge_inst : _GEN_19061 ? _slots_19_io_uop_edge_inst : _GEN_18737 ? _slots_18_io_uop_edge_inst : _GEN_18413 ? _slots_17_io_uop_edge_inst : _GEN_18089 ? _slots_16_io_uop_edge_inst : _GEN_17765 ? _slots_15_io_uop_edge_inst : _GEN_17441 ? _slots_14_io_uop_edge_inst : _GEN_17117 ? _slots_13_io_uop_edge_inst : _GEN_16793 ? _slots_12_io_uop_edge_inst : _GEN_16469 ? _slots_11_io_uop_edge_inst : _GEN_16145 ? _slots_10_io_uop_edge_inst : _GEN_15821 ? _slots_9_io_uop_edge_inst : _GEN_15497 ? _slots_8_io_uop_edge_inst : _GEN_15173 ? _slots_7_io_uop_edge_inst : _GEN_14849 ? _slots_6_io_uop_edge_inst : _GEN_14525 ? _slots_5_io_uop_edge_inst : _GEN_14201 ? _slots_4_io_uop_edge_inst : _GEN_13877 ? _slots_3_io_uop_edge_inst : _GEN_13553 ? _slots_2_io_uop_edge_inst : _GEN_13229 ? _slots_1_io_uop_edge_inst : _GEN_12906 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_0_pc_lob = _GEN_25541 ? _slots_39_io_uop_pc_lob : _GEN_25217 ? _slots_38_io_uop_pc_lob : _GEN_24893 ? _slots_37_io_uop_pc_lob : _GEN_24569 ? _slots_36_io_uop_pc_lob : _GEN_24245 ? _slots_35_io_uop_pc_lob : _GEN_23921 ? _slots_34_io_uop_pc_lob : _GEN_23597 ? _slots_33_io_uop_pc_lob : _GEN_23273 ? _slots_32_io_uop_pc_lob : _GEN_22949 ? _slots_31_io_uop_pc_lob : _GEN_22625 ? _slots_30_io_uop_pc_lob : _GEN_22301 ? _slots_29_io_uop_pc_lob : _GEN_21977 ? _slots_28_io_uop_pc_lob : _GEN_21653 ? _slots_27_io_uop_pc_lob : _GEN_21329 ? _slots_26_io_uop_pc_lob : _GEN_21005 ? _slots_25_io_uop_pc_lob : _GEN_20681 ? _slots_24_io_uop_pc_lob : _GEN_20357 ? _slots_23_io_uop_pc_lob : _GEN_20033 ? _slots_22_io_uop_pc_lob : _GEN_19709 ? _slots_21_io_uop_pc_lob : _GEN_19385 ? _slots_20_io_uop_pc_lob : _GEN_19061 ? _slots_19_io_uop_pc_lob : _GEN_18737 ? _slots_18_io_uop_pc_lob : _GEN_18413 ? _slots_17_io_uop_pc_lob : _GEN_18089 ? _slots_16_io_uop_pc_lob : _GEN_17765 ? _slots_15_io_uop_pc_lob : _GEN_17441 ? _slots_14_io_uop_pc_lob : _GEN_17117 ? _slots_13_io_uop_pc_lob : _GEN_16793 ? _slots_12_io_uop_pc_lob : _GEN_16469 ? _slots_11_io_uop_pc_lob : _GEN_16145 ? _slots_10_io_uop_pc_lob : _GEN_15821 ? _slots_9_io_uop_pc_lob : _GEN_15497 ? _slots_8_io_uop_pc_lob : _GEN_15173 ? _slots_7_io_uop_pc_lob : _GEN_14849 ? _slots_6_io_uop_pc_lob : _GEN_14525 ? _slots_5_io_uop_pc_lob : _GEN_14201 ? _slots_4_io_uop_pc_lob : _GEN_13877 ? _slots_3_io_uop_pc_lob : _GEN_13553 ? _slots_2_io_uop_pc_lob : _GEN_13229 ? _slots_1_io_uop_pc_lob : _GEN_12906 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_0_taken = _GEN_25541 ? _slots_39_io_uop_taken : _GEN_25217 ? _slots_38_io_uop_taken : _GEN_24893 ? _slots_37_io_uop_taken : _GEN_24569 ? _slots_36_io_uop_taken : _GEN_24245 ? _slots_35_io_uop_taken : _GEN_23921 ? _slots_34_io_uop_taken : _GEN_23597 ? _slots_33_io_uop_taken : _GEN_23273 ? _slots_32_io_uop_taken : _GEN_22949 ? _slots_31_io_uop_taken : _GEN_22625 ? _slots_30_io_uop_taken : _GEN_22301 ? _slots_29_io_uop_taken : _GEN_21977 ? _slots_28_io_uop_taken : _GEN_21653 ? _slots_27_io_uop_taken : _GEN_21329 ? _slots_26_io_uop_taken : _GEN_21005 ? _slots_25_io_uop_taken : _GEN_20681 ? _slots_24_io_uop_taken : _GEN_20357 ? _slots_23_io_uop_taken : _GEN_20033 ? _slots_22_io_uop_taken : _GEN_19709 ? _slots_21_io_uop_taken : _GEN_19385 ? _slots_20_io_uop_taken : _GEN_19061 ? _slots_19_io_uop_taken : _GEN_18737 ? _slots_18_io_uop_taken : _GEN_18413 ? _slots_17_io_uop_taken : _GEN_18089 ? _slots_16_io_uop_taken : _GEN_17765 ? _slots_15_io_uop_taken : _GEN_17441 ? _slots_14_io_uop_taken : _GEN_17117 ? _slots_13_io_uop_taken : _GEN_16793 ? _slots_12_io_uop_taken : _GEN_16469 ? _slots_11_io_uop_taken : _GEN_16145 ? _slots_10_io_uop_taken : _GEN_15821 ? _slots_9_io_uop_taken : _GEN_15497 ? _slots_8_io_uop_taken : _GEN_15173 ? _slots_7_io_uop_taken : _GEN_14849 ? _slots_6_io_uop_taken : _GEN_14525 ? _slots_5_io_uop_taken : _GEN_14201 ? _slots_4_io_uop_taken : _GEN_13877 ? _slots_3_io_uop_taken : _GEN_13553 ? _slots_2_io_uop_taken : _GEN_13229 ? _slots_1_io_uop_taken : _GEN_12906 & _slots_0_io_uop_taken;
  assign io_iss_uops_0_imm_packed = _GEN_25541 ? _slots_39_io_uop_imm_packed : _GEN_25217 ? _slots_38_io_uop_imm_packed : _GEN_24893 ? _slots_37_io_uop_imm_packed : _GEN_24569 ? _slots_36_io_uop_imm_packed : _GEN_24245 ? _slots_35_io_uop_imm_packed : _GEN_23921 ? _slots_34_io_uop_imm_packed : _GEN_23597 ? _slots_33_io_uop_imm_packed : _GEN_23273 ? _slots_32_io_uop_imm_packed : _GEN_22949 ? _slots_31_io_uop_imm_packed : _GEN_22625 ? _slots_30_io_uop_imm_packed : _GEN_22301 ? _slots_29_io_uop_imm_packed : _GEN_21977 ? _slots_28_io_uop_imm_packed : _GEN_21653 ? _slots_27_io_uop_imm_packed : _GEN_21329 ? _slots_26_io_uop_imm_packed : _GEN_21005 ? _slots_25_io_uop_imm_packed : _GEN_20681 ? _slots_24_io_uop_imm_packed : _GEN_20357 ? _slots_23_io_uop_imm_packed : _GEN_20033 ? _slots_22_io_uop_imm_packed : _GEN_19709 ? _slots_21_io_uop_imm_packed : _GEN_19385 ? _slots_20_io_uop_imm_packed : _GEN_19061 ? _slots_19_io_uop_imm_packed : _GEN_18737 ? _slots_18_io_uop_imm_packed : _GEN_18413 ? _slots_17_io_uop_imm_packed : _GEN_18089 ? _slots_16_io_uop_imm_packed : _GEN_17765 ? _slots_15_io_uop_imm_packed : _GEN_17441 ? _slots_14_io_uop_imm_packed : _GEN_17117 ? _slots_13_io_uop_imm_packed : _GEN_16793 ? _slots_12_io_uop_imm_packed : _GEN_16469 ? _slots_11_io_uop_imm_packed : _GEN_16145 ? _slots_10_io_uop_imm_packed : _GEN_15821 ? _slots_9_io_uop_imm_packed : _GEN_15497 ? _slots_8_io_uop_imm_packed : _GEN_15173 ? _slots_7_io_uop_imm_packed : _GEN_14849 ? _slots_6_io_uop_imm_packed : _GEN_14525 ? _slots_5_io_uop_imm_packed : _GEN_14201 ? _slots_4_io_uop_imm_packed : _GEN_13877 ? _slots_3_io_uop_imm_packed : _GEN_13553 ? _slots_2_io_uop_imm_packed : _GEN_13229 ? _slots_1_io_uop_imm_packed : _GEN_12906 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_0_rob_idx = _GEN_25541 ? _slots_39_io_uop_rob_idx : _GEN_25217 ? _slots_38_io_uop_rob_idx : _GEN_24893 ? _slots_37_io_uop_rob_idx : _GEN_24569 ? _slots_36_io_uop_rob_idx : _GEN_24245 ? _slots_35_io_uop_rob_idx : _GEN_23921 ? _slots_34_io_uop_rob_idx : _GEN_23597 ? _slots_33_io_uop_rob_idx : _GEN_23273 ? _slots_32_io_uop_rob_idx : _GEN_22949 ? _slots_31_io_uop_rob_idx : _GEN_22625 ? _slots_30_io_uop_rob_idx : _GEN_22301 ? _slots_29_io_uop_rob_idx : _GEN_21977 ? _slots_28_io_uop_rob_idx : _GEN_21653 ? _slots_27_io_uop_rob_idx : _GEN_21329 ? _slots_26_io_uop_rob_idx : _GEN_21005 ? _slots_25_io_uop_rob_idx : _GEN_20681 ? _slots_24_io_uop_rob_idx : _GEN_20357 ? _slots_23_io_uop_rob_idx : _GEN_20033 ? _slots_22_io_uop_rob_idx : _GEN_19709 ? _slots_21_io_uop_rob_idx : _GEN_19385 ? _slots_20_io_uop_rob_idx : _GEN_19061 ? _slots_19_io_uop_rob_idx : _GEN_18737 ? _slots_18_io_uop_rob_idx : _GEN_18413 ? _slots_17_io_uop_rob_idx : _GEN_18089 ? _slots_16_io_uop_rob_idx : _GEN_17765 ? _slots_15_io_uop_rob_idx : _GEN_17441 ? _slots_14_io_uop_rob_idx : _GEN_17117 ? _slots_13_io_uop_rob_idx : _GEN_16793 ? _slots_12_io_uop_rob_idx : _GEN_16469 ? _slots_11_io_uop_rob_idx : _GEN_16145 ? _slots_10_io_uop_rob_idx : _GEN_15821 ? _slots_9_io_uop_rob_idx : _GEN_15497 ? _slots_8_io_uop_rob_idx : _GEN_15173 ? _slots_7_io_uop_rob_idx : _GEN_14849 ? _slots_6_io_uop_rob_idx : _GEN_14525 ? _slots_5_io_uop_rob_idx : _GEN_14201 ? _slots_4_io_uop_rob_idx : _GEN_13877 ? _slots_3_io_uop_rob_idx : _GEN_13553 ? _slots_2_io_uop_rob_idx : _GEN_13229 ? _slots_1_io_uop_rob_idx : _GEN_12906 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_0_ldq_idx = _GEN_25541 ? _slots_39_io_uop_ldq_idx : _GEN_25217 ? _slots_38_io_uop_ldq_idx : _GEN_24893 ? _slots_37_io_uop_ldq_idx : _GEN_24569 ? _slots_36_io_uop_ldq_idx : _GEN_24245 ? _slots_35_io_uop_ldq_idx : _GEN_23921 ? _slots_34_io_uop_ldq_idx : _GEN_23597 ? _slots_33_io_uop_ldq_idx : _GEN_23273 ? _slots_32_io_uop_ldq_idx : _GEN_22949 ? _slots_31_io_uop_ldq_idx : _GEN_22625 ? _slots_30_io_uop_ldq_idx : _GEN_22301 ? _slots_29_io_uop_ldq_idx : _GEN_21977 ? _slots_28_io_uop_ldq_idx : _GEN_21653 ? _slots_27_io_uop_ldq_idx : _GEN_21329 ? _slots_26_io_uop_ldq_idx : _GEN_21005 ? _slots_25_io_uop_ldq_idx : _GEN_20681 ? _slots_24_io_uop_ldq_idx : _GEN_20357 ? _slots_23_io_uop_ldq_idx : _GEN_20033 ? _slots_22_io_uop_ldq_idx : _GEN_19709 ? _slots_21_io_uop_ldq_idx : _GEN_19385 ? _slots_20_io_uop_ldq_idx : _GEN_19061 ? _slots_19_io_uop_ldq_idx : _GEN_18737 ? _slots_18_io_uop_ldq_idx : _GEN_18413 ? _slots_17_io_uop_ldq_idx : _GEN_18089 ? _slots_16_io_uop_ldq_idx : _GEN_17765 ? _slots_15_io_uop_ldq_idx : _GEN_17441 ? _slots_14_io_uop_ldq_idx : _GEN_17117 ? _slots_13_io_uop_ldq_idx : _GEN_16793 ? _slots_12_io_uop_ldq_idx : _GEN_16469 ? _slots_11_io_uop_ldq_idx : _GEN_16145 ? _slots_10_io_uop_ldq_idx : _GEN_15821 ? _slots_9_io_uop_ldq_idx : _GEN_15497 ? _slots_8_io_uop_ldq_idx : _GEN_15173 ? _slots_7_io_uop_ldq_idx : _GEN_14849 ? _slots_6_io_uop_ldq_idx : _GEN_14525 ? _slots_5_io_uop_ldq_idx : _GEN_14201 ? _slots_4_io_uop_ldq_idx : _GEN_13877 ? _slots_3_io_uop_ldq_idx : _GEN_13553 ? _slots_2_io_uop_ldq_idx : _GEN_13229 ? _slots_1_io_uop_ldq_idx : _GEN_12906 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_0_stq_idx = _GEN_25541 ? _slots_39_io_uop_stq_idx : _GEN_25217 ? _slots_38_io_uop_stq_idx : _GEN_24893 ? _slots_37_io_uop_stq_idx : _GEN_24569 ? _slots_36_io_uop_stq_idx : _GEN_24245 ? _slots_35_io_uop_stq_idx : _GEN_23921 ? _slots_34_io_uop_stq_idx : _GEN_23597 ? _slots_33_io_uop_stq_idx : _GEN_23273 ? _slots_32_io_uop_stq_idx : _GEN_22949 ? _slots_31_io_uop_stq_idx : _GEN_22625 ? _slots_30_io_uop_stq_idx : _GEN_22301 ? _slots_29_io_uop_stq_idx : _GEN_21977 ? _slots_28_io_uop_stq_idx : _GEN_21653 ? _slots_27_io_uop_stq_idx : _GEN_21329 ? _slots_26_io_uop_stq_idx : _GEN_21005 ? _slots_25_io_uop_stq_idx : _GEN_20681 ? _slots_24_io_uop_stq_idx : _GEN_20357 ? _slots_23_io_uop_stq_idx : _GEN_20033 ? _slots_22_io_uop_stq_idx : _GEN_19709 ? _slots_21_io_uop_stq_idx : _GEN_19385 ? _slots_20_io_uop_stq_idx : _GEN_19061 ? _slots_19_io_uop_stq_idx : _GEN_18737 ? _slots_18_io_uop_stq_idx : _GEN_18413 ? _slots_17_io_uop_stq_idx : _GEN_18089 ? _slots_16_io_uop_stq_idx : _GEN_17765 ? _slots_15_io_uop_stq_idx : _GEN_17441 ? _slots_14_io_uop_stq_idx : _GEN_17117 ? _slots_13_io_uop_stq_idx : _GEN_16793 ? _slots_12_io_uop_stq_idx : _GEN_16469 ? _slots_11_io_uop_stq_idx : _GEN_16145 ? _slots_10_io_uop_stq_idx : _GEN_15821 ? _slots_9_io_uop_stq_idx : _GEN_15497 ? _slots_8_io_uop_stq_idx : _GEN_15173 ? _slots_7_io_uop_stq_idx : _GEN_14849 ? _slots_6_io_uop_stq_idx : _GEN_14525 ? _slots_5_io_uop_stq_idx : _GEN_14201 ? _slots_4_io_uop_stq_idx : _GEN_13877 ? _slots_3_io_uop_stq_idx : _GEN_13553 ? _slots_2_io_uop_stq_idx : _GEN_13229 ? _slots_1_io_uop_stq_idx : _GEN_12906 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_0_pdst = _GEN_25541 ? _slots_39_io_uop_pdst : _GEN_25217 ? _slots_38_io_uop_pdst : _GEN_24893 ? _slots_37_io_uop_pdst : _GEN_24569 ? _slots_36_io_uop_pdst : _GEN_24245 ? _slots_35_io_uop_pdst : _GEN_23921 ? _slots_34_io_uop_pdst : _GEN_23597 ? _slots_33_io_uop_pdst : _GEN_23273 ? _slots_32_io_uop_pdst : _GEN_22949 ? _slots_31_io_uop_pdst : _GEN_22625 ? _slots_30_io_uop_pdst : _GEN_22301 ? _slots_29_io_uop_pdst : _GEN_21977 ? _slots_28_io_uop_pdst : _GEN_21653 ? _slots_27_io_uop_pdst : _GEN_21329 ? _slots_26_io_uop_pdst : _GEN_21005 ? _slots_25_io_uop_pdst : _GEN_20681 ? _slots_24_io_uop_pdst : _GEN_20357 ? _slots_23_io_uop_pdst : _GEN_20033 ? _slots_22_io_uop_pdst : _GEN_19709 ? _slots_21_io_uop_pdst : _GEN_19385 ? _slots_20_io_uop_pdst : _GEN_19061 ? _slots_19_io_uop_pdst : _GEN_18737 ? _slots_18_io_uop_pdst : _GEN_18413 ? _slots_17_io_uop_pdst : _GEN_18089 ? _slots_16_io_uop_pdst : _GEN_17765 ? _slots_15_io_uop_pdst : _GEN_17441 ? _slots_14_io_uop_pdst : _GEN_17117 ? _slots_13_io_uop_pdst : _GEN_16793 ? _slots_12_io_uop_pdst : _GEN_16469 ? _slots_11_io_uop_pdst : _GEN_16145 ? _slots_10_io_uop_pdst : _GEN_15821 ? _slots_9_io_uop_pdst : _GEN_15497 ? _slots_8_io_uop_pdst : _GEN_15173 ? _slots_7_io_uop_pdst : _GEN_14849 ? _slots_6_io_uop_pdst : _GEN_14525 ? _slots_5_io_uop_pdst : _GEN_14201 ? _slots_4_io_uop_pdst : _GEN_13877 ? _slots_3_io_uop_pdst : _GEN_13553 ? _slots_2_io_uop_pdst : _GEN_13229 ? _slots_1_io_uop_pdst : _GEN_12906 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_0_prs1 = _GEN_25541 ? _slots_39_io_uop_prs1 : _GEN_25217 ? _slots_38_io_uop_prs1 : _GEN_24893 ? _slots_37_io_uop_prs1 : _GEN_24569 ? _slots_36_io_uop_prs1 : _GEN_24245 ? _slots_35_io_uop_prs1 : _GEN_23921 ? _slots_34_io_uop_prs1 : _GEN_23597 ? _slots_33_io_uop_prs1 : _GEN_23273 ? _slots_32_io_uop_prs1 : _GEN_22949 ? _slots_31_io_uop_prs1 : _GEN_22625 ? _slots_30_io_uop_prs1 : _GEN_22301 ? _slots_29_io_uop_prs1 : _GEN_21977 ? _slots_28_io_uop_prs1 : _GEN_21653 ? _slots_27_io_uop_prs1 : _GEN_21329 ? _slots_26_io_uop_prs1 : _GEN_21005 ? _slots_25_io_uop_prs1 : _GEN_20681 ? _slots_24_io_uop_prs1 : _GEN_20357 ? _slots_23_io_uop_prs1 : _GEN_20033 ? _slots_22_io_uop_prs1 : _GEN_19709 ? _slots_21_io_uop_prs1 : _GEN_19385 ? _slots_20_io_uop_prs1 : _GEN_19061 ? _slots_19_io_uop_prs1 : _GEN_18737 ? _slots_18_io_uop_prs1 : _GEN_18413 ? _slots_17_io_uop_prs1 : _GEN_18089 ? _slots_16_io_uop_prs1 : _GEN_17765 ? _slots_15_io_uop_prs1 : _GEN_17441 ? _slots_14_io_uop_prs1 : _GEN_17117 ? _slots_13_io_uop_prs1 : _GEN_16793 ? _slots_12_io_uop_prs1 : _GEN_16469 ? _slots_11_io_uop_prs1 : _GEN_16145 ? _slots_10_io_uop_prs1 : _GEN_15821 ? _slots_9_io_uop_prs1 : _GEN_15497 ? _slots_8_io_uop_prs1 : _GEN_15173 ? _slots_7_io_uop_prs1 : _GEN_14849 ? _slots_6_io_uop_prs1 : _GEN_14525 ? _slots_5_io_uop_prs1 : _GEN_14201 ? _slots_4_io_uop_prs1 : _GEN_13877 ? _slots_3_io_uop_prs1 : _GEN_13553 ? _slots_2_io_uop_prs1 : _GEN_13229 ? _slots_1_io_uop_prs1 : _GEN_12906 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_0_prs2 = _GEN_25541 ? _slots_39_io_uop_prs2 : _GEN_25217 ? _slots_38_io_uop_prs2 : _GEN_24893 ? _slots_37_io_uop_prs2 : _GEN_24569 ? _slots_36_io_uop_prs2 : _GEN_24245 ? _slots_35_io_uop_prs2 : _GEN_23921 ? _slots_34_io_uop_prs2 : _GEN_23597 ? _slots_33_io_uop_prs2 : _GEN_23273 ? _slots_32_io_uop_prs2 : _GEN_22949 ? _slots_31_io_uop_prs2 : _GEN_22625 ? _slots_30_io_uop_prs2 : _GEN_22301 ? _slots_29_io_uop_prs2 : _GEN_21977 ? _slots_28_io_uop_prs2 : _GEN_21653 ? _slots_27_io_uop_prs2 : _GEN_21329 ? _slots_26_io_uop_prs2 : _GEN_21005 ? _slots_25_io_uop_prs2 : _GEN_20681 ? _slots_24_io_uop_prs2 : _GEN_20357 ? _slots_23_io_uop_prs2 : _GEN_20033 ? _slots_22_io_uop_prs2 : _GEN_19709 ? _slots_21_io_uop_prs2 : _GEN_19385 ? _slots_20_io_uop_prs2 : _GEN_19061 ? _slots_19_io_uop_prs2 : _GEN_18737 ? _slots_18_io_uop_prs2 : _GEN_18413 ? _slots_17_io_uop_prs2 : _GEN_18089 ? _slots_16_io_uop_prs2 : _GEN_17765 ? _slots_15_io_uop_prs2 : _GEN_17441 ? _slots_14_io_uop_prs2 : _GEN_17117 ? _slots_13_io_uop_prs2 : _GEN_16793 ? _slots_12_io_uop_prs2 : _GEN_16469 ? _slots_11_io_uop_prs2 : _GEN_16145 ? _slots_10_io_uop_prs2 : _GEN_15821 ? _slots_9_io_uop_prs2 : _GEN_15497 ? _slots_8_io_uop_prs2 : _GEN_15173 ? _slots_7_io_uop_prs2 : _GEN_14849 ? _slots_6_io_uop_prs2 : _GEN_14525 ? _slots_5_io_uop_prs2 : _GEN_14201 ? _slots_4_io_uop_prs2 : _GEN_13877 ? _slots_3_io_uop_prs2 : _GEN_13553 ? _slots_2_io_uop_prs2 : _GEN_13229 ? _slots_1_io_uop_prs2 : _GEN_12906 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_0_bypassable = _GEN_25541 ? _slots_39_io_uop_bypassable : _GEN_25217 ? _slots_38_io_uop_bypassable : _GEN_24893 ? _slots_37_io_uop_bypassable : _GEN_24569 ? _slots_36_io_uop_bypassable : _GEN_24245 ? _slots_35_io_uop_bypassable : _GEN_23921 ? _slots_34_io_uop_bypassable : _GEN_23597 ? _slots_33_io_uop_bypassable : _GEN_23273 ? _slots_32_io_uop_bypassable : _GEN_22949 ? _slots_31_io_uop_bypassable : _GEN_22625 ? _slots_30_io_uop_bypassable : _GEN_22301 ? _slots_29_io_uop_bypassable : _GEN_21977 ? _slots_28_io_uop_bypassable : _GEN_21653 ? _slots_27_io_uop_bypassable : _GEN_21329 ? _slots_26_io_uop_bypassable : _GEN_21005 ? _slots_25_io_uop_bypassable : _GEN_20681 ? _slots_24_io_uop_bypassable : _GEN_20357 ? _slots_23_io_uop_bypassable : _GEN_20033 ? _slots_22_io_uop_bypassable : _GEN_19709 ? _slots_21_io_uop_bypassable : _GEN_19385 ? _slots_20_io_uop_bypassable : _GEN_19061 ? _slots_19_io_uop_bypassable : _GEN_18737 ? _slots_18_io_uop_bypassable : _GEN_18413 ? _slots_17_io_uop_bypassable : _GEN_18089 ? _slots_16_io_uop_bypassable : _GEN_17765 ? _slots_15_io_uop_bypassable : _GEN_17441 ? _slots_14_io_uop_bypassable : _GEN_17117 ? _slots_13_io_uop_bypassable : _GEN_16793 ? _slots_12_io_uop_bypassable : _GEN_16469 ? _slots_11_io_uop_bypassable : _GEN_16145 ? _slots_10_io_uop_bypassable : _GEN_15821 ? _slots_9_io_uop_bypassable : _GEN_15497 ? _slots_8_io_uop_bypassable : _GEN_15173 ? _slots_7_io_uop_bypassable : _GEN_14849 ? _slots_6_io_uop_bypassable : _GEN_14525 ? _slots_5_io_uop_bypassable : _GEN_14201 ? _slots_4_io_uop_bypassable : _GEN_13877 ? _slots_3_io_uop_bypassable : _GEN_13553 ? _slots_2_io_uop_bypassable : _GEN_13229 ? _slots_1_io_uop_bypassable : _GEN_12906 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_0_mem_cmd = _GEN_25541 ? _slots_39_io_uop_mem_cmd : _GEN_25217 ? _slots_38_io_uop_mem_cmd : _GEN_24893 ? _slots_37_io_uop_mem_cmd : _GEN_24569 ? _slots_36_io_uop_mem_cmd : _GEN_24245 ? _slots_35_io_uop_mem_cmd : _GEN_23921 ? _slots_34_io_uop_mem_cmd : _GEN_23597 ? _slots_33_io_uop_mem_cmd : _GEN_23273 ? _slots_32_io_uop_mem_cmd : _GEN_22949 ? _slots_31_io_uop_mem_cmd : _GEN_22625 ? _slots_30_io_uop_mem_cmd : _GEN_22301 ? _slots_29_io_uop_mem_cmd : _GEN_21977 ? _slots_28_io_uop_mem_cmd : _GEN_21653 ? _slots_27_io_uop_mem_cmd : _GEN_21329 ? _slots_26_io_uop_mem_cmd : _GEN_21005 ? _slots_25_io_uop_mem_cmd : _GEN_20681 ? _slots_24_io_uop_mem_cmd : _GEN_20357 ? _slots_23_io_uop_mem_cmd : _GEN_20033 ? _slots_22_io_uop_mem_cmd : _GEN_19709 ? _slots_21_io_uop_mem_cmd : _GEN_19385 ? _slots_20_io_uop_mem_cmd : _GEN_19061 ? _slots_19_io_uop_mem_cmd : _GEN_18737 ? _slots_18_io_uop_mem_cmd : _GEN_18413 ? _slots_17_io_uop_mem_cmd : _GEN_18089 ? _slots_16_io_uop_mem_cmd : _GEN_17765 ? _slots_15_io_uop_mem_cmd : _GEN_17441 ? _slots_14_io_uop_mem_cmd : _GEN_17117 ? _slots_13_io_uop_mem_cmd : _GEN_16793 ? _slots_12_io_uop_mem_cmd : _GEN_16469 ? _slots_11_io_uop_mem_cmd : _GEN_16145 ? _slots_10_io_uop_mem_cmd : _GEN_15821 ? _slots_9_io_uop_mem_cmd : _GEN_15497 ? _slots_8_io_uop_mem_cmd : _GEN_15173 ? _slots_7_io_uop_mem_cmd : _GEN_14849 ? _slots_6_io_uop_mem_cmd : _GEN_14525 ? _slots_5_io_uop_mem_cmd : _GEN_14201 ? _slots_4_io_uop_mem_cmd : _GEN_13877 ? _slots_3_io_uop_mem_cmd : _GEN_13553 ? _slots_2_io_uop_mem_cmd : _GEN_13229 ? _slots_1_io_uop_mem_cmd : _GEN_12906 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_0_is_amo = _GEN_25541 ? _slots_39_io_uop_is_amo : _GEN_25217 ? _slots_38_io_uop_is_amo : _GEN_24893 ? _slots_37_io_uop_is_amo : _GEN_24569 ? _slots_36_io_uop_is_amo : _GEN_24245 ? _slots_35_io_uop_is_amo : _GEN_23921 ? _slots_34_io_uop_is_amo : _GEN_23597 ? _slots_33_io_uop_is_amo : _GEN_23273 ? _slots_32_io_uop_is_amo : _GEN_22949 ? _slots_31_io_uop_is_amo : _GEN_22625 ? _slots_30_io_uop_is_amo : _GEN_22301 ? _slots_29_io_uop_is_amo : _GEN_21977 ? _slots_28_io_uop_is_amo : _GEN_21653 ? _slots_27_io_uop_is_amo : _GEN_21329 ? _slots_26_io_uop_is_amo : _GEN_21005 ? _slots_25_io_uop_is_amo : _GEN_20681 ? _slots_24_io_uop_is_amo : _GEN_20357 ? _slots_23_io_uop_is_amo : _GEN_20033 ? _slots_22_io_uop_is_amo : _GEN_19709 ? _slots_21_io_uop_is_amo : _GEN_19385 ? _slots_20_io_uop_is_amo : _GEN_19061 ? _slots_19_io_uop_is_amo : _GEN_18737 ? _slots_18_io_uop_is_amo : _GEN_18413 ? _slots_17_io_uop_is_amo : _GEN_18089 ? _slots_16_io_uop_is_amo : _GEN_17765 ? _slots_15_io_uop_is_amo : _GEN_17441 ? _slots_14_io_uop_is_amo : _GEN_17117 ? _slots_13_io_uop_is_amo : _GEN_16793 ? _slots_12_io_uop_is_amo : _GEN_16469 ? _slots_11_io_uop_is_amo : _GEN_16145 ? _slots_10_io_uop_is_amo : _GEN_15821 ? _slots_9_io_uop_is_amo : _GEN_15497 ? _slots_8_io_uop_is_amo : _GEN_15173 ? _slots_7_io_uop_is_amo : _GEN_14849 ? _slots_6_io_uop_is_amo : _GEN_14525 ? _slots_5_io_uop_is_amo : _GEN_14201 ? _slots_4_io_uop_is_amo : _GEN_13877 ? _slots_3_io_uop_is_amo : _GEN_13553 ? _slots_2_io_uop_is_amo : _GEN_13229 ? _slots_1_io_uop_is_amo : _GEN_12906 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_0_uses_stq = _GEN_25541 ? _slots_39_io_uop_uses_stq : _GEN_25217 ? _slots_38_io_uop_uses_stq : _GEN_24893 ? _slots_37_io_uop_uses_stq : _GEN_24569 ? _slots_36_io_uop_uses_stq : _GEN_24245 ? _slots_35_io_uop_uses_stq : _GEN_23921 ? _slots_34_io_uop_uses_stq : _GEN_23597 ? _slots_33_io_uop_uses_stq : _GEN_23273 ? _slots_32_io_uop_uses_stq : _GEN_22949 ? _slots_31_io_uop_uses_stq : _GEN_22625 ? _slots_30_io_uop_uses_stq : _GEN_22301 ? _slots_29_io_uop_uses_stq : _GEN_21977 ? _slots_28_io_uop_uses_stq : _GEN_21653 ? _slots_27_io_uop_uses_stq : _GEN_21329 ? _slots_26_io_uop_uses_stq : _GEN_21005 ? _slots_25_io_uop_uses_stq : _GEN_20681 ? _slots_24_io_uop_uses_stq : _GEN_20357 ? _slots_23_io_uop_uses_stq : _GEN_20033 ? _slots_22_io_uop_uses_stq : _GEN_19709 ? _slots_21_io_uop_uses_stq : _GEN_19385 ? _slots_20_io_uop_uses_stq : _GEN_19061 ? _slots_19_io_uop_uses_stq : _GEN_18737 ? _slots_18_io_uop_uses_stq : _GEN_18413 ? _slots_17_io_uop_uses_stq : _GEN_18089 ? _slots_16_io_uop_uses_stq : _GEN_17765 ? _slots_15_io_uop_uses_stq : _GEN_17441 ? _slots_14_io_uop_uses_stq : _GEN_17117 ? _slots_13_io_uop_uses_stq : _GEN_16793 ? _slots_12_io_uop_uses_stq : _GEN_16469 ? _slots_11_io_uop_uses_stq : _GEN_16145 ? _slots_10_io_uop_uses_stq : _GEN_15821 ? _slots_9_io_uop_uses_stq : _GEN_15497 ? _slots_8_io_uop_uses_stq : _GEN_15173 ? _slots_7_io_uop_uses_stq : _GEN_14849 ? _slots_6_io_uop_uses_stq : _GEN_14525 ? _slots_5_io_uop_uses_stq : _GEN_14201 ? _slots_4_io_uop_uses_stq : _GEN_13877 ? _slots_3_io_uop_uses_stq : _GEN_13553 ? _slots_2_io_uop_uses_stq : _GEN_13229 ? _slots_1_io_uop_uses_stq : _GEN_12906 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_0_ldst_val = _GEN_25541 ? _slots_39_io_uop_ldst_val : _GEN_25217 ? _slots_38_io_uop_ldst_val : _GEN_24893 ? _slots_37_io_uop_ldst_val : _GEN_24569 ? _slots_36_io_uop_ldst_val : _GEN_24245 ? _slots_35_io_uop_ldst_val : _GEN_23921 ? _slots_34_io_uop_ldst_val : _GEN_23597 ? _slots_33_io_uop_ldst_val : _GEN_23273 ? _slots_32_io_uop_ldst_val : _GEN_22949 ? _slots_31_io_uop_ldst_val : _GEN_22625 ? _slots_30_io_uop_ldst_val : _GEN_22301 ? _slots_29_io_uop_ldst_val : _GEN_21977 ? _slots_28_io_uop_ldst_val : _GEN_21653 ? _slots_27_io_uop_ldst_val : _GEN_21329 ? _slots_26_io_uop_ldst_val : _GEN_21005 ? _slots_25_io_uop_ldst_val : _GEN_20681 ? _slots_24_io_uop_ldst_val : _GEN_20357 ? _slots_23_io_uop_ldst_val : _GEN_20033 ? _slots_22_io_uop_ldst_val : _GEN_19709 ? _slots_21_io_uop_ldst_val : _GEN_19385 ? _slots_20_io_uop_ldst_val : _GEN_19061 ? _slots_19_io_uop_ldst_val : _GEN_18737 ? _slots_18_io_uop_ldst_val : _GEN_18413 ? _slots_17_io_uop_ldst_val : _GEN_18089 ? _slots_16_io_uop_ldst_val : _GEN_17765 ? _slots_15_io_uop_ldst_val : _GEN_17441 ? _slots_14_io_uop_ldst_val : _GEN_17117 ? _slots_13_io_uop_ldst_val : _GEN_16793 ? _slots_12_io_uop_ldst_val : _GEN_16469 ? _slots_11_io_uop_ldst_val : _GEN_16145 ? _slots_10_io_uop_ldst_val : _GEN_15821 ? _slots_9_io_uop_ldst_val : _GEN_15497 ? _slots_8_io_uop_ldst_val : _GEN_15173 ? _slots_7_io_uop_ldst_val : _GEN_14849 ? _slots_6_io_uop_ldst_val : _GEN_14525 ? _slots_5_io_uop_ldst_val : _GEN_14201 ? _slots_4_io_uop_ldst_val : _GEN_13877 ? _slots_3_io_uop_ldst_val : _GEN_13553 ? _slots_2_io_uop_ldst_val : _GEN_13229 ? _slots_1_io_uop_ldst_val : _GEN_12906 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_0_dst_rtype = _GEN_25541 ? _slots_39_io_uop_dst_rtype : _GEN_25217 ? _slots_38_io_uop_dst_rtype : _GEN_24893 ? _slots_37_io_uop_dst_rtype : _GEN_24569 ? _slots_36_io_uop_dst_rtype : _GEN_24245 ? _slots_35_io_uop_dst_rtype : _GEN_23921 ? _slots_34_io_uop_dst_rtype : _GEN_23597 ? _slots_33_io_uop_dst_rtype : _GEN_23273 ? _slots_32_io_uop_dst_rtype : _GEN_22949 ? _slots_31_io_uop_dst_rtype : _GEN_22625 ? _slots_30_io_uop_dst_rtype : _GEN_22301 ? _slots_29_io_uop_dst_rtype : _GEN_21977 ? _slots_28_io_uop_dst_rtype : _GEN_21653 ? _slots_27_io_uop_dst_rtype : _GEN_21329 ? _slots_26_io_uop_dst_rtype : _GEN_21005 ? _slots_25_io_uop_dst_rtype : _GEN_20681 ? _slots_24_io_uop_dst_rtype : _GEN_20357 ? _slots_23_io_uop_dst_rtype : _GEN_20033 ? _slots_22_io_uop_dst_rtype : _GEN_19709 ? _slots_21_io_uop_dst_rtype : _GEN_19385 ? _slots_20_io_uop_dst_rtype : _GEN_19061 ? _slots_19_io_uop_dst_rtype : _GEN_18737 ? _slots_18_io_uop_dst_rtype : _GEN_18413 ? _slots_17_io_uop_dst_rtype : _GEN_18089 ? _slots_16_io_uop_dst_rtype : _GEN_17765 ? _slots_15_io_uop_dst_rtype : _GEN_17441 ? _slots_14_io_uop_dst_rtype : _GEN_17117 ? _slots_13_io_uop_dst_rtype : _GEN_16793 ? _slots_12_io_uop_dst_rtype : _GEN_16469 ? _slots_11_io_uop_dst_rtype : _GEN_16145 ? _slots_10_io_uop_dst_rtype : _GEN_15821 ? _slots_9_io_uop_dst_rtype : _GEN_15497 ? _slots_8_io_uop_dst_rtype : _GEN_15173 ? _slots_7_io_uop_dst_rtype : _GEN_14849 ? _slots_6_io_uop_dst_rtype : _GEN_14525 ? _slots_5_io_uop_dst_rtype : _GEN_14201 ? _slots_4_io_uop_dst_rtype : _GEN_13877 ? _slots_3_io_uop_dst_rtype : _GEN_13553 ? _slots_2_io_uop_dst_rtype : _GEN_13229 ? _slots_1_io_uop_dst_rtype : _GEN_12906 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_0_lrs1_rtype = _GEN_25541 ? _slots_39_io_uop_lrs1_rtype : _GEN_25217 ? _slots_38_io_uop_lrs1_rtype : _GEN_24893 ? _slots_37_io_uop_lrs1_rtype : _GEN_24569 ? _slots_36_io_uop_lrs1_rtype : _GEN_24245 ? _slots_35_io_uop_lrs1_rtype : _GEN_23921 ? _slots_34_io_uop_lrs1_rtype : _GEN_23597 ? _slots_33_io_uop_lrs1_rtype : _GEN_23273 ? _slots_32_io_uop_lrs1_rtype : _GEN_22949 ? _slots_31_io_uop_lrs1_rtype : _GEN_22625 ? _slots_30_io_uop_lrs1_rtype : _GEN_22301 ? _slots_29_io_uop_lrs1_rtype : _GEN_21977 ? _slots_28_io_uop_lrs1_rtype : _GEN_21653 ? _slots_27_io_uop_lrs1_rtype : _GEN_21329 ? _slots_26_io_uop_lrs1_rtype : _GEN_21005 ? _slots_25_io_uop_lrs1_rtype : _GEN_20681 ? _slots_24_io_uop_lrs1_rtype : _GEN_20357 ? _slots_23_io_uop_lrs1_rtype : _GEN_20033 ? _slots_22_io_uop_lrs1_rtype : _GEN_19709 ? _slots_21_io_uop_lrs1_rtype : _GEN_19385 ? _slots_20_io_uop_lrs1_rtype : _GEN_19061 ? _slots_19_io_uop_lrs1_rtype : _GEN_18737 ? _slots_18_io_uop_lrs1_rtype : _GEN_18413 ? _slots_17_io_uop_lrs1_rtype : _GEN_18089 ? _slots_16_io_uop_lrs1_rtype : _GEN_17765 ? _slots_15_io_uop_lrs1_rtype : _GEN_17441 ? _slots_14_io_uop_lrs1_rtype : _GEN_17117 ? _slots_13_io_uop_lrs1_rtype : _GEN_16793 ? _slots_12_io_uop_lrs1_rtype : _GEN_16469 ? _slots_11_io_uop_lrs1_rtype : _GEN_16145 ? _slots_10_io_uop_lrs1_rtype : _GEN_15821 ? _slots_9_io_uop_lrs1_rtype : _GEN_15497 ? _slots_8_io_uop_lrs1_rtype : _GEN_15173 ? _slots_7_io_uop_lrs1_rtype : _GEN_14849 ? _slots_6_io_uop_lrs1_rtype : _GEN_14525 ? _slots_5_io_uop_lrs1_rtype : _GEN_14201 ? _slots_4_io_uop_lrs1_rtype : _GEN_13877 ? _slots_3_io_uop_lrs1_rtype : _GEN_13553 ? _slots_2_io_uop_lrs1_rtype : _GEN_13229 ? _slots_1_io_uop_lrs1_rtype : _GEN_12906 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_0_lrs2_rtype = _GEN_25541 ? _slots_39_io_uop_lrs2_rtype : _GEN_25217 ? _slots_38_io_uop_lrs2_rtype : _GEN_24893 ? _slots_37_io_uop_lrs2_rtype : _GEN_24569 ? _slots_36_io_uop_lrs2_rtype : _GEN_24245 ? _slots_35_io_uop_lrs2_rtype : _GEN_23921 ? _slots_34_io_uop_lrs2_rtype : _GEN_23597 ? _slots_33_io_uop_lrs2_rtype : _GEN_23273 ? _slots_32_io_uop_lrs2_rtype : _GEN_22949 ? _slots_31_io_uop_lrs2_rtype : _GEN_22625 ? _slots_30_io_uop_lrs2_rtype : _GEN_22301 ? _slots_29_io_uop_lrs2_rtype : _GEN_21977 ? _slots_28_io_uop_lrs2_rtype : _GEN_21653 ? _slots_27_io_uop_lrs2_rtype : _GEN_21329 ? _slots_26_io_uop_lrs2_rtype : _GEN_21005 ? _slots_25_io_uop_lrs2_rtype : _GEN_20681 ? _slots_24_io_uop_lrs2_rtype : _GEN_20357 ? _slots_23_io_uop_lrs2_rtype : _GEN_20033 ? _slots_22_io_uop_lrs2_rtype : _GEN_19709 ? _slots_21_io_uop_lrs2_rtype : _GEN_19385 ? _slots_20_io_uop_lrs2_rtype : _GEN_19061 ? _slots_19_io_uop_lrs2_rtype : _GEN_18737 ? _slots_18_io_uop_lrs2_rtype : _GEN_18413 ? _slots_17_io_uop_lrs2_rtype : _GEN_18089 ? _slots_16_io_uop_lrs2_rtype : _GEN_17765 ? _slots_15_io_uop_lrs2_rtype : _GEN_17441 ? _slots_14_io_uop_lrs2_rtype : _GEN_17117 ? _slots_13_io_uop_lrs2_rtype : _GEN_16793 ? _slots_12_io_uop_lrs2_rtype : _GEN_16469 ? _slots_11_io_uop_lrs2_rtype : _GEN_16145 ? _slots_10_io_uop_lrs2_rtype : _GEN_15821 ? _slots_9_io_uop_lrs2_rtype : _GEN_15497 ? _slots_8_io_uop_lrs2_rtype : _GEN_15173 ? _slots_7_io_uop_lrs2_rtype : _GEN_14849 ? _slots_6_io_uop_lrs2_rtype : _GEN_14525 ? _slots_5_io_uop_lrs2_rtype : _GEN_14201 ? _slots_4_io_uop_lrs2_rtype : _GEN_13877 ? _slots_3_io_uop_lrs2_rtype : _GEN_13553 ? _slots_2_io_uop_lrs2_rtype : _GEN_13229 ? _slots_1_io_uop_lrs2_rtype : _GEN_12906 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_0_fp_val = _GEN_25541 ? _slots_39_io_uop_fp_val : _GEN_25217 ? _slots_38_io_uop_fp_val : _GEN_24893 ? _slots_37_io_uop_fp_val : _GEN_24569 ? _slots_36_io_uop_fp_val : _GEN_24245 ? _slots_35_io_uop_fp_val : _GEN_23921 ? _slots_34_io_uop_fp_val : _GEN_23597 ? _slots_33_io_uop_fp_val : _GEN_23273 ? _slots_32_io_uop_fp_val : _GEN_22949 ? _slots_31_io_uop_fp_val : _GEN_22625 ? _slots_30_io_uop_fp_val : _GEN_22301 ? _slots_29_io_uop_fp_val : _GEN_21977 ? _slots_28_io_uop_fp_val : _GEN_21653 ? _slots_27_io_uop_fp_val : _GEN_21329 ? _slots_26_io_uop_fp_val : _GEN_21005 ? _slots_25_io_uop_fp_val : _GEN_20681 ? _slots_24_io_uop_fp_val : _GEN_20357 ? _slots_23_io_uop_fp_val : _GEN_20033 ? _slots_22_io_uop_fp_val : _GEN_19709 ? _slots_21_io_uop_fp_val : _GEN_19385 ? _slots_20_io_uop_fp_val : _GEN_19061 ? _slots_19_io_uop_fp_val : _GEN_18737 ? _slots_18_io_uop_fp_val : _GEN_18413 ? _slots_17_io_uop_fp_val : _GEN_18089 ? _slots_16_io_uop_fp_val : _GEN_17765 ? _slots_15_io_uop_fp_val : _GEN_17441 ? _slots_14_io_uop_fp_val : _GEN_17117 ? _slots_13_io_uop_fp_val : _GEN_16793 ? _slots_12_io_uop_fp_val : _GEN_16469 ? _slots_11_io_uop_fp_val : _GEN_16145 ? _slots_10_io_uop_fp_val : _GEN_15821 ? _slots_9_io_uop_fp_val : _GEN_15497 ? _slots_8_io_uop_fp_val : _GEN_15173 ? _slots_7_io_uop_fp_val : _GEN_14849 ? _slots_6_io_uop_fp_val : _GEN_14525 ? _slots_5_io_uop_fp_val : _GEN_14201 ? _slots_4_io_uop_fp_val : _GEN_13877 ? _slots_3_io_uop_fp_val : _GEN_13553 ? _slots_2_io_uop_fp_val : _GEN_13229 ? _slots_1_io_uop_fp_val : _GEN_12906 & _slots_0_io_uop_fp_val;
  assign io_iss_uops_1_uopc = _GEN_596 ? _slots_39_io_uop_uopc : _GEN_586 ? _slots_38_io_uop_uopc : _GEN_599 ? _slots_37_io_uop_uopc : _GEN_561 ? _slots_36_io_uop_uopc : _GEN_547 ? _slots_35_io_uop_uopc : _GEN_530 ? _slots_34_io_uop_uopc : _GEN_516 ? _slots_33_io_uop_uopc : _GEN_533 ? _slots_32_io_uop_uopc : _GEN_491 ? _slots_31_io_uop_uopc : _GEN_477 ? _slots_30_io_uop_uopc : _GEN_460 ? _slots_29_io_uop_uopc : _GEN_446 ? _slots_28_io_uop_uopc : _GEN_463 ? _slots_27_io_uop_uopc : _GEN_421 ? _slots_26_io_uop_uopc : _GEN_407 ? _slots_25_io_uop_uopc : _GEN_390 ? _slots_24_io_uop_uopc : _GEN_376 ? _slots_23_io_uop_uopc : _GEN_393 ? _slots_22_io_uop_uopc : _GEN_351 ? _slots_21_io_uop_uopc : _GEN_337 ? _slots_20_io_uop_uopc : _GEN_320 ? _slots_19_io_uop_uopc : _GEN_306 ? _slots_18_io_uop_uopc : _GEN_323 ? _slots_17_io_uop_uopc : _GEN_281 ? _slots_16_io_uop_uopc : _GEN_267 ? _slots_15_io_uop_uopc : _GEN_250 ? _slots_14_io_uop_uopc : _GEN_236 ? _slots_13_io_uop_uopc : _GEN_253 ? _slots_12_io_uop_uopc : _GEN_211 ? _slots_11_io_uop_uopc : _GEN_197 ? _slots_10_io_uop_uopc : _GEN_180 ? _slots_9_io_uop_uopc : _GEN_166 ? _slots_8_io_uop_uopc : _GEN_183 ? _slots_7_io_uop_uopc : _GEN_141 ? _slots_6_io_uop_uopc : _GEN_127 ? _slots_5_io_uop_uopc : _GEN_110 ? _slots_4_io_uop_uopc : _GEN_94 ? _slots_3_io_uop_uopc : _GEN_113 ? _slots_2_io_uop_uopc : _GEN_44 ? _slots_1_io_uop_uopc : _GEN_12987 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_1_is_rvc = _GEN_596 ? _slots_39_io_uop_is_rvc : _GEN_586 ? _slots_38_io_uop_is_rvc : _GEN_599 ? _slots_37_io_uop_is_rvc : _GEN_561 ? _slots_36_io_uop_is_rvc : _GEN_547 ? _slots_35_io_uop_is_rvc : _GEN_530 ? _slots_34_io_uop_is_rvc : _GEN_516 ? _slots_33_io_uop_is_rvc : _GEN_533 ? _slots_32_io_uop_is_rvc : _GEN_491 ? _slots_31_io_uop_is_rvc : _GEN_477 ? _slots_30_io_uop_is_rvc : _GEN_460 ? _slots_29_io_uop_is_rvc : _GEN_446 ? _slots_28_io_uop_is_rvc : _GEN_463 ? _slots_27_io_uop_is_rvc : _GEN_421 ? _slots_26_io_uop_is_rvc : _GEN_407 ? _slots_25_io_uop_is_rvc : _GEN_390 ? _slots_24_io_uop_is_rvc : _GEN_376 ? _slots_23_io_uop_is_rvc : _GEN_393 ? _slots_22_io_uop_is_rvc : _GEN_351 ? _slots_21_io_uop_is_rvc : _GEN_337 ? _slots_20_io_uop_is_rvc : _GEN_320 ? _slots_19_io_uop_is_rvc : _GEN_306 ? _slots_18_io_uop_is_rvc : _GEN_323 ? _slots_17_io_uop_is_rvc : _GEN_281 ? _slots_16_io_uop_is_rvc : _GEN_267 ? _slots_15_io_uop_is_rvc : _GEN_250 ? _slots_14_io_uop_is_rvc : _GEN_236 ? _slots_13_io_uop_is_rvc : _GEN_253 ? _slots_12_io_uop_is_rvc : _GEN_211 ? _slots_11_io_uop_is_rvc : _GEN_197 ? _slots_10_io_uop_is_rvc : _GEN_180 ? _slots_9_io_uop_is_rvc : _GEN_166 ? _slots_8_io_uop_is_rvc : _GEN_183 ? _slots_7_io_uop_is_rvc : _GEN_141 ? _slots_6_io_uop_is_rvc : _GEN_127 ? _slots_5_io_uop_is_rvc : _GEN_110 ? _slots_4_io_uop_is_rvc : _GEN_94 ? _slots_3_io_uop_is_rvc : _GEN_113 ? _slots_2_io_uop_is_rvc : _GEN_44 ? _slots_1_io_uop_is_rvc : _GEN_12987 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_1_fu_code = _GEN_596 ? _slots_39_io_uop_fu_code : _GEN_586 ? _slots_38_io_uop_fu_code : _GEN_599 ? _slots_37_io_uop_fu_code : _GEN_561 ? _slots_36_io_uop_fu_code : _GEN_547 ? _slots_35_io_uop_fu_code : _GEN_530 ? _slots_34_io_uop_fu_code : _GEN_516 ? _slots_33_io_uop_fu_code : _GEN_533 ? _slots_32_io_uop_fu_code : _GEN_491 ? _slots_31_io_uop_fu_code : _GEN_477 ? _slots_30_io_uop_fu_code : _GEN_460 ? _slots_29_io_uop_fu_code : _GEN_446 ? _slots_28_io_uop_fu_code : _GEN_463 ? _slots_27_io_uop_fu_code : _GEN_421 ? _slots_26_io_uop_fu_code : _GEN_407 ? _slots_25_io_uop_fu_code : _GEN_390 ? _slots_24_io_uop_fu_code : _GEN_376 ? _slots_23_io_uop_fu_code : _GEN_393 ? _slots_22_io_uop_fu_code : _GEN_351 ? _slots_21_io_uop_fu_code : _GEN_337 ? _slots_20_io_uop_fu_code : _GEN_320 ? _slots_19_io_uop_fu_code : _GEN_306 ? _slots_18_io_uop_fu_code : _GEN_323 ? _slots_17_io_uop_fu_code : _GEN_281 ? _slots_16_io_uop_fu_code : _GEN_267 ? _slots_15_io_uop_fu_code : _GEN_250 ? _slots_14_io_uop_fu_code : _GEN_236 ? _slots_13_io_uop_fu_code : _GEN_253 ? _slots_12_io_uop_fu_code : _GEN_211 ? _slots_11_io_uop_fu_code : _GEN_197 ? _slots_10_io_uop_fu_code : _GEN_180 ? _slots_9_io_uop_fu_code : _GEN_166 ? _slots_8_io_uop_fu_code : _GEN_183 ? _slots_7_io_uop_fu_code : _GEN_141 ? _slots_6_io_uop_fu_code : _GEN_127 ? _slots_5_io_uop_fu_code : _GEN_110 ? _slots_4_io_uop_fu_code : _GEN_94 ? _slots_3_io_uop_fu_code : _GEN_113 ? _slots_2_io_uop_fu_code : _GEN_44 ? _slots_1_io_uop_fu_code : _GEN_12987 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_1_iw_p1_poisoned = _GEN_596 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_586 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_599 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_561 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_547 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_530 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_516 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_533 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_491 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_477 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_460 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_446 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_463 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_421 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_407 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_390 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_376 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_393 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_351 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_337 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_320 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_306 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_323 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_281 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_267 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_250 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_236 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_253 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_211 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_197 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_180 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_166 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_183 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_141 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_127 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_110 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_94 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_113 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_44 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_12987 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_1_iw_p2_poisoned = _GEN_596 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_586 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_599 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_561 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_547 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_530 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_516 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_533 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_491 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_477 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_460 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_446 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_463 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_421 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_407 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_390 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_376 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_393 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_351 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_337 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_320 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_306 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_323 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_281 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_267 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_250 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_236 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_253 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_211 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_197 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_180 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_166 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_183 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_141 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_127 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_110 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_94 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_113 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_44 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_12987 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_1_is_br = _GEN_596 ? _slots_39_io_uop_is_br : _GEN_586 ? _slots_38_io_uop_is_br : _GEN_599 ? _slots_37_io_uop_is_br : _GEN_561 ? _slots_36_io_uop_is_br : _GEN_547 ? _slots_35_io_uop_is_br : _GEN_530 ? _slots_34_io_uop_is_br : _GEN_516 ? _slots_33_io_uop_is_br : _GEN_533 ? _slots_32_io_uop_is_br : _GEN_491 ? _slots_31_io_uop_is_br : _GEN_477 ? _slots_30_io_uop_is_br : _GEN_460 ? _slots_29_io_uop_is_br : _GEN_446 ? _slots_28_io_uop_is_br : _GEN_463 ? _slots_27_io_uop_is_br : _GEN_421 ? _slots_26_io_uop_is_br : _GEN_407 ? _slots_25_io_uop_is_br : _GEN_390 ? _slots_24_io_uop_is_br : _GEN_376 ? _slots_23_io_uop_is_br : _GEN_393 ? _slots_22_io_uop_is_br : _GEN_351 ? _slots_21_io_uop_is_br : _GEN_337 ? _slots_20_io_uop_is_br : _GEN_320 ? _slots_19_io_uop_is_br : _GEN_306 ? _slots_18_io_uop_is_br : _GEN_323 ? _slots_17_io_uop_is_br : _GEN_281 ? _slots_16_io_uop_is_br : _GEN_267 ? _slots_15_io_uop_is_br : _GEN_250 ? _slots_14_io_uop_is_br : _GEN_236 ? _slots_13_io_uop_is_br : _GEN_253 ? _slots_12_io_uop_is_br : _GEN_211 ? _slots_11_io_uop_is_br : _GEN_197 ? _slots_10_io_uop_is_br : _GEN_180 ? _slots_9_io_uop_is_br : _GEN_166 ? _slots_8_io_uop_is_br : _GEN_183 ? _slots_7_io_uop_is_br : _GEN_141 ? _slots_6_io_uop_is_br : _GEN_127 ? _slots_5_io_uop_is_br : _GEN_110 ? _slots_4_io_uop_is_br : _GEN_94 ? _slots_3_io_uop_is_br : _GEN_113 ? _slots_2_io_uop_is_br : _GEN_44 ? _slots_1_io_uop_is_br : _GEN_12987 & _slots_0_io_uop_is_br;
  assign io_iss_uops_1_is_jalr = _GEN_596 ? _slots_39_io_uop_is_jalr : _GEN_586 ? _slots_38_io_uop_is_jalr : _GEN_599 ? _slots_37_io_uop_is_jalr : _GEN_561 ? _slots_36_io_uop_is_jalr : _GEN_547 ? _slots_35_io_uop_is_jalr : _GEN_530 ? _slots_34_io_uop_is_jalr : _GEN_516 ? _slots_33_io_uop_is_jalr : _GEN_533 ? _slots_32_io_uop_is_jalr : _GEN_491 ? _slots_31_io_uop_is_jalr : _GEN_477 ? _slots_30_io_uop_is_jalr : _GEN_460 ? _slots_29_io_uop_is_jalr : _GEN_446 ? _slots_28_io_uop_is_jalr : _GEN_463 ? _slots_27_io_uop_is_jalr : _GEN_421 ? _slots_26_io_uop_is_jalr : _GEN_407 ? _slots_25_io_uop_is_jalr : _GEN_390 ? _slots_24_io_uop_is_jalr : _GEN_376 ? _slots_23_io_uop_is_jalr : _GEN_393 ? _slots_22_io_uop_is_jalr : _GEN_351 ? _slots_21_io_uop_is_jalr : _GEN_337 ? _slots_20_io_uop_is_jalr : _GEN_320 ? _slots_19_io_uop_is_jalr : _GEN_306 ? _slots_18_io_uop_is_jalr : _GEN_323 ? _slots_17_io_uop_is_jalr : _GEN_281 ? _slots_16_io_uop_is_jalr : _GEN_267 ? _slots_15_io_uop_is_jalr : _GEN_250 ? _slots_14_io_uop_is_jalr : _GEN_236 ? _slots_13_io_uop_is_jalr : _GEN_253 ? _slots_12_io_uop_is_jalr : _GEN_211 ? _slots_11_io_uop_is_jalr : _GEN_197 ? _slots_10_io_uop_is_jalr : _GEN_180 ? _slots_9_io_uop_is_jalr : _GEN_166 ? _slots_8_io_uop_is_jalr : _GEN_183 ? _slots_7_io_uop_is_jalr : _GEN_141 ? _slots_6_io_uop_is_jalr : _GEN_127 ? _slots_5_io_uop_is_jalr : _GEN_110 ? _slots_4_io_uop_is_jalr : _GEN_94 ? _slots_3_io_uop_is_jalr : _GEN_113 ? _slots_2_io_uop_is_jalr : _GEN_44 ? _slots_1_io_uop_is_jalr : _GEN_12987 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_1_is_jal = _GEN_596 ? _slots_39_io_uop_is_jal : _GEN_586 ? _slots_38_io_uop_is_jal : _GEN_599 ? _slots_37_io_uop_is_jal : _GEN_561 ? _slots_36_io_uop_is_jal : _GEN_547 ? _slots_35_io_uop_is_jal : _GEN_530 ? _slots_34_io_uop_is_jal : _GEN_516 ? _slots_33_io_uop_is_jal : _GEN_533 ? _slots_32_io_uop_is_jal : _GEN_491 ? _slots_31_io_uop_is_jal : _GEN_477 ? _slots_30_io_uop_is_jal : _GEN_460 ? _slots_29_io_uop_is_jal : _GEN_446 ? _slots_28_io_uop_is_jal : _GEN_463 ? _slots_27_io_uop_is_jal : _GEN_421 ? _slots_26_io_uop_is_jal : _GEN_407 ? _slots_25_io_uop_is_jal : _GEN_390 ? _slots_24_io_uop_is_jal : _GEN_376 ? _slots_23_io_uop_is_jal : _GEN_393 ? _slots_22_io_uop_is_jal : _GEN_351 ? _slots_21_io_uop_is_jal : _GEN_337 ? _slots_20_io_uop_is_jal : _GEN_320 ? _slots_19_io_uop_is_jal : _GEN_306 ? _slots_18_io_uop_is_jal : _GEN_323 ? _slots_17_io_uop_is_jal : _GEN_281 ? _slots_16_io_uop_is_jal : _GEN_267 ? _slots_15_io_uop_is_jal : _GEN_250 ? _slots_14_io_uop_is_jal : _GEN_236 ? _slots_13_io_uop_is_jal : _GEN_253 ? _slots_12_io_uop_is_jal : _GEN_211 ? _slots_11_io_uop_is_jal : _GEN_197 ? _slots_10_io_uop_is_jal : _GEN_180 ? _slots_9_io_uop_is_jal : _GEN_166 ? _slots_8_io_uop_is_jal : _GEN_183 ? _slots_7_io_uop_is_jal : _GEN_141 ? _slots_6_io_uop_is_jal : _GEN_127 ? _slots_5_io_uop_is_jal : _GEN_110 ? _slots_4_io_uop_is_jal : _GEN_94 ? _slots_3_io_uop_is_jal : _GEN_113 ? _slots_2_io_uop_is_jal : _GEN_44 ? _slots_1_io_uop_is_jal : _GEN_12987 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_1_is_sfb = _GEN_596 ? _slots_39_io_uop_is_sfb : _GEN_586 ? _slots_38_io_uop_is_sfb : _GEN_599 ? _slots_37_io_uop_is_sfb : _GEN_561 ? _slots_36_io_uop_is_sfb : _GEN_547 ? _slots_35_io_uop_is_sfb : _GEN_530 ? _slots_34_io_uop_is_sfb : _GEN_516 ? _slots_33_io_uop_is_sfb : _GEN_533 ? _slots_32_io_uop_is_sfb : _GEN_491 ? _slots_31_io_uop_is_sfb : _GEN_477 ? _slots_30_io_uop_is_sfb : _GEN_460 ? _slots_29_io_uop_is_sfb : _GEN_446 ? _slots_28_io_uop_is_sfb : _GEN_463 ? _slots_27_io_uop_is_sfb : _GEN_421 ? _slots_26_io_uop_is_sfb : _GEN_407 ? _slots_25_io_uop_is_sfb : _GEN_390 ? _slots_24_io_uop_is_sfb : _GEN_376 ? _slots_23_io_uop_is_sfb : _GEN_393 ? _slots_22_io_uop_is_sfb : _GEN_351 ? _slots_21_io_uop_is_sfb : _GEN_337 ? _slots_20_io_uop_is_sfb : _GEN_320 ? _slots_19_io_uop_is_sfb : _GEN_306 ? _slots_18_io_uop_is_sfb : _GEN_323 ? _slots_17_io_uop_is_sfb : _GEN_281 ? _slots_16_io_uop_is_sfb : _GEN_267 ? _slots_15_io_uop_is_sfb : _GEN_250 ? _slots_14_io_uop_is_sfb : _GEN_236 ? _slots_13_io_uop_is_sfb : _GEN_253 ? _slots_12_io_uop_is_sfb : _GEN_211 ? _slots_11_io_uop_is_sfb : _GEN_197 ? _slots_10_io_uop_is_sfb : _GEN_180 ? _slots_9_io_uop_is_sfb : _GEN_166 ? _slots_8_io_uop_is_sfb : _GEN_183 ? _slots_7_io_uop_is_sfb : _GEN_141 ? _slots_6_io_uop_is_sfb : _GEN_127 ? _slots_5_io_uop_is_sfb : _GEN_110 ? _slots_4_io_uop_is_sfb : _GEN_94 ? _slots_3_io_uop_is_sfb : _GEN_113 ? _slots_2_io_uop_is_sfb : _GEN_44 ? _slots_1_io_uop_is_sfb : _GEN_12987 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_1_br_mask = _GEN_596 ? _slots_39_io_uop_br_mask : _GEN_586 ? _slots_38_io_uop_br_mask : _GEN_599 ? _slots_37_io_uop_br_mask : _GEN_561 ? _slots_36_io_uop_br_mask : _GEN_547 ? _slots_35_io_uop_br_mask : _GEN_530 ? _slots_34_io_uop_br_mask : _GEN_516 ? _slots_33_io_uop_br_mask : _GEN_533 ? _slots_32_io_uop_br_mask : _GEN_491 ? _slots_31_io_uop_br_mask : _GEN_477 ? _slots_30_io_uop_br_mask : _GEN_460 ? _slots_29_io_uop_br_mask : _GEN_446 ? _slots_28_io_uop_br_mask : _GEN_463 ? _slots_27_io_uop_br_mask : _GEN_421 ? _slots_26_io_uop_br_mask : _GEN_407 ? _slots_25_io_uop_br_mask : _GEN_390 ? _slots_24_io_uop_br_mask : _GEN_376 ? _slots_23_io_uop_br_mask : _GEN_393 ? _slots_22_io_uop_br_mask : _GEN_351 ? _slots_21_io_uop_br_mask : _GEN_337 ? _slots_20_io_uop_br_mask : _GEN_320 ? _slots_19_io_uop_br_mask : _GEN_306 ? _slots_18_io_uop_br_mask : _GEN_323 ? _slots_17_io_uop_br_mask : _GEN_281 ? _slots_16_io_uop_br_mask : _GEN_267 ? _slots_15_io_uop_br_mask : _GEN_250 ? _slots_14_io_uop_br_mask : _GEN_236 ? _slots_13_io_uop_br_mask : _GEN_253 ? _slots_12_io_uop_br_mask : _GEN_211 ? _slots_11_io_uop_br_mask : _GEN_197 ? _slots_10_io_uop_br_mask : _GEN_180 ? _slots_9_io_uop_br_mask : _GEN_166 ? _slots_8_io_uop_br_mask : _GEN_183 ? _slots_7_io_uop_br_mask : _GEN_141 ? _slots_6_io_uop_br_mask : _GEN_127 ? _slots_5_io_uop_br_mask : _GEN_110 ? _slots_4_io_uop_br_mask : _GEN_94 ? _slots_3_io_uop_br_mask : _GEN_113 ? _slots_2_io_uop_br_mask : _GEN_44 ? _slots_1_io_uop_br_mask : _GEN_12987 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_1_br_tag = _GEN_596 ? _slots_39_io_uop_br_tag : _GEN_586 ? _slots_38_io_uop_br_tag : _GEN_599 ? _slots_37_io_uop_br_tag : _GEN_561 ? _slots_36_io_uop_br_tag : _GEN_547 ? _slots_35_io_uop_br_tag : _GEN_530 ? _slots_34_io_uop_br_tag : _GEN_516 ? _slots_33_io_uop_br_tag : _GEN_533 ? _slots_32_io_uop_br_tag : _GEN_491 ? _slots_31_io_uop_br_tag : _GEN_477 ? _slots_30_io_uop_br_tag : _GEN_460 ? _slots_29_io_uop_br_tag : _GEN_446 ? _slots_28_io_uop_br_tag : _GEN_463 ? _slots_27_io_uop_br_tag : _GEN_421 ? _slots_26_io_uop_br_tag : _GEN_407 ? _slots_25_io_uop_br_tag : _GEN_390 ? _slots_24_io_uop_br_tag : _GEN_376 ? _slots_23_io_uop_br_tag : _GEN_393 ? _slots_22_io_uop_br_tag : _GEN_351 ? _slots_21_io_uop_br_tag : _GEN_337 ? _slots_20_io_uop_br_tag : _GEN_320 ? _slots_19_io_uop_br_tag : _GEN_306 ? _slots_18_io_uop_br_tag : _GEN_323 ? _slots_17_io_uop_br_tag : _GEN_281 ? _slots_16_io_uop_br_tag : _GEN_267 ? _slots_15_io_uop_br_tag : _GEN_250 ? _slots_14_io_uop_br_tag : _GEN_236 ? _slots_13_io_uop_br_tag : _GEN_253 ? _slots_12_io_uop_br_tag : _GEN_211 ? _slots_11_io_uop_br_tag : _GEN_197 ? _slots_10_io_uop_br_tag : _GEN_180 ? _slots_9_io_uop_br_tag : _GEN_166 ? _slots_8_io_uop_br_tag : _GEN_183 ? _slots_7_io_uop_br_tag : _GEN_141 ? _slots_6_io_uop_br_tag : _GEN_127 ? _slots_5_io_uop_br_tag : _GEN_110 ? _slots_4_io_uop_br_tag : _GEN_94 ? _slots_3_io_uop_br_tag : _GEN_113 ? _slots_2_io_uop_br_tag : _GEN_44 ? _slots_1_io_uop_br_tag : _GEN_12987 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_1_ftq_idx = _GEN_596 ? _slots_39_io_uop_ftq_idx : _GEN_586 ? _slots_38_io_uop_ftq_idx : _GEN_599 ? _slots_37_io_uop_ftq_idx : _GEN_561 ? _slots_36_io_uop_ftq_idx : _GEN_547 ? _slots_35_io_uop_ftq_idx : _GEN_530 ? _slots_34_io_uop_ftq_idx : _GEN_516 ? _slots_33_io_uop_ftq_idx : _GEN_533 ? _slots_32_io_uop_ftq_idx : _GEN_491 ? _slots_31_io_uop_ftq_idx : _GEN_477 ? _slots_30_io_uop_ftq_idx : _GEN_460 ? _slots_29_io_uop_ftq_idx : _GEN_446 ? _slots_28_io_uop_ftq_idx : _GEN_463 ? _slots_27_io_uop_ftq_idx : _GEN_421 ? _slots_26_io_uop_ftq_idx : _GEN_407 ? _slots_25_io_uop_ftq_idx : _GEN_390 ? _slots_24_io_uop_ftq_idx : _GEN_376 ? _slots_23_io_uop_ftq_idx : _GEN_393 ? _slots_22_io_uop_ftq_idx : _GEN_351 ? _slots_21_io_uop_ftq_idx : _GEN_337 ? _slots_20_io_uop_ftq_idx : _GEN_320 ? _slots_19_io_uop_ftq_idx : _GEN_306 ? _slots_18_io_uop_ftq_idx : _GEN_323 ? _slots_17_io_uop_ftq_idx : _GEN_281 ? _slots_16_io_uop_ftq_idx : _GEN_267 ? _slots_15_io_uop_ftq_idx : _GEN_250 ? _slots_14_io_uop_ftq_idx : _GEN_236 ? _slots_13_io_uop_ftq_idx : _GEN_253 ? _slots_12_io_uop_ftq_idx : _GEN_211 ? _slots_11_io_uop_ftq_idx : _GEN_197 ? _slots_10_io_uop_ftq_idx : _GEN_180 ? _slots_9_io_uop_ftq_idx : _GEN_166 ? _slots_8_io_uop_ftq_idx : _GEN_183 ? _slots_7_io_uop_ftq_idx : _GEN_141 ? _slots_6_io_uop_ftq_idx : _GEN_127 ? _slots_5_io_uop_ftq_idx : _GEN_110 ? _slots_4_io_uop_ftq_idx : _GEN_94 ? _slots_3_io_uop_ftq_idx : _GEN_113 ? _slots_2_io_uop_ftq_idx : _GEN_44 ? _slots_1_io_uop_ftq_idx : _GEN_12987 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_1_edge_inst = _GEN_596 ? _slots_39_io_uop_edge_inst : _GEN_586 ? _slots_38_io_uop_edge_inst : _GEN_599 ? _slots_37_io_uop_edge_inst : _GEN_561 ? _slots_36_io_uop_edge_inst : _GEN_547 ? _slots_35_io_uop_edge_inst : _GEN_530 ? _slots_34_io_uop_edge_inst : _GEN_516 ? _slots_33_io_uop_edge_inst : _GEN_533 ? _slots_32_io_uop_edge_inst : _GEN_491 ? _slots_31_io_uop_edge_inst : _GEN_477 ? _slots_30_io_uop_edge_inst : _GEN_460 ? _slots_29_io_uop_edge_inst : _GEN_446 ? _slots_28_io_uop_edge_inst : _GEN_463 ? _slots_27_io_uop_edge_inst : _GEN_421 ? _slots_26_io_uop_edge_inst : _GEN_407 ? _slots_25_io_uop_edge_inst : _GEN_390 ? _slots_24_io_uop_edge_inst : _GEN_376 ? _slots_23_io_uop_edge_inst : _GEN_393 ? _slots_22_io_uop_edge_inst : _GEN_351 ? _slots_21_io_uop_edge_inst : _GEN_337 ? _slots_20_io_uop_edge_inst : _GEN_320 ? _slots_19_io_uop_edge_inst : _GEN_306 ? _slots_18_io_uop_edge_inst : _GEN_323 ? _slots_17_io_uop_edge_inst : _GEN_281 ? _slots_16_io_uop_edge_inst : _GEN_267 ? _slots_15_io_uop_edge_inst : _GEN_250 ? _slots_14_io_uop_edge_inst : _GEN_236 ? _slots_13_io_uop_edge_inst : _GEN_253 ? _slots_12_io_uop_edge_inst : _GEN_211 ? _slots_11_io_uop_edge_inst : _GEN_197 ? _slots_10_io_uop_edge_inst : _GEN_180 ? _slots_9_io_uop_edge_inst : _GEN_166 ? _slots_8_io_uop_edge_inst : _GEN_183 ? _slots_7_io_uop_edge_inst : _GEN_141 ? _slots_6_io_uop_edge_inst : _GEN_127 ? _slots_5_io_uop_edge_inst : _GEN_110 ? _slots_4_io_uop_edge_inst : _GEN_94 ? _slots_3_io_uop_edge_inst : _GEN_113 ? _slots_2_io_uop_edge_inst : _GEN_44 ? _slots_1_io_uop_edge_inst : _GEN_12987 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_1_pc_lob = _GEN_596 ? _slots_39_io_uop_pc_lob : _GEN_586 ? _slots_38_io_uop_pc_lob : _GEN_599 ? _slots_37_io_uop_pc_lob : _GEN_561 ? _slots_36_io_uop_pc_lob : _GEN_547 ? _slots_35_io_uop_pc_lob : _GEN_530 ? _slots_34_io_uop_pc_lob : _GEN_516 ? _slots_33_io_uop_pc_lob : _GEN_533 ? _slots_32_io_uop_pc_lob : _GEN_491 ? _slots_31_io_uop_pc_lob : _GEN_477 ? _slots_30_io_uop_pc_lob : _GEN_460 ? _slots_29_io_uop_pc_lob : _GEN_446 ? _slots_28_io_uop_pc_lob : _GEN_463 ? _slots_27_io_uop_pc_lob : _GEN_421 ? _slots_26_io_uop_pc_lob : _GEN_407 ? _slots_25_io_uop_pc_lob : _GEN_390 ? _slots_24_io_uop_pc_lob : _GEN_376 ? _slots_23_io_uop_pc_lob : _GEN_393 ? _slots_22_io_uop_pc_lob : _GEN_351 ? _slots_21_io_uop_pc_lob : _GEN_337 ? _slots_20_io_uop_pc_lob : _GEN_320 ? _slots_19_io_uop_pc_lob : _GEN_306 ? _slots_18_io_uop_pc_lob : _GEN_323 ? _slots_17_io_uop_pc_lob : _GEN_281 ? _slots_16_io_uop_pc_lob : _GEN_267 ? _slots_15_io_uop_pc_lob : _GEN_250 ? _slots_14_io_uop_pc_lob : _GEN_236 ? _slots_13_io_uop_pc_lob : _GEN_253 ? _slots_12_io_uop_pc_lob : _GEN_211 ? _slots_11_io_uop_pc_lob : _GEN_197 ? _slots_10_io_uop_pc_lob : _GEN_180 ? _slots_9_io_uop_pc_lob : _GEN_166 ? _slots_8_io_uop_pc_lob : _GEN_183 ? _slots_7_io_uop_pc_lob : _GEN_141 ? _slots_6_io_uop_pc_lob : _GEN_127 ? _slots_5_io_uop_pc_lob : _GEN_110 ? _slots_4_io_uop_pc_lob : _GEN_94 ? _slots_3_io_uop_pc_lob : _GEN_113 ? _slots_2_io_uop_pc_lob : _GEN_44 ? _slots_1_io_uop_pc_lob : _GEN_12987 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_1_taken = _GEN_596 ? _slots_39_io_uop_taken : _GEN_586 ? _slots_38_io_uop_taken : _GEN_599 ? _slots_37_io_uop_taken : _GEN_561 ? _slots_36_io_uop_taken : _GEN_547 ? _slots_35_io_uop_taken : _GEN_530 ? _slots_34_io_uop_taken : _GEN_516 ? _slots_33_io_uop_taken : _GEN_533 ? _slots_32_io_uop_taken : _GEN_491 ? _slots_31_io_uop_taken : _GEN_477 ? _slots_30_io_uop_taken : _GEN_460 ? _slots_29_io_uop_taken : _GEN_446 ? _slots_28_io_uop_taken : _GEN_463 ? _slots_27_io_uop_taken : _GEN_421 ? _slots_26_io_uop_taken : _GEN_407 ? _slots_25_io_uop_taken : _GEN_390 ? _slots_24_io_uop_taken : _GEN_376 ? _slots_23_io_uop_taken : _GEN_393 ? _slots_22_io_uop_taken : _GEN_351 ? _slots_21_io_uop_taken : _GEN_337 ? _slots_20_io_uop_taken : _GEN_320 ? _slots_19_io_uop_taken : _GEN_306 ? _slots_18_io_uop_taken : _GEN_323 ? _slots_17_io_uop_taken : _GEN_281 ? _slots_16_io_uop_taken : _GEN_267 ? _slots_15_io_uop_taken : _GEN_250 ? _slots_14_io_uop_taken : _GEN_236 ? _slots_13_io_uop_taken : _GEN_253 ? _slots_12_io_uop_taken : _GEN_211 ? _slots_11_io_uop_taken : _GEN_197 ? _slots_10_io_uop_taken : _GEN_180 ? _slots_9_io_uop_taken : _GEN_166 ? _slots_8_io_uop_taken : _GEN_183 ? _slots_7_io_uop_taken : _GEN_141 ? _slots_6_io_uop_taken : _GEN_127 ? _slots_5_io_uop_taken : _GEN_110 ? _slots_4_io_uop_taken : _GEN_94 ? _slots_3_io_uop_taken : _GEN_113 ? _slots_2_io_uop_taken : _GEN_44 ? _slots_1_io_uop_taken : _GEN_12987 & _slots_0_io_uop_taken;
  assign io_iss_uops_1_imm_packed = _GEN_596 ? _slots_39_io_uop_imm_packed : _GEN_586 ? _slots_38_io_uop_imm_packed : _GEN_599 ? _slots_37_io_uop_imm_packed : _GEN_561 ? _slots_36_io_uop_imm_packed : _GEN_547 ? _slots_35_io_uop_imm_packed : _GEN_530 ? _slots_34_io_uop_imm_packed : _GEN_516 ? _slots_33_io_uop_imm_packed : _GEN_533 ? _slots_32_io_uop_imm_packed : _GEN_491 ? _slots_31_io_uop_imm_packed : _GEN_477 ? _slots_30_io_uop_imm_packed : _GEN_460 ? _slots_29_io_uop_imm_packed : _GEN_446 ? _slots_28_io_uop_imm_packed : _GEN_463 ? _slots_27_io_uop_imm_packed : _GEN_421 ? _slots_26_io_uop_imm_packed : _GEN_407 ? _slots_25_io_uop_imm_packed : _GEN_390 ? _slots_24_io_uop_imm_packed : _GEN_376 ? _slots_23_io_uop_imm_packed : _GEN_393 ? _slots_22_io_uop_imm_packed : _GEN_351 ? _slots_21_io_uop_imm_packed : _GEN_337 ? _slots_20_io_uop_imm_packed : _GEN_320 ? _slots_19_io_uop_imm_packed : _GEN_306 ? _slots_18_io_uop_imm_packed : _GEN_323 ? _slots_17_io_uop_imm_packed : _GEN_281 ? _slots_16_io_uop_imm_packed : _GEN_267 ? _slots_15_io_uop_imm_packed : _GEN_250 ? _slots_14_io_uop_imm_packed : _GEN_236 ? _slots_13_io_uop_imm_packed : _GEN_253 ? _slots_12_io_uop_imm_packed : _GEN_211 ? _slots_11_io_uop_imm_packed : _GEN_197 ? _slots_10_io_uop_imm_packed : _GEN_180 ? _slots_9_io_uop_imm_packed : _GEN_166 ? _slots_8_io_uop_imm_packed : _GEN_183 ? _slots_7_io_uop_imm_packed : _GEN_141 ? _slots_6_io_uop_imm_packed : _GEN_127 ? _slots_5_io_uop_imm_packed : _GEN_110 ? _slots_4_io_uop_imm_packed : _GEN_94 ? _slots_3_io_uop_imm_packed : _GEN_113 ? _slots_2_io_uop_imm_packed : _GEN_44 ? _slots_1_io_uop_imm_packed : _GEN_12987 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_1_rob_idx = _GEN_596 ? _slots_39_io_uop_rob_idx : _GEN_586 ? _slots_38_io_uop_rob_idx : _GEN_599 ? _slots_37_io_uop_rob_idx : _GEN_561 ? _slots_36_io_uop_rob_idx : _GEN_547 ? _slots_35_io_uop_rob_idx : _GEN_530 ? _slots_34_io_uop_rob_idx : _GEN_516 ? _slots_33_io_uop_rob_idx : _GEN_533 ? _slots_32_io_uop_rob_idx : _GEN_491 ? _slots_31_io_uop_rob_idx : _GEN_477 ? _slots_30_io_uop_rob_idx : _GEN_460 ? _slots_29_io_uop_rob_idx : _GEN_446 ? _slots_28_io_uop_rob_idx : _GEN_463 ? _slots_27_io_uop_rob_idx : _GEN_421 ? _slots_26_io_uop_rob_idx : _GEN_407 ? _slots_25_io_uop_rob_idx : _GEN_390 ? _slots_24_io_uop_rob_idx : _GEN_376 ? _slots_23_io_uop_rob_idx : _GEN_393 ? _slots_22_io_uop_rob_idx : _GEN_351 ? _slots_21_io_uop_rob_idx : _GEN_337 ? _slots_20_io_uop_rob_idx : _GEN_320 ? _slots_19_io_uop_rob_idx : _GEN_306 ? _slots_18_io_uop_rob_idx : _GEN_323 ? _slots_17_io_uop_rob_idx : _GEN_281 ? _slots_16_io_uop_rob_idx : _GEN_267 ? _slots_15_io_uop_rob_idx : _GEN_250 ? _slots_14_io_uop_rob_idx : _GEN_236 ? _slots_13_io_uop_rob_idx : _GEN_253 ? _slots_12_io_uop_rob_idx : _GEN_211 ? _slots_11_io_uop_rob_idx : _GEN_197 ? _slots_10_io_uop_rob_idx : _GEN_180 ? _slots_9_io_uop_rob_idx : _GEN_166 ? _slots_8_io_uop_rob_idx : _GEN_183 ? _slots_7_io_uop_rob_idx : _GEN_141 ? _slots_6_io_uop_rob_idx : _GEN_127 ? _slots_5_io_uop_rob_idx : _GEN_110 ? _slots_4_io_uop_rob_idx : _GEN_94 ? _slots_3_io_uop_rob_idx : _GEN_113 ? _slots_2_io_uop_rob_idx : _GEN_44 ? _slots_1_io_uop_rob_idx : _GEN_12987 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_1_ldq_idx = _GEN_596 ? _slots_39_io_uop_ldq_idx : _GEN_586 ? _slots_38_io_uop_ldq_idx : _GEN_599 ? _slots_37_io_uop_ldq_idx : _GEN_561 ? _slots_36_io_uop_ldq_idx : _GEN_547 ? _slots_35_io_uop_ldq_idx : _GEN_530 ? _slots_34_io_uop_ldq_idx : _GEN_516 ? _slots_33_io_uop_ldq_idx : _GEN_533 ? _slots_32_io_uop_ldq_idx : _GEN_491 ? _slots_31_io_uop_ldq_idx : _GEN_477 ? _slots_30_io_uop_ldq_idx : _GEN_460 ? _slots_29_io_uop_ldq_idx : _GEN_446 ? _slots_28_io_uop_ldq_idx : _GEN_463 ? _slots_27_io_uop_ldq_idx : _GEN_421 ? _slots_26_io_uop_ldq_idx : _GEN_407 ? _slots_25_io_uop_ldq_idx : _GEN_390 ? _slots_24_io_uop_ldq_idx : _GEN_376 ? _slots_23_io_uop_ldq_idx : _GEN_393 ? _slots_22_io_uop_ldq_idx : _GEN_351 ? _slots_21_io_uop_ldq_idx : _GEN_337 ? _slots_20_io_uop_ldq_idx : _GEN_320 ? _slots_19_io_uop_ldq_idx : _GEN_306 ? _slots_18_io_uop_ldq_idx : _GEN_323 ? _slots_17_io_uop_ldq_idx : _GEN_281 ? _slots_16_io_uop_ldq_idx : _GEN_267 ? _slots_15_io_uop_ldq_idx : _GEN_250 ? _slots_14_io_uop_ldq_idx : _GEN_236 ? _slots_13_io_uop_ldq_idx : _GEN_253 ? _slots_12_io_uop_ldq_idx : _GEN_211 ? _slots_11_io_uop_ldq_idx : _GEN_197 ? _slots_10_io_uop_ldq_idx : _GEN_180 ? _slots_9_io_uop_ldq_idx : _GEN_166 ? _slots_8_io_uop_ldq_idx : _GEN_183 ? _slots_7_io_uop_ldq_idx : _GEN_141 ? _slots_6_io_uop_ldq_idx : _GEN_127 ? _slots_5_io_uop_ldq_idx : _GEN_110 ? _slots_4_io_uop_ldq_idx : _GEN_94 ? _slots_3_io_uop_ldq_idx : _GEN_113 ? _slots_2_io_uop_ldq_idx : _GEN_44 ? _slots_1_io_uop_ldq_idx : _GEN_12987 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_1_stq_idx = _GEN_596 ? _slots_39_io_uop_stq_idx : _GEN_586 ? _slots_38_io_uop_stq_idx : _GEN_599 ? _slots_37_io_uop_stq_idx : _GEN_561 ? _slots_36_io_uop_stq_idx : _GEN_547 ? _slots_35_io_uop_stq_idx : _GEN_530 ? _slots_34_io_uop_stq_idx : _GEN_516 ? _slots_33_io_uop_stq_idx : _GEN_533 ? _slots_32_io_uop_stq_idx : _GEN_491 ? _slots_31_io_uop_stq_idx : _GEN_477 ? _slots_30_io_uop_stq_idx : _GEN_460 ? _slots_29_io_uop_stq_idx : _GEN_446 ? _slots_28_io_uop_stq_idx : _GEN_463 ? _slots_27_io_uop_stq_idx : _GEN_421 ? _slots_26_io_uop_stq_idx : _GEN_407 ? _slots_25_io_uop_stq_idx : _GEN_390 ? _slots_24_io_uop_stq_idx : _GEN_376 ? _slots_23_io_uop_stq_idx : _GEN_393 ? _slots_22_io_uop_stq_idx : _GEN_351 ? _slots_21_io_uop_stq_idx : _GEN_337 ? _slots_20_io_uop_stq_idx : _GEN_320 ? _slots_19_io_uop_stq_idx : _GEN_306 ? _slots_18_io_uop_stq_idx : _GEN_323 ? _slots_17_io_uop_stq_idx : _GEN_281 ? _slots_16_io_uop_stq_idx : _GEN_267 ? _slots_15_io_uop_stq_idx : _GEN_250 ? _slots_14_io_uop_stq_idx : _GEN_236 ? _slots_13_io_uop_stq_idx : _GEN_253 ? _slots_12_io_uop_stq_idx : _GEN_211 ? _slots_11_io_uop_stq_idx : _GEN_197 ? _slots_10_io_uop_stq_idx : _GEN_180 ? _slots_9_io_uop_stq_idx : _GEN_166 ? _slots_8_io_uop_stq_idx : _GEN_183 ? _slots_7_io_uop_stq_idx : _GEN_141 ? _slots_6_io_uop_stq_idx : _GEN_127 ? _slots_5_io_uop_stq_idx : _GEN_110 ? _slots_4_io_uop_stq_idx : _GEN_94 ? _slots_3_io_uop_stq_idx : _GEN_113 ? _slots_2_io_uop_stq_idx : _GEN_44 ? _slots_1_io_uop_stq_idx : _GEN_12987 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_1_pdst = _GEN_596 ? _slots_39_io_uop_pdst : _GEN_586 ? _slots_38_io_uop_pdst : _GEN_599 ? _slots_37_io_uop_pdst : _GEN_561 ? _slots_36_io_uop_pdst : _GEN_547 ? _slots_35_io_uop_pdst : _GEN_530 ? _slots_34_io_uop_pdst : _GEN_516 ? _slots_33_io_uop_pdst : _GEN_533 ? _slots_32_io_uop_pdst : _GEN_491 ? _slots_31_io_uop_pdst : _GEN_477 ? _slots_30_io_uop_pdst : _GEN_460 ? _slots_29_io_uop_pdst : _GEN_446 ? _slots_28_io_uop_pdst : _GEN_463 ? _slots_27_io_uop_pdst : _GEN_421 ? _slots_26_io_uop_pdst : _GEN_407 ? _slots_25_io_uop_pdst : _GEN_390 ? _slots_24_io_uop_pdst : _GEN_376 ? _slots_23_io_uop_pdst : _GEN_393 ? _slots_22_io_uop_pdst : _GEN_351 ? _slots_21_io_uop_pdst : _GEN_337 ? _slots_20_io_uop_pdst : _GEN_320 ? _slots_19_io_uop_pdst : _GEN_306 ? _slots_18_io_uop_pdst : _GEN_323 ? _slots_17_io_uop_pdst : _GEN_281 ? _slots_16_io_uop_pdst : _GEN_267 ? _slots_15_io_uop_pdst : _GEN_250 ? _slots_14_io_uop_pdst : _GEN_236 ? _slots_13_io_uop_pdst : _GEN_253 ? _slots_12_io_uop_pdst : _GEN_211 ? _slots_11_io_uop_pdst : _GEN_197 ? _slots_10_io_uop_pdst : _GEN_180 ? _slots_9_io_uop_pdst : _GEN_166 ? _slots_8_io_uop_pdst : _GEN_183 ? _slots_7_io_uop_pdst : _GEN_141 ? _slots_6_io_uop_pdst : _GEN_127 ? _slots_5_io_uop_pdst : _GEN_110 ? _slots_4_io_uop_pdst : _GEN_94 ? _slots_3_io_uop_pdst : _GEN_113 ? _slots_2_io_uop_pdst : _GEN_44 ? _slots_1_io_uop_pdst : _GEN_12987 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_1_prs1 = _GEN_596 ? _slots_39_io_uop_prs1 : _GEN_586 ? _slots_38_io_uop_prs1 : _GEN_599 ? _slots_37_io_uop_prs1 : _GEN_561 ? _slots_36_io_uop_prs1 : _GEN_547 ? _slots_35_io_uop_prs1 : _GEN_530 ? _slots_34_io_uop_prs1 : _GEN_516 ? _slots_33_io_uop_prs1 : _GEN_533 ? _slots_32_io_uop_prs1 : _GEN_491 ? _slots_31_io_uop_prs1 : _GEN_477 ? _slots_30_io_uop_prs1 : _GEN_460 ? _slots_29_io_uop_prs1 : _GEN_446 ? _slots_28_io_uop_prs1 : _GEN_463 ? _slots_27_io_uop_prs1 : _GEN_421 ? _slots_26_io_uop_prs1 : _GEN_407 ? _slots_25_io_uop_prs1 : _GEN_390 ? _slots_24_io_uop_prs1 : _GEN_376 ? _slots_23_io_uop_prs1 : _GEN_393 ? _slots_22_io_uop_prs1 : _GEN_351 ? _slots_21_io_uop_prs1 : _GEN_337 ? _slots_20_io_uop_prs1 : _GEN_320 ? _slots_19_io_uop_prs1 : _GEN_306 ? _slots_18_io_uop_prs1 : _GEN_323 ? _slots_17_io_uop_prs1 : _GEN_281 ? _slots_16_io_uop_prs1 : _GEN_267 ? _slots_15_io_uop_prs1 : _GEN_250 ? _slots_14_io_uop_prs1 : _GEN_236 ? _slots_13_io_uop_prs1 : _GEN_253 ? _slots_12_io_uop_prs1 : _GEN_211 ? _slots_11_io_uop_prs1 : _GEN_197 ? _slots_10_io_uop_prs1 : _GEN_180 ? _slots_9_io_uop_prs1 : _GEN_166 ? _slots_8_io_uop_prs1 : _GEN_183 ? _slots_7_io_uop_prs1 : _GEN_141 ? _slots_6_io_uop_prs1 : _GEN_127 ? _slots_5_io_uop_prs1 : _GEN_110 ? _slots_4_io_uop_prs1 : _GEN_94 ? _slots_3_io_uop_prs1 : _GEN_113 ? _slots_2_io_uop_prs1 : _GEN_44 ? _slots_1_io_uop_prs1 : _GEN_12987 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_1_prs2 = _GEN_596 ? _slots_39_io_uop_prs2 : _GEN_586 ? _slots_38_io_uop_prs2 : _GEN_599 ? _slots_37_io_uop_prs2 : _GEN_561 ? _slots_36_io_uop_prs2 : _GEN_547 ? _slots_35_io_uop_prs2 : _GEN_530 ? _slots_34_io_uop_prs2 : _GEN_516 ? _slots_33_io_uop_prs2 : _GEN_533 ? _slots_32_io_uop_prs2 : _GEN_491 ? _slots_31_io_uop_prs2 : _GEN_477 ? _slots_30_io_uop_prs2 : _GEN_460 ? _slots_29_io_uop_prs2 : _GEN_446 ? _slots_28_io_uop_prs2 : _GEN_463 ? _slots_27_io_uop_prs2 : _GEN_421 ? _slots_26_io_uop_prs2 : _GEN_407 ? _slots_25_io_uop_prs2 : _GEN_390 ? _slots_24_io_uop_prs2 : _GEN_376 ? _slots_23_io_uop_prs2 : _GEN_393 ? _slots_22_io_uop_prs2 : _GEN_351 ? _slots_21_io_uop_prs2 : _GEN_337 ? _slots_20_io_uop_prs2 : _GEN_320 ? _slots_19_io_uop_prs2 : _GEN_306 ? _slots_18_io_uop_prs2 : _GEN_323 ? _slots_17_io_uop_prs2 : _GEN_281 ? _slots_16_io_uop_prs2 : _GEN_267 ? _slots_15_io_uop_prs2 : _GEN_250 ? _slots_14_io_uop_prs2 : _GEN_236 ? _slots_13_io_uop_prs2 : _GEN_253 ? _slots_12_io_uop_prs2 : _GEN_211 ? _slots_11_io_uop_prs2 : _GEN_197 ? _slots_10_io_uop_prs2 : _GEN_180 ? _slots_9_io_uop_prs2 : _GEN_166 ? _slots_8_io_uop_prs2 : _GEN_183 ? _slots_7_io_uop_prs2 : _GEN_141 ? _slots_6_io_uop_prs2 : _GEN_127 ? _slots_5_io_uop_prs2 : _GEN_110 ? _slots_4_io_uop_prs2 : _GEN_94 ? _slots_3_io_uop_prs2 : _GEN_113 ? _slots_2_io_uop_prs2 : _GEN_44 ? _slots_1_io_uop_prs2 : _GEN_12987 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_1_bypassable = _GEN_596 ? _slots_39_io_uop_bypassable : _GEN_586 ? _slots_38_io_uop_bypassable : _GEN_599 ? _slots_37_io_uop_bypassable : _GEN_561 ? _slots_36_io_uop_bypassable : _GEN_547 ? _slots_35_io_uop_bypassable : _GEN_530 ? _slots_34_io_uop_bypassable : _GEN_516 ? _slots_33_io_uop_bypassable : _GEN_533 ? _slots_32_io_uop_bypassable : _GEN_491 ? _slots_31_io_uop_bypassable : _GEN_477 ? _slots_30_io_uop_bypassable : _GEN_460 ? _slots_29_io_uop_bypassable : _GEN_446 ? _slots_28_io_uop_bypassable : _GEN_463 ? _slots_27_io_uop_bypassable : _GEN_421 ? _slots_26_io_uop_bypassable : _GEN_407 ? _slots_25_io_uop_bypassable : _GEN_390 ? _slots_24_io_uop_bypassable : _GEN_376 ? _slots_23_io_uop_bypassable : _GEN_393 ? _slots_22_io_uop_bypassable : _GEN_351 ? _slots_21_io_uop_bypassable : _GEN_337 ? _slots_20_io_uop_bypassable : _GEN_320 ? _slots_19_io_uop_bypassable : _GEN_306 ? _slots_18_io_uop_bypassable : _GEN_323 ? _slots_17_io_uop_bypassable : _GEN_281 ? _slots_16_io_uop_bypassable : _GEN_267 ? _slots_15_io_uop_bypassable : _GEN_250 ? _slots_14_io_uop_bypassable : _GEN_236 ? _slots_13_io_uop_bypassable : _GEN_253 ? _slots_12_io_uop_bypassable : _GEN_211 ? _slots_11_io_uop_bypassable : _GEN_197 ? _slots_10_io_uop_bypassable : _GEN_180 ? _slots_9_io_uop_bypassable : _GEN_166 ? _slots_8_io_uop_bypassable : _GEN_183 ? _slots_7_io_uop_bypassable : _GEN_141 ? _slots_6_io_uop_bypassable : _GEN_127 ? _slots_5_io_uop_bypassable : _GEN_110 ? _slots_4_io_uop_bypassable : _GEN_94 ? _slots_3_io_uop_bypassable : _GEN_113 ? _slots_2_io_uop_bypassable : _GEN_44 ? _slots_1_io_uop_bypassable : _GEN_12987 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_1_mem_cmd = _GEN_596 ? _slots_39_io_uop_mem_cmd : _GEN_586 ? _slots_38_io_uop_mem_cmd : _GEN_599 ? _slots_37_io_uop_mem_cmd : _GEN_561 ? _slots_36_io_uop_mem_cmd : _GEN_547 ? _slots_35_io_uop_mem_cmd : _GEN_530 ? _slots_34_io_uop_mem_cmd : _GEN_516 ? _slots_33_io_uop_mem_cmd : _GEN_533 ? _slots_32_io_uop_mem_cmd : _GEN_491 ? _slots_31_io_uop_mem_cmd : _GEN_477 ? _slots_30_io_uop_mem_cmd : _GEN_460 ? _slots_29_io_uop_mem_cmd : _GEN_446 ? _slots_28_io_uop_mem_cmd : _GEN_463 ? _slots_27_io_uop_mem_cmd : _GEN_421 ? _slots_26_io_uop_mem_cmd : _GEN_407 ? _slots_25_io_uop_mem_cmd : _GEN_390 ? _slots_24_io_uop_mem_cmd : _GEN_376 ? _slots_23_io_uop_mem_cmd : _GEN_393 ? _slots_22_io_uop_mem_cmd : _GEN_351 ? _slots_21_io_uop_mem_cmd : _GEN_337 ? _slots_20_io_uop_mem_cmd : _GEN_320 ? _slots_19_io_uop_mem_cmd : _GEN_306 ? _slots_18_io_uop_mem_cmd : _GEN_323 ? _slots_17_io_uop_mem_cmd : _GEN_281 ? _slots_16_io_uop_mem_cmd : _GEN_267 ? _slots_15_io_uop_mem_cmd : _GEN_250 ? _slots_14_io_uop_mem_cmd : _GEN_236 ? _slots_13_io_uop_mem_cmd : _GEN_253 ? _slots_12_io_uop_mem_cmd : _GEN_211 ? _slots_11_io_uop_mem_cmd : _GEN_197 ? _slots_10_io_uop_mem_cmd : _GEN_180 ? _slots_9_io_uop_mem_cmd : _GEN_166 ? _slots_8_io_uop_mem_cmd : _GEN_183 ? _slots_7_io_uop_mem_cmd : _GEN_141 ? _slots_6_io_uop_mem_cmd : _GEN_127 ? _slots_5_io_uop_mem_cmd : _GEN_110 ? _slots_4_io_uop_mem_cmd : _GEN_94 ? _slots_3_io_uop_mem_cmd : _GEN_113 ? _slots_2_io_uop_mem_cmd : _GEN_44 ? _slots_1_io_uop_mem_cmd : _GEN_12987 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_1_is_amo = _GEN_596 ? _slots_39_io_uop_is_amo : _GEN_586 ? _slots_38_io_uop_is_amo : _GEN_599 ? _slots_37_io_uop_is_amo : _GEN_561 ? _slots_36_io_uop_is_amo : _GEN_547 ? _slots_35_io_uop_is_amo : _GEN_530 ? _slots_34_io_uop_is_amo : _GEN_516 ? _slots_33_io_uop_is_amo : _GEN_533 ? _slots_32_io_uop_is_amo : _GEN_491 ? _slots_31_io_uop_is_amo : _GEN_477 ? _slots_30_io_uop_is_amo : _GEN_460 ? _slots_29_io_uop_is_amo : _GEN_446 ? _slots_28_io_uop_is_amo : _GEN_463 ? _slots_27_io_uop_is_amo : _GEN_421 ? _slots_26_io_uop_is_amo : _GEN_407 ? _slots_25_io_uop_is_amo : _GEN_390 ? _slots_24_io_uop_is_amo : _GEN_376 ? _slots_23_io_uop_is_amo : _GEN_393 ? _slots_22_io_uop_is_amo : _GEN_351 ? _slots_21_io_uop_is_amo : _GEN_337 ? _slots_20_io_uop_is_amo : _GEN_320 ? _slots_19_io_uop_is_amo : _GEN_306 ? _slots_18_io_uop_is_amo : _GEN_323 ? _slots_17_io_uop_is_amo : _GEN_281 ? _slots_16_io_uop_is_amo : _GEN_267 ? _slots_15_io_uop_is_amo : _GEN_250 ? _slots_14_io_uop_is_amo : _GEN_236 ? _slots_13_io_uop_is_amo : _GEN_253 ? _slots_12_io_uop_is_amo : _GEN_211 ? _slots_11_io_uop_is_amo : _GEN_197 ? _slots_10_io_uop_is_amo : _GEN_180 ? _slots_9_io_uop_is_amo : _GEN_166 ? _slots_8_io_uop_is_amo : _GEN_183 ? _slots_7_io_uop_is_amo : _GEN_141 ? _slots_6_io_uop_is_amo : _GEN_127 ? _slots_5_io_uop_is_amo : _GEN_110 ? _slots_4_io_uop_is_amo : _GEN_94 ? _slots_3_io_uop_is_amo : _GEN_113 ? _slots_2_io_uop_is_amo : _GEN_44 ? _slots_1_io_uop_is_amo : _GEN_12987 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_1_uses_stq = _GEN_596 ? _slots_39_io_uop_uses_stq : _GEN_586 ? _slots_38_io_uop_uses_stq : _GEN_599 ? _slots_37_io_uop_uses_stq : _GEN_561 ? _slots_36_io_uop_uses_stq : _GEN_547 ? _slots_35_io_uop_uses_stq : _GEN_530 ? _slots_34_io_uop_uses_stq : _GEN_516 ? _slots_33_io_uop_uses_stq : _GEN_533 ? _slots_32_io_uop_uses_stq : _GEN_491 ? _slots_31_io_uop_uses_stq : _GEN_477 ? _slots_30_io_uop_uses_stq : _GEN_460 ? _slots_29_io_uop_uses_stq : _GEN_446 ? _slots_28_io_uop_uses_stq : _GEN_463 ? _slots_27_io_uop_uses_stq : _GEN_421 ? _slots_26_io_uop_uses_stq : _GEN_407 ? _slots_25_io_uop_uses_stq : _GEN_390 ? _slots_24_io_uop_uses_stq : _GEN_376 ? _slots_23_io_uop_uses_stq : _GEN_393 ? _slots_22_io_uop_uses_stq : _GEN_351 ? _slots_21_io_uop_uses_stq : _GEN_337 ? _slots_20_io_uop_uses_stq : _GEN_320 ? _slots_19_io_uop_uses_stq : _GEN_306 ? _slots_18_io_uop_uses_stq : _GEN_323 ? _slots_17_io_uop_uses_stq : _GEN_281 ? _slots_16_io_uop_uses_stq : _GEN_267 ? _slots_15_io_uop_uses_stq : _GEN_250 ? _slots_14_io_uop_uses_stq : _GEN_236 ? _slots_13_io_uop_uses_stq : _GEN_253 ? _slots_12_io_uop_uses_stq : _GEN_211 ? _slots_11_io_uop_uses_stq : _GEN_197 ? _slots_10_io_uop_uses_stq : _GEN_180 ? _slots_9_io_uop_uses_stq : _GEN_166 ? _slots_8_io_uop_uses_stq : _GEN_183 ? _slots_7_io_uop_uses_stq : _GEN_141 ? _slots_6_io_uop_uses_stq : _GEN_127 ? _slots_5_io_uop_uses_stq : _GEN_110 ? _slots_4_io_uop_uses_stq : _GEN_94 ? _slots_3_io_uop_uses_stq : _GEN_113 ? _slots_2_io_uop_uses_stq : _GEN_44 ? _slots_1_io_uop_uses_stq : _GEN_12987 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_1_ldst_val = _GEN_596 ? _slots_39_io_uop_ldst_val : _GEN_586 ? _slots_38_io_uop_ldst_val : _GEN_599 ? _slots_37_io_uop_ldst_val : _GEN_561 ? _slots_36_io_uop_ldst_val : _GEN_547 ? _slots_35_io_uop_ldst_val : _GEN_530 ? _slots_34_io_uop_ldst_val : _GEN_516 ? _slots_33_io_uop_ldst_val : _GEN_533 ? _slots_32_io_uop_ldst_val : _GEN_491 ? _slots_31_io_uop_ldst_val : _GEN_477 ? _slots_30_io_uop_ldst_val : _GEN_460 ? _slots_29_io_uop_ldst_val : _GEN_446 ? _slots_28_io_uop_ldst_val : _GEN_463 ? _slots_27_io_uop_ldst_val : _GEN_421 ? _slots_26_io_uop_ldst_val : _GEN_407 ? _slots_25_io_uop_ldst_val : _GEN_390 ? _slots_24_io_uop_ldst_val : _GEN_376 ? _slots_23_io_uop_ldst_val : _GEN_393 ? _slots_22_io_uop_ldst_val : _GEN_351 ? _slots_21_io_uop_ldst_val : _GEN_337 ? _slots_20_io_uop_ldst_val : _GEN_320 ? _slots_19_io_uop_ldst_val : _GEN_306 ? _slots_18_io_uop_ldst_val : _GEN_323 ? _slots_17_io_uop_ldst_val : _GEN_281 ? _slots_16_io_uop_ldst_val : _GEN_267 ? _slots_15_io_uop_ldst_val : _GEN_250 ? _slots_14_io_uop_ldst_val : _GEN_236 ? _slots_13_io_uop_ldst_val : _GEN_253 ? _slots_12_io_uop_ldst_val : _GEN_211 ? _slots_11_io_uop_ldst_val : _GEN_197 ? _slots_10_io_uop_ldst_val : _GEN_180 ? _slots_9_io_uop_ldst_val : _GEN_166 ? _slots_8_io_uop_ldst_val : _GEN_183 ? _slots_7_io_uop_ldst_val : _GEN_141 ? _slots_6_io_uop_ldst_val : _GEN_127 ? _slots_5_io_uop_ldst_val : _GEN_110 ? _slots_4_io_uop_ldst_val : _GEN_94 ? _slots_3_io_uop_ldst_val : _GEN_113 ? _slots_2_io_uop_ldst_val : _GEN_44 ? _slots_1_io_uop_ldst_val : _GEN_12987 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_1_dst_rtype = _GEN_596 ? _slots_39_io_uop_dst_rtype : _GEN_586 ? _slots_38_io_uop_dst_rtype : _GEN_599 ? _slots_37_io_uop_dst_rtype : _GEN_561 ? _slots_36_io_uop_dst_rtype : _GEN_547 ? _slots_35_io_uop_dst_rtype : _GEN_530 ? _slots_34_io_uop_dst_rtype : _GEN_516 ? _slots_33_io_uop_dst_rtype : _GEN_533 ? _slots_32_io_uop_dst_rtype : _GEN_491 ? _slots_31_io_uop_dst_rtype : _GEN_477 ? _slots_30_io_uop_dst_rtype : _GEN_460 ? _slots_29_io_uop_dst_rtype : _GEN_446 ? _slots_28_io_uop_dst_rtype : _GEN_463 ? _slots_27_io_uop_dst_rtype : _GEN_421 ? _slots_26_io_uop_dst_rtype : _GEN_407 ? _slots_25_io_uop_dst_rtype : _GEN_390 ? _slots_24_io_uop_dst_rtype : _GEN_376 ? _slots_23_io_uop_dst_rtype : _GEN_393 ? _slots_22_io_uop_dst_rtype : _GEN_351 ? _slots_21_io_uop_dst_rtype : _GEN_337 ? _slots_20_io_uop_dst_rtype : _GEN_320 ? _slots_19_io_uop_dst_rtype : _GEN_306 ? _slots_18_io_uop_dst_rtype : _GEN_323 ? _slots_17_io_uop_dst_rtype : _GEN_281 ? _slots_16_io_uop_dst_rtype : _GEN_267 ? _slots_15_io_uop_dst_rtype : _GEN_250 ? _slots_14_io_uop_dst_rtype : _GEN_236 ? _slots_13_io_uop_dst_rtype : _GEN_253 ? _slots_12_io_uop_dst_rtype : _GEN_211 ? _slots_11_io_uop_dst_rtype : _GEN_197 ? _slots_10_io_uop_dst_rtype : _GEN_180 ? _slots_9_io_uop_dst_rtype : _GEN_166 ? _slots_8_io_uop_dst_rtype : _GEN_183 ? _slots_7_io_uop_dst_rtype : _GEN_141 ? _slots_6_io_uop_dst_rtype : _GEN_127 ? _slots_5_io_uop_dst_rtype : _GEN_110 ? _slots_4_io_uop_dst_rtype : _GEN_94 ? _slots_3_io_uop_dst_rtype : _GEN_113 ? _slots_2_io_uop_dst_rtype : _GEN_44 ? _slots_1_io_uop_dst_rtype : _GEN_12987 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_1_lrs1_rtype = _GEN_596 ? _slots_39_io_uop_lrs1_rtype : _GEN_586 ? _slots_38_io_uop_lrs1_rtype : _GEN_599 ? _slots_37_io_uop_lrs1_rtype : _GEN_561 ? _slots_36_io_uop_lrs1_rtype : _GEN_547 ? _slots_35_io_uop_lrs1_rtype : _GEN_530 ? _slots_34_io_uop_lrs1_rtype : _GEN_516 ? _slots_33_io_uop_lrs1_rtype : _GEN_533 ? _slots_32_io_uop_lrs1_rtype : _GEN_491 ? _slots_31_io_uop_lrs1_rtype : _GEN_477 ? _slots_30_io_uop_lrs1_rtype : _GEN_460 ? _slots_29_io_uop_lrs1_rtype : _GEN_446 ? _slots_28_io_uop_lrs1_rtype : _GEN_463 ? _slots_27_io_uop_lrs1_rtype : _GEN_421 ? _slots_26_io_uop_lrs1_rtype : _GEN_407 ? _slots_25_io_uop_lrs1_rtype : _GEN_390 ? _slots_24_io_uop_lrs1_rtype : _GEN_376 ? _slots_23_io_uop_lrs1_rtype : _GEN_393 ? _slots_22_io_uop_lrs1_rtype : _GEN_351 ? _slots_21_io_uop_lrs1_rtype : _GEN_337 ? _slots_20_io_uop_lrs1_rtype : _GEN_320 ? _slots_19_io_uop_lrs1_rtype : _GEN_306 ? _slots_18_io_uop_lrs1_rtype : _GEN_323 ? _slots_17_io_uop_lrs1_rtype : _GEN_281 ? _slots_16_io_uop_lrs1_rtype : _GEN_267 ? _slots_15_io_uop_lrs1_rtype : _GEN_250 ? _slots_14_io_uop_lrs1_rtype : _GEN_236 ? _slots_13_io_uop_lrs1_rtype : _GEN_253 ? _slots_12_io_uop_lrs1_rtype : _GEN_211 ? _slots_11_io_uop_lrs1_rtype : _GEN_197 ? _slots_10_io_uop_lrs1_rtype : _GEN_180 ? _slots_9_io_uop_lrs1_rtype : _GEN_166 ? _slots_8_io_uop_lrs1_rtype : _GEN_183 ? _slots_7_io_uop_lrs1_rtype : _GEN_141 ? _slots_6_io_uop_lrs1_rtype : _GEN_127 ? _slots_5_io_uop_lrs1_rtype : _GEN_110 ? _slots_4_io_uop_lrs1_rtype : _GEN_94 ? _slots_3_io_uop_lrs1_rtype : _GEN_113 ? _slots_2_io_uop_lrs1_rtype : _GEN_44 ? _slots_1_io_uop_lrs1_rtype : _GEN_12987 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_1_lrs2_rtype = _GEN_596 ? _slots_39_io_uop_lrs2_rtype : _GEN_586 ? _slots_38_io_uop_lrs2_rtype : _GEN_599 ? _slots_37_io_uop_lrs2_rtype : _GEN_561 ? _slots_36_io_uop_lrs2_rtype : _GEN_547 ? _slots_35_io_uop_lrs2_rtype : _GEN_530 ? _slots_34_io_uop_lrs2_rtype : _GEN_516 ? _slots_33_io_uop_lrs2_rtype : _GEN_533 ? _slots_32_io_uop_lrs2_rtype : _GEN_491 ? _slots_31_io_uop_lrs2_rtype : _GEN_477 ? _slots_30_io_uop_lrs2_rtype : _GEN_460 ? _slots_29_io_uop_lrs2_rtype : _GEN_446 ? _slots_28_io_uop_lrs2_rtype : _GEN_463 ? _slots_27_io_uop_lrs2_rtype : _GEN_421 ? _slots_26_io_uop_lrs2_rtype : _GEN_407 ? _slots_25_io_uop_lrs2_rtype : _GEN_390 ? _slots_24_io_uop_lrs2_rtype : _GEN_376 ? _slots_23_io_uop_lrs2_rtype : _GEN_393 ? _slots_22_io_uop_lrs2_rtype : _GEN_351 ? _slots_21_io_uop_lrs2_rtype : _GEN_337 ? _slots_20_io_uop_lrs2_rtype : _GEN_320 ? _slots_19_io_uop_lrs2_rtype : _GEN_306 ? _slots_18_io_uop_lrs2_rtype : _GEN_323 ? _slots_17_io_uop_lrs2_rtype : _GEN_281 ? _slots_16_io_uop_lrs2_rtype : _GEN_267 ? _slots_15_io_uop_lrs2_rtype : _GEN_250 ? _slots_14_io_uop_lrs2_rtype : _GEN_236 ? _slots_13_io_uop_lrs2_rtype : _GEN_253 ? _slots_12_io_uop_lrs2_rtype : _GEN_211 ? _slots_11_io_uop_lrs2_rtype : _GEN_197 ? _slots_10_io_uop_lrs2_rtype : _GEN_180 ? _slots_9_io_uop_lrs2_rtype : _GEN_166 ? _slots_8_io_uop_lrs2_rtype : _GEN_183 ? _slots_7_io_uop_lrs2_rtype : _GEN_141 ? _slots_6_io_uop_lrs2_rtype : _GEN_127 ? _slots_5_io_uop_lrs2_rtype : _GEN_110 ? _slots_4_io_uop_lrs2_rtype : _GEN_94 ? _slots_3_io_uop_lrs2_rtype : _GEN_113 ? _slots_2_io_uop_lrs2_rtype : _GEN_44 ? _slots_1_io_uop_lrs2_rtype : _GEN_12987 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_2_uopc = _GEN_595 ? _slots_39_io_uop_uopc : _GEN_584 ? _slots_38_io_uop_uopc : _GEN_598 ? _slots_37_io_uop_uopc : _GEN_559 ? _slots_36_io_uop_uopc : _GEN_545 ? _slots_35_io_uop_uopc : _GEN_528 ? _slots_34_io_uop_uopc : _GEN_514 ? _slots_33_io_uop_uopc : _GEN_532 ? _slots_32_io_uop_uopc : _GEN_489 ? _slots_31_io_uop_uopc : _GEN_475 ? _slots_30_io_uop_uopc : _GEN_458 ? _slots_29_io_uop_uopc : _GEN_444 ? _slots_28_io_uop_uopc : _GEN_462 ? _slots_27_io_uop_uopc : _GEN_419 ? _slots_26_io_uop_uopc : _GEN_405 ? _slots_25_io_uop_uopc : _GEN_388 ? _slots_24_io_uop_uopc : _GEN_374 ? _slots_23_io_uop_uopc : _GEN_392 ? _slots_22_io_uop_uopc : _GEN_349 ? _slots_21_io_uop_uopc : _GEN_335 ? _slots_20_io_uop_uopc : _GEN_318 ? _slots_19_io_uop_uopc : _GEN_304 ? _slots_18_io_uop_uopc : _GEN_322 ? _slots_17_io_uop_uopc : _GEN_279 ? _slots_16_io_uop_uopc : _GEN_265 ? _slots_15_io_uop_uopc : _GEN_248 ? _slots_14_io_uop_uopc : _GEN_234 ? _slots_13_io_uop_uopc : _GEN_252 ? _slots_12_io_uop_uopc : _GEN_209 ? _slots_11_io_uop_uopc : _GEN_195 ? _slots_10_io_uop_uopc : _GEN_178 ? _slots_9_io_uop_uopc : _GEN_164 ? _slots_8_io_uop_uopc : _GEN_182 ? _slots_7_io_uop_uopc : _GEN_139 ? _slots_6_io_uop_uopc : _GEN_125 ? _slots_5_io_uop_uopc : _GEN_108 ? _slots_4_io_uop_uopc : _GEN_90 ? _slots_3_io_uop_uopc : _GEN_112 ? _slots_2_io_uop_uopc : _GEN_40 ? _slots_1_io_uop_uopc : _GEN_13068 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_2_is_rvc = _GEN_595 ? _slots_39_io_uop_is_rvc : _GEN_584 ? _slots_38_io_uop_is_rvc : _GEN_598 ? _slots_37_io_uop_is_rvc : _GEN_559 ? _slots_36_io_uop_is_rvc : _GEN_545 ? _slots_35_io_uop_is_rvc : _GEN_528 ? _slots_34_io_uop_is_rvc : _GEN_514 ? _slots_33_io_uop_is_rvc : _GEN_532 ? _slots_32_io_uop_is_rvc : _GEN_489 ? _slots_31_io_uop_is_rvc : _GEN_475 ? _slots_30_io_uop_is_rvc : _GEN_458 ? _slots_29_io_uop_is_rvc : _GEN_444 ? _slots_28_io_uop_is_rvc : _GEN_462 ? _slots_27_io_uop_is_rvc : _GEN_419 ? _slots_26_io_uop_is_rvc : _GEN_405 ? _slots_25_io_uop_is_rvc : _GEN_388 ? _slots_24_io_uop_is_rvc : _GEN_374 ? _slots_23_io_uop_is_rvc : _GEN_392 ? _slots_22_io_uop_is_rvc : _GEN_349 ? _slots_21_io_uop_is_rvc : _GEN_335 ? _slots_20_io_uop_is_rvc : _GEN_318 ? _slots_19_io_uop_is_rvc : _GEN_304 ? _slots_18_io_uop_is_rvc : _GEN_322 ? _slots_17_io_uop_is_rvc : _GEN_279 ? _slots_16_io_uop_is_rvc : _GEN_265 ? _slots_15_io_uop_is_rvc : _GEN_248 ? _slots_14_io_uop_is_rvc : _GEN_234 ? _slots_13_io_uop_is_rvc : _GEN_252 ? _slots_12_io_uop_is_rvc : _GEN_209 ? _slots_11_io_uop_is_rvc : _GEN_195 ? _slots_10_io_uop_is_rvc : _GEN_178 ? _slots_9_io_uop_is_rvc : _GEN_164 ? _slots_8_io_uop_is_rvc : _GEN_182 ? _slots_7_io_uop_is_rvc : _GEN_139 ? _slots_6_io_uop_is_rvc : _GEN_125 ? _slots_5_io_uop_is_rvc : _GEN_108 ? _slots_4_io_uop_is_rvc : _GEN_90 ? _slots_3_io_uop_is_rvc : _GEN_112 ? _slots_2_io_uop_is_rvc : _GEN_40 ? _slots_1_io_uop_is_rvc : _GEN_13068 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_2_fu_code = _GEN_595 ? _slots_39_io_uop_fu_code : _GEN_584 ? _slots_38_io_uop_fu_code : _GEN_598 ? _slots_37_io_uop_fu_code : _GEN_559 ? _slots_36_io_uop_fu_code : _GEN_545 ? _slots_35_io_uop_fu_code : _GEN_528 ? _slots_34_io_uop_fu_code : _GEN_514 ? _slots_33_io_uop_fu_code : _GEN_532 ? _slots_32_io_uop_fu_code : _GEN_489 ? _slots_31_io_uop_fu_code : _GEN_475 ? _slots_30_io_uop_fu_code : _GEN_458 ? _slots_29_io_uop_fu_code : _GEN_444 ? _slots_28_io_uop_fu_code : _GEN_462 ? _slots_27_io_uop_fu_code : _GEN_419 ? _slots_26_io_uop_fu_code : _GEN_405 ? _slots_25_io_uop_fu_code : _GEN_388 ? _slots_24_io_uop_fu_code : _GEN_374 ? _slots_23_io_uop_fu_code : _GEN_392 ? _slots_22_io_uop_fu_code : _GEN_349 ? _slots_21_io_uop_fu_code : _GEN_335 ? _slots_20_io_uop_fu_code : _GEN_318 ? _slots_19_io_uop_fu_code : _GEN_304 ? _slots_18_io_uop_fu_code : _GEN_322 ? _slots_17_io_uop_fu_code : _GEN_279 ? _slots_16_io_uop_fu_code : _GEN_265 ? _slots_15_io_uop_fu_code : _GEN_248 ? _slots_14_io_uop_fu_code : _GEN_234 ? _slots_13_io_uop_fu_code : _GEN_252 ? _slots_12_io_uop_fu_code : _GEN_209 ? _slots_11_io_uop_fu_code : _GEN_195 ? _slots_10_io_uop_fu_code : _GEN_178 ? _slots_9_io_uop_fu_code : _GEN_164 ? _slots_8_io_uop_fu_code : _GEN_182 ? _slots_7_io_uop_fu_code : _GEN_139 ? _slots_6_io_uop_fu_code : _GEN_125 ? _slots_5_io_uop_fu_code : _GEN_108 ? _slots_4_io_uop_fu_code : _GEN_90 ? _slots_3_io_uop_fu_code : _GEN_112 ? _slots_2_io_uop_fu_code : _GEN_40 ? _slots_1_io_uop_fu_code : _GEN_13068 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_2_iw_p1_poisoned = _GEN_595 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_584 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_598 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_559 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_545 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_528 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_514 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_532 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_489 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_475 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_458 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_444 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_462 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_419 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_405 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_388 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_374 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_392 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_349 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_335 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_318 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_304 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_322 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_279 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_265 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_248 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_234 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_252 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_209 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_195 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_178 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_164 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_182 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_139 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_125 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_108 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_90 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_112 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_40 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_13068 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_2_iw_p2_poisoned = _GEN_595 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_584 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_598 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_559 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_545 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_528 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_514 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_532 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_489 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_475 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_458 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_444 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_462 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_419 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_405 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_388 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_374 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_392 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_349 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_335 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_318 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_304 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_322 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_279 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_265 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_248 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_234 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_252 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_209 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_195 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_178 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_164 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_182 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_139 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_125 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_108 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_90 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_112 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_40 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_13068 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_2_is_br = _GEN_595 ? _slots_39_io_uop_is_br : _GEN_584 ? _slots_38_io_uop_is_br : _GEN_598 ? _slots_37_io_uop_is_br : _GEN_559 ? _slots_36_io_uop_is_br : _GEN_545 ? _slots_35_io_uop_is_br : _GEN_528 ? _slots_34_io_uop_is_br : _GEN_514 ? _slots_33_io_uop_is_br : _GEN_532 ? _slots_32_io_uop_is_br : _GEN_489 ? _slots_31_io_uop_is_br : _GEN_475 ? _slots_30_io_uop_is_br : _GEN_458 ? _slots_29_io_uop_is_br : _GEN_444 ? _slots_28_io_uop_is_br : _GEN_462 ? _slots_27_io_uop_is_br : _GEN_419 ? _slots_26_io_uop_is_br : _GEN_405 ? _slots_25_io_uop_is_br : _GEN_388 ? _slots_24_io_uop_is_br : _GEN_374 ? _slots_23_io_uop_is_br : _GEN_392 ? _slots_22_io_uop_is_br : _GEN_349 ? _slots_21_io_uop_is_br : _GEN_335 ? _slots_20_io_uop_is_br : _GEN_318 ? _slots_19_io_uop_is_br : _GEN_304 ? _slots_18_io_uop_is_br : _GEN_322 ? _slots_17_io_uop_is_br : _GEN_279 ? _slots_16_io_uop_is_br : _GEN_265 ? _slots_15_io_uop_is_br : _GEN_248 ? _slots_14_io_uop_is_br : _GEN_234 ? _slots_13_io_uop_is_br : _GEN_252 ? _slots_12_io_uop_is_br : _GEN_209 ? _slots_11_io_uop_is_br : _GEN_195 ? _slots_10_io_uop_is_br : _GEN_178 ? _slots_9_io_uop_is_br : _GEN_164 ? _slots_8_io_uop_is_br : _GEN_182 ? _slots_7_io_uop_is_br : _GEN_139 ? _slots_6_io_uop_is_br : _GEN_125 ? _slots_5_io_uop_is_br : _GEN_108 ? _slots_4_io_uop_is_br : _GEN_90 ? _slots_3_io_uop_is_br : _GEN_112 ? _slots_2_io_uop_is_br : _GEN_40 ? _slots_1_io_uop_is_br : _GEN_13068 & _slots_0_io_uop_is_br;
  assign io_iss_uops_2_is_jalr = _GEN_595 ? _slots_39_io_uop_is_jalr : _GEN_584 ? _slots_38_io_uop_is_jalr : _GEN_598 ? _slots_37_io_uop_is_jalr : _GEN_559 ? _slots_36_io_uop_is_jalr : _GEN_545 ? _slots_35_io_uop_is_jalr : _GEN_528 ? _slots_34_io_uop_is_jalr : _GEN_514 ? _slots_33_io_uop_is_jalr : _GEN_532 ? _slots_32_io_uop_is_jalr : _GEN_489 ? _slots_31_io_uop_is_jalr : _GEN_475 ? _slots_30_io_uop_is_jalr : _GEN_458 ? _slots_29_io_uop_is_jalr : _GEN_444 ? _slots_28_io_uop_is_jalr : _GEN_462 ? _slots_27_io_uop_is_jalr : _GEN_419 ? _slots_26_io_uop_is_jalr : _GEN_405 ? _slots_25_io_uop_is_jalr : _GEN_388 ? _slots_24_io_uop_is_jalr : _GEN_374 ? _slots_23_io_uop_is_jalr : _GEN_392 ? _slots_22_io_uop_is_jalr : _GEN_349 ? _slots_21_io_uop_is_jalr : _GEN_335 ? _slots_20_io_uop_is_jalr : _GEN_318 ? _slots_19_io_uop_is_jalr : _GEN_304 ? _slots_18_io_uop_is_jalr : _GEN_322 ? _slots_17_io_uop_is_jalr : _GEN_279 ? _slots_16_io_uop_is_jalr : _GEN_265 ? _slots_15_io_uop_is_jalr : _GEN_248 ? _slots_14_io_uop_is_jalr : _GEN_234 ? _slots_13_io_uop_is_jalr : _GEN_252 ? _slots_12_io_uop_is_jalr : _GEN_209 ? _slots_11_io_uop_is_jalr : _GEN_195 ? _slots_10_io_uop_is_jalr : _GEN_178 ? _slots_9_io_uop_is_jalr : _GEN_164 ? _slots_8_io_uop_is_jalr : _GEN_182 ? _slots_7_io_uop_is_jalr : _GEN_139 ? _slots_6_io_uop_is_jalr : _GEN_125 ? _slots_5_io_uop_is_jalr : _GEN_108 ? _slots_4_io_uop_is_jalr : _GEN_90 ? _slots_3_io_uop_is_jalr : _GEN_112 ? _slots_2_io_uop_is_jalr : _GEN_40 ? _slots_1_io_uop_is_jalr : _GEN_13068 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_2_is_jal = _GEN_595 ? _slots_39_io_uop_is_jal : _GEN_584 ? _slots_38_io_uop_is_jal : _GEN_598 ? _slots_37_io_uop_is_jal : _GEN_559 ? _slots_36_io_uop_is_jal : _GEN_545 ? _slots_35_io_uop_is_jal : _GEN_528 ? _slots_34_io_uop_is_jal : _GEN_514 ? _slots_33_io_uop_is_jal : _GEN_532 ? _slots_32_io_uop_is_jal : _GEN_489 ? _slots_31_io_uop_is_jal : _GEN_475 ? _slots_30_io_uop_is_jal : _GEN_458 ? _slots_29_io_uop_is_jal : _GEN_444 ? _slots_28_io_uop_is_jal : _GEN_462 ? _slots_27_io_uop_is_jal : _GEN_419 ? _slots_26_io_uop_is_jal : _GEN_405 ? _slots_25_io_uop_is_jal : _GEN_388 ? _slots_24_io_uop_is_jal : _GEN_374 ? _slots_23_io_uop_is_jal : _GEN_392 ? _slots_22_io_uop_is_jal : _GEN_349 ? _slots_21_io_uop_is_jal : _GEN_335 ? _slots_20_io_uop_is_jal : _GEN_318 ? _slots_19_io_uop_is_jal : _GEN_304 ? _slots_18_io_uop_is_jal : _GEN_322 ? _slots_17_io_uop_is_jal : _GEN_279 ? _slots_16_io_uop_is_jal : _GEN_265 ? _slots_15_io_uop_is_jal : _GEN_248 ? _slots_14_io_uop_is_jal : _GEN_234 ? _slots_13_io_uop_is_jal : _GEN_252 ? _slots_12_io_uop_is_jal : _GEN_209 ? _slots_11_io_uop_is_jal : _GEN_195 ? _slots_10_io_uop_is_jal : _GEN_178 ? _slots_9_io_uop_is_jal : _GEN_164 ? _slots_8_io_uop_is_jal : _GEN_182 ? _slots_7_io_uop_is_jal : _GEN_139 ? _slots_6_io_uop_is_jal : _GEN_125 ? _slots_5_io_uop_is_jal : _GEN_108 ? _slots_4_io_uop_is_jal : _GEN_90 ? _slots_3_io_uop_is_jal : _GEN_112 ? _slots_2_io_uop_is_jal : _GEN_40 ? _slots_1_io_uop_is_jal : _GEN_13068 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_2_is_sfb = _GEN_595 ? _slots_39_io_uop_is_sfb : _GEN_584 ? _slots_38_io_uop_is_sfb : _GEN_598 ? _slots_37_io_uop_is_sfb : _GEN_559 ? _slots_36_io_uop_is_sfb : _GEN_545 ? _slots_35_io_uop_is_sfb : _GEN_528 ? _slots_34_io_uop_is_sfb : _GEN_514 ? _slots_33_io_uop_is_sfb : _GEN_532 ? _slots_32_io_uop_is_sfb : _GEN_489 ? _slots_31_io_uop_is_sfb : _GEN_475 ? _slots_30_io_uop_is_sfb : _GEN_458 ? _slots_29_io_uop_is_sfb : _GEN_444 ? _slots_28_io_uop_is_sfb : _GEN_462 ? _slots_27_io_uop_is_sfb : _GEN_419 ? _slots_26_io_uop_is_sfb : _GEN_405 ? _slots_25_io_uop_is_sfb : _GEN_388 ? _slots_24_io_uop_is_sfb : _GEN_374 ? _slots_23_io_uop_is_sfb : _GEN_392 ? _slots_22_io_uop_is_sfb : _GEN_349 ? _slots_21_io_uop_is_sfb : _GEN_335 ? _slots_20_io_uop_is_sfb : _GEN_318 ? _slots_19_io_uop_is_sfb : _GEN_304 ? _slots_18_io_uop_is_sfb : _GEN_322 ? _slots_17_io_uop_is_sfb : _GEN_279 ? _slots_16_io_uop_is_sfb : _GEN_265 ? _slots_15_io_uop_is_sfb : _GEN_248 ? _slots_14_io_uop_is_sfb : _GEN_234 ? _slots_13_io_uop_is_sfb : _GEN_252 ? _slots_12_io_uop_is_sfb : _GEN_209 ? _slots_11_io_uop_is_sfb : _GEN_195 ? _slots_10_io_uop_is_sfb : _GEN_178 ? _slots_9_io_uop_is_sfb : _GEN_164 ? _slots_8_io_uop_is_sfb : _GEN_182 ? _slots_7_io_uop_is_sfb : _GEN_139 ? _slots_6_io_uop_is_sfb : _GEN_125 ? _slots_5_io_uop_is_sfb : _GEN_108 ? _slots_4_io_uop_is_sfb : _GEN_90 ? _slots_3_io_uop_is_sfb : _GEN_112 ? _slots_2_io_uop_is_sfb : _GEN_40 ? _slots_1_io_uop_is_sfb : _GEN_13068 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_2_br_mask = _GEN_595 ? _slots_39_io_uop_br_mask : _GEN_584 ? _slots_38_io_uop_br_mask : _GEN_598 ? _slots_37_io_uop_br_mask : _GEN_559 ? _slots_36_io_uop_br_mask : _GEN_545 ? _slots_35_io_uop_br_mask : _GEN_528 ? _slots_34_io_uop_br_mask : _GEN_514 ? _slots_33_io_uop_br_mask : _GEN_532 ? _slots_32_io_uop_br_mask : _GEN_489 ? _slots_31_io_uop_br_mask : _GEN_475 ? _slots_30_io_uop_br_mask : _GEN_458 ? _slots_29_io_uop_br_mask : _GEN_444 ? _slots_28_io_uop_br_mask : _GEN_462 ? _slots_27_io_uop_br_mask : _GEN_419 ? _slots_26_io_uop_br_mask : _GEN_405 ? _slots_25_io_uop_br_mask : _GEN_388 ? _slots_24_io_uop_br_mask : _GEN_374 ? _slots_23_io_uop_br_mask : _GEN_392 ? _slots_22_io_uop_br_mask : _GEN_349 ? _slots_21_io_uop_br_mask : _GEN_335 ? _slots_20_io_uop_br_mask : _GEN_318 ? _slots_19_io_uop_br_mask : _GEN_304 ? _slots_18_io_uop_br_mask : _GEN_322 ? _slots_17_io_uop_br_mask : _GEN_279 ? _slots_16_io_uop_br_mask : _GEN_265 ? _slots_15_io_uop_br_mask : _GEN_248 ? _slots_14_io_uop_br_mask : _GEN_234 ? _slots_13_io_uop_br_mask : _GEN_252 ? _slots_12_io_uop_br_mask : _GEN_209 ? _slots_11_io_uop_br_mask : _GEN_195 ? _slots_10_io_uop_br_mask : _GEN_178 ? _slots_9_io_uop_br_mask : _GEN_164 ? _slots_8_io_uop_br_mask : _GEN_182 ? _slots_7_io_uop_br_mask : _GEN_139 ? _slots_6_io_uop_br_mask : _GEN_125 ? _slots_5_io_uop_br_mask : _GEN_108 ? _slots_4_io_uop_br_mask : _GEN_90 ? _slots_3_io_uop_br_mask : _GEN_112 ? _slots_2_io_uop_br_mask : _GEN_40 ? _slots_1_io_uop_br_mask : _GEN_13068 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_2_br_tag = _GEN_595 ? _slots_39_io_uop_br_tag : _GEN_584 ? _slots_38_io_uop_br_tag : _GEN_598 ? _slots_37_io_uop_br_tag : _GEN_559 ? _slots_36_io_uop_br_tag : _GEN_545 ? _slots_35_io_uop_br_tag : _GEN_528 ? _slots_34_io_uop_br_tag : _GEN_514 ? _slots_33_io_uop_br_tag : _GEN_532 ? _slots_32_io_uop_br_tag : _GEN_489 ? _slots_31_io_uop_br_tag : _GEN_475 ? _slots_30_io_uop_br_tag : _GEN_458 ? _slots_29_io_uop_br_tag : _GEN_444 ? _slots_28_io_uop_br_tag : _GEN_462 ? _slots_27_io_uop_br_tag : _GEN_419 ? _slots_26_io_uop_br_tag : _GEN_405 ? _slots_25_io_uop_br_tag : _GEN_388 ? _slots_24_io_uop_br_tag : _GEN_374 ? _slots_23_io_uop_br_tag : _GEN_392 ? _slots_22_io_uop_br_tag : _GEN_349 ? _slots_21_io_uop_br_tag : _GEN_335 ? _slots_20_io_uop_br_tag : _GEN_318 ? _slots_19_io_uop_br_tag : _GEN_304 ? _slots_18_io_uop_br_tag : _GEN_322 ? _slots_17_io_uop_br_tag : _GEN_279 ? _slots_16_io_uop_br_tag : _GEN_265 ? _slots_15_io_uop_br_tag : _GEN_248 ? _slots_14_io_uop_br_tag : _GEN_234 ? _slots_13_io_uop_br_tag : _GEN_252 ? _slots_12_io_uop_br_tag : _GEN_209 ? _slots_11_io_uop_br_tag : _GEN_195 ? _slots_10_io_uop_br_tag : _GEN_178 ? _slots_9_io_uop_br_tag : _GEN_164 ? _slots_8_io_uop_br_tag : _GEN_182 ? _slots_7_io_uop_br_tag : _GEN_139 ? _slots_6_io_uop_br_tag : _GEN_125 ? _slots_5_io_uop_br_tag : _GEN_108 ? _slots_4_io_uop_br_tag : _GEN_90 ? _slots_3_io_uop_br_tag : _GEN_112 ? _slots_2_io_uop_br_tag : _GEN_40 ? _slots_1_io_uop_br_tag : _GEN_13068 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_2_ftq_idx = _GEN_595 ? _slots_39_io_uop_ftq_idx : _GEN_584 ? _slots_38_io_uop_ftq_idx : _GEN_598 ? _slots_37_io_uop_ftq_idx : _GEN_559 ? _slots_36_io_uop_ftq_idx : _GEN_545 ? _slots_35_io_uop_ftq_idx : _GEN_528 ? _slots_34_io_uop_ftq_idx : _GEN_514 ? _slots_33_io_uop_ftq_idx : _GEN_532 ? _slots_32_io_uop_ftq_idx : _GEN_489 ? _slots_31_io_uop_ftq_idx : _GEN_475 ? _slots_30_io_uop_ftq_idx : _GEN_458 ? _slots_29_io_uop_ftq_idx : _GEN_444 ? _slots_28_io_uop_ftq_idx : _GEN_462 ? _slots_27_io_uop_ftq_idx : _GEN_419 ? _slots_26_io_uop_ftq_idx : _GEN_405 ? _slots_25_io_uop_ftq_idx : _GEN_388 ? _slots_24_io_uop_ftq_idx : _GEN_374 ? _slots_23_io_uop_ftq_idx : _GEN_392 ? _slots_22_io_uop_ftq_idx : _GEN_349 ? _slots_21_io_uop_ftq_idx : _GEN_335 ? _slots_20_io_uop_ftq_idx : _GEN_318 ? _slots_19_io_uop_ftq_idx : _GEN_304 ? _slots_18_io_uop_ftq_idx : _GEN_322 ? _slots_17_io_uop_ftq_idx : _GEN_279 ? _slots_16_io_uop_ftq_idx : _GEN_265 ? _slots_15_io_uop_ftq_idx : _GEN_248 ? _slots_14_io_uop_ftq_idx : _GEN_234 ? _slots_13_io_uop_ftq_idx : _GEN_252 ? _slots_12_io_uop_ftq_idx : _GEN_209 ? _slots_11_io_uop_ftq_idx : _GEN_195 ? _slots_10_io_uop_ftq_idx : _GEN_178 ? _slots_9_io_uop_ftq_idx : _GEN_164 ? _slots_8_io_uop_ftq_idx : _GEN_182 ? _slots_7_io_uop_ftq_idx : _GEN_139 ? _slots_6_io_uop_ftq_idx : _GEN_125 ? _slots_5_io_uop_ftq_idx : _GEN_108 ? _slots_4_io_uop_ftq_idx : _GEN_90 ? _slots_3_io_uop_ftq_idx : _GEN_112 ? _slots_2_io_uop_ftq_idx : _GEN_40 ? _slots_1_io_uop_ftq_idx : _GEN_13068 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_2_edge_inst = _GEN_595 ? _slots_39_io_uop_edge_inst : _GEN_584 ? _slots_38_io_uop_edge_inst : _GEN_598 ? _slots_37_io_uop_edge_inst : _GEN_559 ? _slots_36_io_uop_edge_inst : _GEN_545 ? _slots_35_io_uop_edge_inst : _GEN_528 ? _slots_34_io_uop_edge_inst : _GEN_514 ? _slots_33_io_uop_edge_inst : _GEN_532 ? _slots_32_io_uop_edge_inst : _GEN_489 ? _slots_31_io_uop_edge_inst : _GEN_475 ? _slots_30_io_uop_edge_inst : _GEN_458 ? _slots_29_io_uop_edge_inst : _GEN_444 ? _slots_28_io_uop_edge_inst : _GEN_462 ? _slots_27_io_uop_edge_inst : _GEN_419 ? _slots_26_io_uop_edge_inst : _GEN_405 ? _slots_25_io_uop_edge_inst : _GEN_388 ? _slots_24_io_uop_edge_inst : _GEN_374 ? _slots_23_io_uop_edge_inst : _GEN_392 ? _slots_22_io_uop_edge_inst : _GEN_349 ? _slots_21_io_uop_edge_inst : _GEN_335 ? _slots_20_io_uop_edge_inst : _GEN_318 ? _slots_19_io_uop_edge_inst : _GEN_304 ? _slots_18_io_uop_edge_inst : _GEN_322 ? _slots_17_io_uop_edge_inst : _GEN_279 ? _slots_16_io_uop_edge_inst : _GEN_265 ? _slots_15_io_uop_edge_inst : _GEN_248 ? _slots_14_io_uop_edge_inst : _GEN_234 ? _slots_13_io_uop_edge_inst : _GEN_252 ? _slots_12_io_uop_edge_inst : _GEN_209 ? _slots_11_io_uop_edge_inst : _GEN_195 ? _slots_10_io_uop_edge_inst : _GEN_178 ? _slots_9_io_uop_edge_inst : _GEN_164 ? _slots_8_io_uop_edge_inst : _GEN_182 ? _slots_7_io_uop_edge_inst : _GEN_139 ? _slots_6_io_uop_edge_inst : _GEN_125 ? _slots_5_io_uop_edge_inst : _GEN_108 ? _slots_4_io_uop_edge_inst : _GEN_90 ? _slots_3_io_uop_edge_inst : _GEN_112 ? _slots_2_io_uop_edge_inst : _GEN_40 ? _slots_1_io_uop_edge_inst : _GEN_13068 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_2_pc_lob = _GEN_595 ? _slots_39_io_uop_pc_lob : _GEN_584 ? _slots_38_io_uop_pc_lob : _GEN_598 ? _slots_37_io_uop_pc_lob : _GEN_559 ? _slots_36_io_uop_pc_lob : _GEN_545 ? _slots_35_io_uop_pc_lob : _GEN_528 ? _slots_34_io_uop_pc_lob : _GEN_514 ? _slots_33_io_uop_pc_lob : _GEN_532 ? _slots_32_io_uop_pc_lob : _GEN_489 ? _slots_31_io_uop_pc_lob : _GEN_475 ? _slots_30_io_uop_pc_lob : _GEN_458 ? _slots_29_io_uop_pc_lob : _GEN_444 ? _slots_28_io_uop_pc_lob : _GEN_462 ? _slots_27_io_uop_pc_lob : _GEN_419 ? _slots_26_io_uop_pc_lob : _GEN_405 ? _slots_25_io_uop_pc_lob : _GEN_388 ? _slots_24_io_uop_pc_lob : _GEN_374 ? _slots_23_io_uop_pc_lob : _GEN_392 ? _slots_22_io_uop_pc_lob : _GEN_349 ? _slots_21_io_uop_pc_lob : _GEN_335 ? _slots_20_io_uop_pc_lob : _GEN_318 ? _slots_19_io_uop_pc_lob : _GEN_304 ? _slots_18_io_uop_pc_lob : _GEN_322 ? _slots_17_io_uop_pc_lob : _GEN_279 ? _slots_16_io_uop_pc_lob : _GEN_265 ? _slots_15_io_uop_pc_lob : _GEN_248 ? _slots_14_io_uop_pc_lob : _GEN_234 ? _slots_13_io_uop_pc_lob : _GEN_252 ? _slots_12_io_uop_pc_lob : _GEN_209 ? _slots_11_io_uop_pc_lob : _GEN_195 ? _slots_10_io_uop_pc_lob : _GEN_178 ? _slots_9_io_uop_pc_lob : _GEN_164 ? _slots_8_io_uop_pc_lob : _GEN_182 ? _slots_7_io_uop_pc_lob : _GEN_139 ? _slots_6_io_uop_pc_lob : _GEN_125 ? _slots_5_io_uop_pc_lob : _GEN_108 ? _slots_4_io_uop_pc_lob : _GEN_90 ? _slots_3_io_uop_pc_lob : _GEN_112 ? _slots_2_io_uop_pc_lob : _GEN_40 ? _slots_1_io_uop_pc_lob : _GEN_13068 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_2_taken = _GEN_595 ? _slots_39_io_uop_taken : _GEN_584 ? _slots_38_io_uop_taken : _GEN_598 ? _slots_37_io_uop_taken : _GEN_559 ? _slots_36_io_uop_taken : _GEN_545 ? _slots_35_io_uop_taken : _GEN_528 ? _slots_34_io_uop_taken : _GEN_514 ? _slots_33_io_uop_taken : _GEN_532 ? _slots_32_io_uop_taken : _GEN_489 ? _slots_31_io_uop_taken : _GEN_475 ? _slots_30_io_uop_taken : _GEN_458 ? _slots_29_io_uop_taken : _GEN_444 ? _slots_28_io_uop_taken : _GEN_462 ? _slots_27_io_uop_taken : _GEN_419 ? _slots_26_io_uop_taken : _GEN_405 ? _slots_25_io_uop_taken : _GEN_388 ? _slots_24_io_uop_taken : _GEN_374 ? _slots_23_io_uop_taken : _GEN_392 ? _slots_22_io_uop_taken : _GEN_349 ? _slots_21_io_uop_taken : _GEN_335 ? _slots_20_io_uop_taken : _GEN_318 ? _slots_19_io_uop_taken : _GEN_304 ? _slots_18_io_uop_taken : _GEN_322 ? _slots_17_io_uop_taken : _GEN_279 ? _slots_16_io_uop_taken : _GEN_265 ? _slots_15_io_uop_taken : _GEN_248 ? _slots_14_io_uop_taken : _GEN_234 ? _slots_13_io_uop_taken : _GEN_252 ? _slots_12_io_uop_taken : _GEN_209 ? _slots_11_io_uop_taken : _GEN_195 ? _slots_10_io_uop_taken : _GEN_178 ? _slots_9_io_uop_taken : _GEN_164 ? _slots_8_io_uop_taken : _GEN_182 ? _slots_7_io_uop_taken : _GEN_139 ? _slots_6_io_uop_taken : _GEN_125 ? _slots_5_io_uop_taken : _GEN_108 ? _slots_4_io_uop_taken : _GEN_90 ? _slots_3_io_uop_taken : _GEN_112 ? _slots_2_io_uop_taken : _GEN_40 ? _slots_1_io_uop_taken : _GEN_13068 & _slots_0_io_uop_taken;
  assign io_iss_uops_2_imm_packed = _GEN_595 ? _slots_39_io_uop_imm_packed : _GEN_584 ? _slots_38_io_uop_imm_packed : _GEN_598 ? _slots_37_io_uop_imm_packed : _GEN_559 ? _slots_36_io_uop_imm_packed : _GEN_545 ? _slots_35_io_uop_imm_packed : _GEN_528 ? _slots_34_io_uop_imm_packed : _GEN_514 ? _slots_33_io_uop_imm_packed : _GEN_532 ? _slots_32_io_uop_imm_packed : _GEN_489 ? _slots_31_io_uop_imm_packed : _GEN_475 ? _slots_30_io_uop_imm_packed : _GEN_458 ? _slots_29_io_uop_imm_packed : _GEN_444 ? _slots_28_io_uop_imm_packed : _GEN_462 ? _slots_27_io_uop_imm_packed : _GEN_419 ? _slots_26_io_uop_imm_packed : _GEN_405 ? _slots_25_io_uop_imm_packed : _GEN_388 ? _slots_24_io_uop_imm_packed : _GEN_374 ? _slots_23_io_uop_imm_packed : _GEN_392 ? _slots_22_io_uop_imm_packed : _GEN_349 ? _slots_21_io_uop_imm_packed : _GEN_335 ? _slots_20_io_uop_imm_packed : _GEN_318 ? _slots_19_io_uop_imm_packed : _GEN_304 ? _slots_18_io_uop_imm_packed : _GEN_322 ? _slots_17_io_uop_imm_packed : _GEN_279 ? _slots_16_io_uop_imm_packed : _GEN_265 ? _slots_15_io_uop_imm_packed : _GEN_248 ? _slots_14_io_uop_imm_packed : _GEN_234 ? _slots_13_io_uop_imm_packed : _GEN_252 ? _slots_12_io_uop_imm_packed : _GEN_209 ? _slots_11_io_uop_imm_packed : _GEN_195 ? _slots_10_io_uop_imm_packed : _GEN_178 ? _slots_9_io_uop_imm_packed : _GEN_164 ? _slots_8_io_uop_imm_packed : _GEN_182 ? _slots_7_io_uop_imm_packed : _GEN_139 ? _slots_6_io_uop_imm_packed : _GEN_125 ? _slots_5_io_uop_imm_packed : _GEN_108 ? _slots_4_io_uop_imm_packed : _GEN_90 ? _slots_3_io_uop_imm_packed : _GEN_112 ? _slots_2_io_uop_imm_packed : _GEN_40 ? _slots_1_io_uop_imm_packed : _GEN_13068 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_2_rob_idx = _GEN_595 ? _slots_39_io_uop_rob_idx : _GEN_584 ? _slots_38_io_uop_rob_idx : _GEN_598 ? _slots_37_io_uop_rob_idx : _GEN_559 ? _slots_36_io_uop_rob_idx : _GEN_545 ? _slots_35_io_uop_rob_idx : _GEN_528 ? _slots_34_io_uop_rob_idx : _GEN_514 ? _slots_33_io_uop_rob_idx : _GEN_532 ? _slots_32_io_uop_rob_idx : _GEN_489 ? _slots_31_io_uop_rob_idx : _GEN_475 ? _slots_30_io_uop_rob_idx : _GEN_458 ? _slots_29_io_uop_rob_idx : _GEN_444 ? _slots_28_io_uop_rob_idx : _GEN_462 ? _slots_27_io_uop_rob_idx : _GEN_419 ? _slots_26_io_uop_rob_idx : _GEN_405 ? _slots_25_io_uop_rob_idx : _GEN_388 ? _slots_24_io_uop_rob_idx : _GEN_374 ? _slots_23_io_uop_rob_idx : _GEN_392 ? _slots_22_io_uop_rob_idx : _GEN_349 ? _slots_21_io_uop_rob_idx : _GEN_335 ? _slots_20_io_uop_rob_idx : _GEN_318 ? _slots_19_io_uop_rob_idx : _GEN_304 ? _slots_18_io_uop_rob_idx : _GEN_322 ? _slots_17_io_uop_rob_idx : _GEN_279 ? _slots_16_io_uop_rob_idx : _GEN_265 ? _slots_15_io_uop_rob_idx : _GEN_248 ? _slots_14_io_uop_rob_idx : _GEN_234 ? _slots_13_io_uop_rob_idx : _GEN_252 ? _slots_12_io_uop_rob_idx : _GEN_209 ? _slots_11_io_uop_rob_idx : _GEN_195 ? _slots_10_io_uop_rob_idx : _GEN_178 ? _slots_9_io_uop_rob_idx : _GEN_164 ? _slots_8_io_uop_rob_idx : _GEN_182 ? _slots_7_io_uop_rob_idx : _GEN_139 ? _slots_6_io_uop_rob_idx : _GEN_125 ? _slots_5_io_uop_rob_idx : _GEN_108 ? _slots_4_io_uop_rob_idx : _GEN_90 ? _slots_3_io_uop_rob_idx : _GEN_112 ? _slots_2_io_uop_rob_idx : _GEN_40 ? _slots_1_io_uop_rob_idx : _GEN_13068 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_2_ldq_idx = _GEN_595 ? _slots_39_io_uop_ldq_idx : _GEN_584 ? _slots_38_io_uop_ldq_idx : _GEN_598 ? _slots_37_io_uop_ldq_idx : _GEN_559 ? _slots_36_io_uop_ldq_idx : _GEN_545 ? _slots_35_io_uop_ldq_idx : _GEN_528 ? _slots_34_io_uop_ldq_idx : _GEN_514 ? _slots_33_io_uop_ldq_idx : _GEN_532 ? _slots_32_io_uop_ldq_idx : _GEN_489 ? _slots_31_io_uop_ldq_idx : _GEN_475 ? _slots_30_io_uop_ldq_idx : _GEN_458 ? _slots_29_io_uop_ldq_idx : _GEN_444 ? _slots_28_io_uop_ldq_idx : _GEN_462 ? _slots_27_io_uop_ldq_idx : _GEN_419 ? _slots_26_io_uop_ldq_idx : _GEN_405 ? _slots_25_io_uop_ldq_idx : _GEN_388 ? _slots_24_io_uop_ldq_idx : _GEN_374 ? _slots_23_io_uop_ldq_idx : _GEN_392 ? _slots_22_io_uop_ldq_idx : _GEN_349 ? _slots_21_io_uop_ldq_idx : _GEN_335 ? _slots_20_io_uop_ldq_idx : _GEN_318 ? _slots_19_io_uop_ldq_idx : _GEN_304 ? _slots_18_io_uop_ldq_idx : _GEN_322 ? _slots_17_io_uop_ldq_idx : _GEN_279 ? _slots_16_io_uop_ldq_idx : _GEN_265 ? _slots_15_io_uop_ldq_idx : _GEN_248 ? _slots_14_io_uop_ldq_idx : _GEN_234 ? _slots_13_io_uop_ldq_idx : _GEN_252 ? _slots_12_io_uop_ldq_idx : _GEN_209 ? _slots_11_io_uop_ldq_idx : _GEN_195 ? _slots_10_io_uop_ldq_idx : _GEN_178 ? _slots_9_io_uop_ldq_idx : _GEN_164 ? _slots_8_io_uop_ldq_idx : _GEN_182 ? _slots_7_io_uop_ldq_idx : _GEN_139 ? _slots_6_io_uop_ldq_idx : _GEN_125 ? _slots_5_io_uop_ldq_idx : _GEN_108 ? _slots_4_io_uop_ldq_idx : _GEN_90 ? _slots_3_io_uop_ldq_idx : _GEN_112 ? _slots_2_io_uop_ldq_idx : _GEN_40 ? _slots_1_io_uop_ldq_idx : _GEN_13068 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_2_stq_idx = _GEN_595 ? _slots_39_io_uop_stq_idx : _GEN_584 ? _slots_38_io_uop_stq_idx : _GEN_598 ? _slots_37_io_uop_stq_idx : _GEN_559 ? _slots_36_io_uop_stq_idx : _GEN_545 ? _slots_35_io_uop_stq_idx : _GEN_528 ? _slots_34_io_uop_stq_idx : _GEN_514 ? _slots_33_io_uop_stq_idx : _GEN_532 ? _slots_32_io_uop_stq_idx : _GEN_489 ? _slots_31_io_uop_stq_idx : _GEN_475 ? _slots_30_io_uop_stq_idx : _GEN_458 ? _slots_29_io_uop_stq_idx : _GEN_444 ? _slots_28_io_uop_stq_idx : _GEN_462 ? _slots_27_io_uop_stq_idx : _GEN_419 ? _slots_26_io_uop_stq_idx : _GEN_405 ? _slots_25_io_uop_stq_idx : _GEN_388 ? _slots_24_io_uop_stq_idx : _GEN_374 ? _slots_23_io_uop_stq_idx : _GEN_392 ? _slots_22_io_uop_stq_idx : _GEN_349 ? _slots_21_io_uop_stq_idx : _GEN_335 ? _slots_20_io_uop_stq_idx : _GEN_318 ? _slots_19_io_uop_stq_idx : _GEN_304 ? _slots_18_io_uop_stq_idx : _GEN_322 ? _slots_17_io_uop_stq_idx : _GEN_279 ? _slots_16_io_uop_stq_idx : _GEN_265 ? _slots_15_io_uop_stq_idx : _GEN_248 ? _slots_14_io_uop_stq_idx : _GEN_234 ? _slots_13_io_uop_stq_idx : _GEN_252 ? _slots_12_io_uop_stq_idx : _GEN_209 ? _slots_11_io_uop_stq_idx : _GEN_195 ? _slots_10_io_uop_stq_idx : _GEN_178 ? _slots_9_io_uop_stq_idx : _GEN_164 ? _slots_8_io_uop_stq_idx : _GEN_182 ? _slots_7_io_uop_stq_idx : _GEN_139 ? _slots_6_io_uop_stq_idx : _GEN_125 ? _slots_5_io_uop_stq_idx : _GEN_108 ? _slots_4_io_uop_stq_idx : _GEN_90 ? _slots_3_io_uop_stq_idx : _GEN_112 ? _slots_2_io_uop_stq_idx : _GEN_40 ? _slots_1_io_uop_stq_idx : _GEN_13068 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_2_pdst = _GEN_595 ? _slots_39_io_uop_pdst : _GEN_584 ? _slots_38_io_uop_pdst : _GEN_598 ? _slots_37_io_uop_pdst : _GEN_559 ? _slots_36_io_uop_pdst : _GEN_545 ? _slots_35_io_uop_pdst : _GEN_528 ? _slots_34_io_uop_pdst : _GEN_514 ? _slots_33_io_uop_pdst : _GEN_532 ? _slots_32_io_uop_pdst : _GEN_489 ? _slots_31_io_uop_pdst : _GEN_475 ? _slots_30_io_uop_pdst : _GEN_458 ? _slots_29_io_uop_pdst : _GEN_444 ? _slots_28_io_uop_pdst : _GEN_462 ? _slots_27_io_uop_pdst : _GEN_419 ? _slots_26_io_uop_pdst : _GEN_405 ? _slots_25_io_uop_pdst : _GEN_388 ? _slots_24_io_uop_pdst : _GEN_374 ? _slots_23_io_uop_pdst : _GEN_392 ? _slots_22_io_uop_pdst : _GEN_349 ? _slots_21_io_uop_pdst : _GEN_335 ? _slots_20_io_uop_pdst : _GEN_318 ? _slots_19_io_uop_pdst : _GEN_304 ? _slots_18_io_uop_pdst : _GEN_322 ? _slots_17_io_uop_pdst : _GEN_279 ? _slots_16_io_uop_pdst : _GEN_265 ? _slots_15_io_uop_pdst : _GEN_248 ? _slots_14_io_uop_pdst : _GEN_234 ? _slots_13_io_uop_pdst : _GEN_252 ? _slots_12_io_uop_pdst : _GEN_209 ? _slots_11_io_uop_pdst : _GEN_195 ? _slots_10_io_uop_pdst : _GEN_178 ? _slots_9_io_uop_pdst : _GEN_164 ? _slots_8_io_uop_pdst : _GEN_182 ? _slots_7_io_uop_pdst : _GEN_139 ? _slots_6_io_uop_pdst : _GEN_125 ? _slots_5_io_uop_pdst : _GEN_108 ? _slots_4_io_uop_pdst : _GEN_90 ? _slots_3_io_uop_pdst : _GEN_112 ? _slots_2_io_uop_pdst : _GEN_40 ? _slots_1_io_uop_pdst : _GEN_13068 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_2_prs1 = _GEN_595 ? _slots_39_io_uop_prs1 : _GEN_584 ? _slots_38_io_uop_prs1 : _GEN_598 ? _slots_37_io_uop_prs1 : _GEN_559 ? _slots_36_io_uop_prs1 : _GEN_545 ? _slots_35_io_uop_prs1 : _GEN_528 ? _slots_34_io_uop_prs1 : _GEN_514 ? _slots_33_io_uop_prs1 : _GEN_532 ? _slots_32_io_uop_prs1 : _GEN_489 ? _slots_31_io_uop_prs1 : _GEN_475 ? _slots_30_io_uop_prs1 : _GEN_458 ? _slots_29_io_uop_prs1 : _GEN_444 ? _slots_28_io_uop_prs1 : _GEN_462 ? _slots_27_io_uop_prs1 : _GEN_419 ? _slots_26_io_uop_prs1 : _GEN_405 ? _slots_25_io_uop_prs1 : _GEN_388 ? _slots_24_io_uop_prs1 : _GEN_374 ? _slots_23_io_uop_prs1 : _GEN_392 ? _slots_22_io_uop_prs1 : _GEN_349 ? _slots_21_io_uop_prs1 : _GEN_335 ? _slots_20_io_uop_prs1 : _GEN_318 ? _slots_19_io_uop_prs1 : _GEN_304 ? _slots_18_io_uop_prs1 : _GEN_322 ? _slots_17_io_uop_prs1 : _GEN_279 ? _slots_16_io_uop_prs1 : _GEN_265 ? _slots_15_io_uop_prs1 : _GEN_248 ? _slots_14_io_uop_prs1 : _GEN_234 ? _slots_13_io_uop_prs1 : _GEN_252 ? _slots_12_io_uop_prs1 : _GEN_209 ? _slots_11_io_uop_prs1 : _GEN_195 ? _slots_10_io_uop_prs1 : _GEN_178 ? _slots_9_io_uop_prs1 : _GEN_164 ? _slots_8_io_uop_prs1 : _GEN_182 ? _slots_7_io_uop_prs1 : _GEN_139 ? _slots_6_io_uop_prs1 : _GEN_125 ? _slots_5_io_uop_prs1 : _GEN_108 ? _slots_4_io_uop_prs1 : _GEN_90 ? _slots_3_io_uop_prs1 : _GEN_112 ? _slots_2_io_uop_prs1 : _GEN_40 ? _slots_1_io_uop_prs1 : _GEN_13068 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_2_prs2 = _GEN_595 ? _slots_39_io_uop_prs2 : _GEN_584 ? _slots_38_io_uop_prs2 : _GEN_598 ? _slots_37_io_uop_prs2 : _GEN_559 ? _slots_36_io_uop_prs2 : _GEN_545 ? _slots_35_io_uop_prs2 : _GEN_528 ? _slots_34_io_uop_prs2 : _GEN_514 ? _slots_33_io_uop_prs2 : _GEN_532 ? _slots_32_io_uop_prs2 : _GEN_489 ? _slots_31_io_uop_prs2 : _GEN_475 ? _slots_30_io_uop_prs2 : _GEN_458 ? _slots_29_io_uop_prs2 : _GEN_444 ? _slots_28_io_uop_prs2 : _GEN_462 ? _slots_27_io_uop_prs2 : _GEN_419 ? _slots_26_io_uop_prs2 : _GEN_405 ? _slots_25_io_uop_prs2 : _GEN_388 ? _slots_24_io_uop_prs2 : _GEN_374 ? _slots_23_io_uop_prs2 : _GEN_392 ? _slots_22_io_uop_prs2 : _GEN_349 ? _slots_21_io_uop_prs2 : _GEN_335 ? _slots_20_io_uop_prs2 : _GEN_318 ? _slots_19_io_uop_prs2 : _GEN_304 ? _slots_18_io_uop_prs2 : _GEN_322 ? _slots_17_io_uop_prs2 : _GEN_279 ? _slots_16_io_uop_prs2 : _GEN_265 ? _slots_15_io_uop_prs2 : _GEN_248 ? _slots_14_io_uop_prs2 : _GEN_234 ? _slots_13_io_uop_prs2 : _GEN_252 ? _slots_12_io_uop_prs2 : _GEN_209 ? _slots_11_io_uop_prs2 : _GEN_195 ? _slots_10_io_uop_prs2 : _GEN_178 ? _slots_9_io_uop_prs2 : _GEN_164 ? _slots_8_io_uop_prs2 : _GEN_182 ? _slots_7_io_uop_prs2 : _GEN_139 ? _slots_6_io_uop_prs2 : _GEN_125 ? _slots_5_io_uop_prs2 : _GEN_108 ? _slots_4_io_uop_prs2 : _GEN_90 ? _slots_3_io_uop_prs2 : _GEN_112 ? _slots_2_io_uop_prs2 : _GEN_40 ? _slots_1_io_uop_prs2 : _GEN_13068 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_2_bypassable = _GEN_595 ? _slots_39_io_uop_bypassable : _GEN_584 ? _slots_38_io_uop_bypassable : _GEN_598 ? _slots_37_io_uop_bypassable : _GEN_559 ? _slots_36_io_uop_bypassable : _GEN_545 ? _slots_35_io_uop_bypassable : _GEN_528 ? _slots_34_io_uop_bypassable : _GEN_514 ? _slots_33_io_uop_bypassable : _GEN_532 ? _slots_32_io_uop_bypassable : _GEN_489 ? _slots_31_io_uop_bypassable : _GEN_475 ? _slots_30_io_uop_bypassable : _GEN_458 ? _slots_29_io_uop_bypassable : _GEN_444 ? _slots_28_io_uop_bypassable : _GEN_462 ? _slots_27_io_uop_bypassable : _GEN_419 ? _slots_26_io_uop_bypassable : _GEN_405 ? _slots_25_io_uop_bypassable : _GEN_388 ? _slots_24_io_uop_bypassable : _GEN_374 ? _slots_23_io_uop_bypassable : _GEN_392 ? _slots_22_io_uop_bypassable : _GEN_349 ? _slots_21_io_uop_bypassable : _GEN_335 ? _slots_20_io_uop_bypassable : _GEN_318 ? _slots_19_io_uop_bypassable : _GEN_304 ? _slots_18_io_uop_bypassable : _GEN_322 ? _slots_17_io_uop_bypassable : _GEN_279 ? _slots_16_io_uop_bypassable : _GEN_265 ? _slots_15_io_uop_bypassable : _GEN_248 ? _slots_14_io_uop_bypassable : _GEN_234 ? _slots_13_io_uop_bypassable : _GEN_252 ? _slots_12_io_uop_bypassable : _GEN_209 ? _slots_11_io_uop_bypassable : _GEN_195 ? _slots_10_io_uop_bypassable : _GEN_178 ? _slots_9_io_uop_bypassable : _GEN_164 ? _slots_8_io_uop_bypassable : _GEN_182 ? _slots_7_io_uop_bypassable : _GEN_139 ? _slots_6_io_uop_bypassable : _GEN_125 ? _slots_5_io_uop_bypassable : _GEN_108 ? _slots_4_io_uop_bypassable : _GEN_90 ? _slots_3_io_uop_bypassable : _GEN_112 ? _slots_2_io_uop_bypassable : _GEN_40 ? _slots_1_io_uop_bypassable : _GEN_13068 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_2_mem_cmd = _GEN_595 ? _slots_39_io_uop_mem_cmd : _GEN_584 ? _slots_38_io_uop_mem_cmd : _GEN_598 ? _slots_37_io_uop_mem_cmd : _GEN_559 ? _slots_36_io_uop_mem_cmd : _GEN_545 ? _slots_35_io_uop_mem_cmd : _GEN_528 ? _slots_34_io_uop_mem_cmd : _GEN_514 ? _slots_33_io_uop_mem_cmd : _GEN_532 ? _slots_32_io_uop_mem_cmd : _GEN_489 ? _slots_31_io_uop_mem_cmd : _GEN_475 ? _slots_30_io_uop_mem_cmd : _GEN_458 ? _slots_29_io_uop_mem_cmd : _GEN_444 ? _slots_28_io_uop_mem_cmd : _GEN_462 ? _slots_27_io_uop_mem_cmd : _GEN_419 ? _slots_26_io_uop_mem_cmd : _GEN_405 ? _slots_25_io_uop_mem_cmd : _GEN_388 ? _slots_24_io_uop_mem_cmd : _GEN_374 ? _slots_23_io_uop_mem_cmd : _GEN_392 ? _slots_22_io_uop_mem_cmd : _GEN_349 ? _slots_21_io_uop_mem_cmd : _GEN_335 ? _slots_20_io_uop_mem_cmd : _GEN_318 ? _slots_19_io_uop_mem_cmd : _GEN_304 ? _slots_18_io_uop_mem_cmd : _GEN_322 ? _slots_17_io_uop_mem_cmd : _GEN_279 ? _slots_16_io_uop_mem_cmd : _GEN_265 ? _slots_15_io_uop_mem_cmd : _GEN_248 ? _slots_14_io_uop_mem_cmd : _GEN_234 ? _slots_13_io_uop_mem_cmd : _GEN_252 ? _slots_12_io_uop_mem_cmd : _GEN_209 ? _slots_11_io_uop_mem_cmd : _GEN_195 ? _slots_10_io_uop_mem_cmd : _GEN_178 ? _slots_9_io_uop_mem_cmd : _GEN_164 ? _slots_8_io_uop_mem_cmd : _GEN_182 ? _slots_7_io_uop_mem_cmd : _GEN_139 ? _slots_6_io_uop_mem_cmd : _GEN_125 ? _slots_5_io_uop_mem_cmd : _GEN_108 ? _slots_4_io_uop_mem_cmd : _GEN_90 ? _slots_3_io_uop_mem_cmd : _GEN_112 ? _slots_2_io_uop_mem_cmd : _GEN_40 ? _slots_1_io_uop_mem_cmd : _GEN_13068 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_2_is_amo = _GEN_595 ? _slots_39_io_uop_is_amo : _GEN_584 ? _slots_38_io_uop_is_amo : _GEN_598 ? _slots_37_io_uop_is_amo : _GEN_559 ? _slots_36_io_uop_is_amo : _GEN_545 ? _slots_35_io_uop_is_amo : _GEN_528 ? _slots_34_io_uop_is_amo : _GEN_514 ? _slots_33_io_uop_is_amo : _GEN_532 ? _slots_32_io_uop_is_amo : _GEN_489 ? _slots_31_io_uop_is_amo : _GEN_475 ? _slots_30_io_uop_is_amo : _GEN_458 ? _slots_29_io_uop_is_amo : _GEN_444 ? _slots_28_io_uop_is_amo : _GEN_462 ? _slots_27_io_uop_is_amo : _GEN_419 ? _slots_26_io_uop_is_amo : _GEN_405 ? _slots_25_io_uop_is_amo : _GEN_388 ? _slots_24_io_uop_is_amo : _GEN_374 ? _slots_23_io_uop_is_amo : _GEN_392 ? _slots_22_io_uop_is_amo : _GEN_349 ? _slots_21_io_uop_is_amo : _GEN_335 ? _slots_20_io_uop_is_amo : _GEN_318 ? _slots_19_io_uop_is_amo : _GEN_304 ? _slots_18_io_uop_is_amo : _GEN_322 ? _slots_17_io_uop_is_amo : _GEN_279 ? _slots_16_io_uop_is_amo : _GEN_265 ? _slots_15_io_uop_is_amo : _GEN_248 ? _slots_14_io_uop_is_amo : _GEN_234 ? _slots_13_io_uop_is_amo : _GEN_252 ? _slots_12_io_uop_is_amo : _GEN_209 ? _slots_11_io_uop_is_amo : _GEN_195 ? _slots_10_io_uop_is_amo : _GEN_178 ? _slots_9_io_uop_is_amo : _GEN_164 ? _slots_8_io_uop_is_amo : _GEN_182 ? _slots_7_io_uop_is_amo : _GEN_139 ? _slots_6_io_uop_is_amo : _GEN_125 ? _slots_5_io_uop_is_amo : _GEN_108 ? _slots_4_io_uop_is_amo : _GEN_90 ? _slots_3_io_uop_is_amo : _GEN_112 ? _slots_2_io_uop_is_amo : _GEN_40 ? _slots_1_io_uop_is_amo : _GEN_13068 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_2_uses_stq = _GEN_595 ? _slots_39_io_uop_uses_stq : _GEN_584 ? _slots_38_io_uop_uses_stq : _GEN_598 ? _slots_37_io_uop_uses_stq : _GEN_559 ? _slots_36_io_uop_uses_stq : _GEN_545 ? _slots_35_io_uop_uses_stq : _GEN_528 ? _slots_34_io_uop_uses_stq : _GEN_514 ? _slots_33_io_uop_uses_stq : _GEN_532 ? _slots_32_io_uop_uses_stq : _GEN_489 ? _slots_31_io_uop_uses_stq : _GEN_475 ? _slots_30_io_uop_uses_stq : _GEN_458 ? _slots_29_io_uop_uses_stq : _GEN_444 ? _slots_28_io_uop_uses_stq : _GEN_462 ? _slots_27_io_uop_uses_stq : _GEN_419 ? _slots_26_io_uop_uses_stq : _GEN_405 ? _slots_25_io_uop_uses_stq : _GEN_388 ? _slots_24_io_uop_uses_stq : _GEN_374 ? _slots_23_io_uop_uses_stq : _GEN_392 ? _slots_22_io_uop_uses_stq : _GEN_349 ? _slots_21_io_uop_uses_stq : _GEN_335 ? _slots_20_io_uop_uses_stq : _GEN_318 ? _slots_19_io_uop_uses_stq : _GEN_304 ? _slots_18_io_uop_uses_stq : _GEN_322 ? _slots_17_io_uop_uses_stq : _GEN_279 ? _slots_16_io_uop_uses_stq : _GEN_265 ? _slots_15_io_uop_uses_stq : _GEN_248 ? _slots_14_io_uop_uses_stq : _GEN_234 ? _slots_13_io_uop_uses_stq : _GEN_252 ? _slots_12_io_uop_uses_stq : _GEN_209 ? _slots_11_io_uop_uses_stq : _GEN_195 ? _slots_10_io_uop_uses_stq : _GEN_178 ? _slots_9_io_uop_uses_stq : _GEN_164 ? _slots_8_io_uop_uses_stq : _GEN_182 ? _slots_7_io_uop_uses_stq : _GEN_139 ? _slots_6_io_uop_uses_stq : _GEN_125 ? _slots_5_io_uop_uses_stq : _GEN_108 ? _slots_4_io_uop_uses_stq : _GEN_90 ? _slots_3_io_uop_uses_stq : _GEN_112 ? _slots_2_io_uop_uses_stq : _GEN_40 ? _slots_1_io_uop_uses_stq : _GEN_13068 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_2_ldst_val = _GEN_595 ? _slots_39_io_uop_ldst_val : _GEN_584 ? _slots_38_io_uop_ldst_val : _GEN_598 ? _slots_37_io_uop_ldst_val : _GEN_559 ? _slots_36_io_uop_ldst_val : _GEN_545 ? _slots_35_io_uop_ldst_val : _GEN_528 ? _slots_34_io_uop_ldst_val : _GEN_514 ? _slots_33_io_uop_ldst_val : _GEN_532 ? _slots_32_io_uop_ldst_val : _GEN_489 ? _slots_31_io_uop_ldst_val : _GEN_475 ? _slots_30_io_uop_ldst_val : _GEN_458 ? _slots_29_io_uop_ldst_val : _GEN_444 ? _slots_28_io_uop_ldst_val : _GEN_462 ? _slots_27_io_uop_ldst_val : _GEN_419 ? _slots_26_io_uop_ldst_val : _GEN_405 ? _slots_25_io_uop_ldst_val : _GEN_388 ? _slots_24_io_uop_ldst_val : _GEN_374 ? _slots_23_io_uop_ldst_val : _GEN_392 ? _slots_22_io_uop_ldst_val : _GEN_349 ? _slots_21_io_uop_ldst_val : _GEN_335 ? _slots_20_io_uop_ldst_val : _GEN_318 ? _slots_19_io_uop_ldst_val : _GEN_304 ? _slots_18_io_uop_ldst_val : _GEN_322 ? _slots_17_io_uop_ldst_val : _GEN_279 ? _slots_16_io_uop_ldst_val : _GEN_265 ? _slots_15_io_uop_ldst_val : _GEN_248 ? _slots_14_io_uop_ldst_val : _GEN_234 ? _slots_13_io_uop_ldst_val : _GEN_252 ? _slots_12_io_uop_ldst_val : _GEN_209 ? _slots_11_io_uop_ldst_val : _GEN_195 ? _slots_10_io_uop_ldst_val : _GEN_178 ? _slots_9_io_uop_ldst_val : _GEN_164 ? _slots_8_io_uop_ldst_val : _GEN_182 ? _slots_7_io_uop_ldst_val : _GEN_139 ? _slots_6_io_uop_ldst_val : _GEN_125 ? _slots_5_io_uop_ldst_val : _GEN_108 ? _slots_4_io_uop_ldst_val : _GEN_90 ? _slots_3_io_uop_ldst_val : _GEN_112 ? _slots_2_io_uop_ldst_val : _GEN_40 ? _slots_1_io_uop_ldst_val : _GEN_13068 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_2_dst_rtype = _GEN_595 ? _slots_39_io_uop_dst_rtype : _GEN_584 ? _slots_38_io_uop_dst_rtype : _GEN_598 ? _slots_37_io_uop_dst_rtype : _GEN_559 ? _slots_36_io_uop_dst_rtype : _GEN_545 ? _slots_35_io_uop_dst_rtype : _GEN_528 ? _slots_34_io_uop_dst_rtype : _GEN_514 ? _slots_33_io_uop_dst_rtype : _GEN_532 ? _slots_32_io_uop_dst_rtype : _GEN_489 ? _slots_31_io_uop_dst_rtype : _GEN_475 ? _slots_30_io_uop_dst_rtype : _GEN_458 ? _slots_29_io_uop_dst_rtype : _GEN_444 ? _slots_28_io_uop_dst_rtype : _GEN_462 ? _slots_27_io_uop_dst_rtype : _GEN_419 ? _slots_26_io_uop_dst_rtype : _GEN_405 ? _slots_25_io_uop_dst_rtype : _GEN_388 ? _slots_24_io_uop_dst_rtype : _GEN_374 ? _slots_23_io_uop_dst_rtype : _GEN_392 ? _slots_22_io_uop_dst_rtype : _GEN_349 ? _slots_21_io_uop_dst_rtype : _GEN_335 ? _slots_20_io_uop_dst_rtype : _GEN_318 ? _slots_19_io_uop_dst_rtype : _GEN_304 ? _slots_18_io_uop_dst_rtype : _GEN_322 ? _slots_17_io_uop_dst_rtype : _GEN_279 ? _slots_16_io_uop_dst_rtype : _GEN_265 ? _slots_15_io_uop_dst_rtype : _GEN_248 ? _slots_14_io_uop_dst_rtype : _GEN_234 ? _slots_13_io_uop_dst_rtype : _GEN_252 ? _slots_12_io_uop_dst_rtype : _GEN_209 ? _slots_11_io_uop_dst_rtype : _GEN_195 ? _slots_10_io_uop_dst_rtype : _GEN_178 ? _slots_9_io_uop_dst_rtype : _GEN_164 ? _slots_8_io_uop_dst_rtype : _GEN_182 ? _slots_7_io_uop_dst_rtype : _GEN_139 ? _slots_6_io_uop_dst_rtype : _GEN_125 ? _slots_5_io_uop_dst_rtype : _GEN_108 ? _slots_4_io_uop_dst_rtype : _GEN_90 ? _slots_3_io_uop_dst_rtype : _GEN_112 ? _slots_2_io_uop_dst_rtype : _GEN_40 ? _slots_1_io_uop_dst_rtype : _GEN_13068 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_2_lrs1_rtype = _GEN_595 ? _slots_39_io_uop_lrs1_rtype : _GEN_584 ? _slots_38_io_uop_lrs1_rtype : _GEN_598 ? _slots_37_io_uop_lrs1_rtype : _GEN_559 ? _slots_36_io_uop_lrs1_rtype : _GEN_545 ? _slots_35_io_uop_lrs1_rtype : _GEN_528 ? _slots_34_io_uop_lrs1_rtype : _GEN_514 ? _slots_33_io_uop_lrs1_rtype : _GEN_532 ? _slots_32_io_uop_lrs1_rtype : _GEN_489 ? _slots_31_io_uop_lrs1_rtype : _GEN_475 ? _slots_30_io_uop_lrs1_rtype : _GEN_458 ? _slots_29_io_uop_lrs1_rtype : _GEN_444 ? _slots_28_io_uop_lrs1_rtype : _GEN_462 ? _slots_27_io_uop_lrs1_rtype : _GEN_419 ? _slots_26_io_uop_lrs1_rtype : _GEN_405 ? _slots_25_io_uop_lrs1_rtype : _GEN_388 ? _slots_24_io_uop_lrs1_rtype : _GEN_374 ? _slots_23_io_uop_lrs1_rtype : _GEN_392 ? _slots_22_io_uop_lrs1_rtype : _GEN_349 ? _slots_21_io_uop_lrs1_rtype : _GEN_335 ? _slots_20_io_uop_lrs1_rtype : _GEN_318 ? _slots_19_io_uop_lrs1_rtype : _GEN_304 ? _slots_18_io_uop_lrs1_rtype : _GEN_322 ? _slots_17_io_uop_lrs1_rtype : _GEN_279 ? _slots_16_io_uop_lrs1_rtype : _GEN_265 ? _slots_15_io_uop_lrs1_rtype : _GEN_248 ? _slots_14_io_uop_lrs1_rtype : _GEN_234 ? _slots_13_io_uop_lrs1_rtype : _GEN_252 ? _slots_12_io_uop_lrs1_rtype : _GEN_209 ? _slots_11_io_uop_lrs1_rtype : _GEN_195 ? _slots_10_io_uop_lrs1_rtype : _GEN_178 ? _slots_9_io_uop_lrs1_rtype : _GEN_164 ? _slots_8_io_uop_lrs1_rtype : _GEN_182 ? _slots_7_io_uop_lrs1_rtype : _GEN_139 ? _slots_6_io_uop_lrs1_rtype : _GEN_125 ? _slots_5_io_uop_lrs1_rtype : _GEN_108 ? _slots_4_io_uop_lrs1_rtype : _GEN_90 ? _slots_3_io_uop_lrs1_rtype : _GEN_112 ? _slots_2_io_uop_lrs1_rtype : _GEN_40 ? _slots_1_io_uop_lrs1_rtype : _GEN_13068 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_2_lrs2_rtype = _GEN_595 ? _slots_39_io_uop_lrs2_rtype : _GEN_584 ? _slots_38_io_uop_lrs2_rtype : _GEN_598 ? _slots_37_io_uop_lrs2_rtype : _GEN_559 ? _slots_36_io_uop_lrs2_rtype : _GEN_545 ? _slots_35_io_uop_lrs2_rtype : _GEN_528 ? _slots_34_io_uop_lrs2_rtype : _GEN_514 ? _slots_33_io_uop_lrs2_rtype : _GEN_532 ? _slots_32_io_uop_lrs2_rtype : _GEN_489 ? _slots_31_io_uop_lrs2_rtype : _GEN_475 ? _slots_30_io_uop_lrs2_rtype : _GEN_458 ? _slots_29_io_uop_lrs2_rtype : _GEN_444 ? _slots_28_io_uop_lrs2_rtype : _GEN_462 ? _slots_27_io_uop_lrs2_rtype : _GEN_419 ? _slots_26_io_uop_lrs2_rtype : _GEN_405 ? _slots_25_io_uop_lrs2_rtype : _GEN_388 ? _slots_24_io_uop_lrs2_rtype : _GEN_374 ? _slots_23_io_uop_lrs2_rtype : _GEN_392 ? _slots_22_io_uop_lrs2_rtype : _GEN_349 ? _slots_21_io_uop_lrs2_rtype : _GEN_335 ? _slots_20_io_uop_lrs2_rtype : _GEN_318 ? _slots_19_io_uop_lrs2_rtype : _GEN_304 ? _slots_18_io_uop_lrs2_rtype : _GEN_322 ? _slots_17_io_uop_lrs2_rtype : _GEN_279 ? _slots_16_io_uop_lrs2_rtype : _GEN_265 ? _slots_15_io_uop_lrs2_rtype : _GEN_248 ? _slots_14_io_uop_lrs2_rtype : _GEN_234 ? _slots_13_io_uop_lrs2_rtype : _GEN_252 ? _slots_12_io_uop_lrs2_rtype : _GEN_209 ? _slots_11_io_uop_lrs2_rtype : _GEN_195 ? _slots_10_io_uop_lrs2_rtype : _GEN_178 ? _slots_9_io_uop_lrs2_rtype : _GEN_164 ? _slots_8_io_uop_lrs2_rtype : _GEN_182 ? _slots_7_io_uop_lrs2_rtype : _GEN_139 ? _slots_6_io_uop_lrs2_rtype : _GEN_125 ? _slots_5_io_uop_lrs2_rtype : _GEN_108 ? _slots_4_io_uop_lrs2_rtype : _GEN_90 ? _slots_3_io_uop_lrs2_rtype : _GEN_112 ? _slots_2_io_uop_lrs2_rtype : _GEN_40 ? _slots_1_io_uop_lrs2_rtype : _GEN_13068 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
  assign io_iss_uops_3_uopc = _GEN_594 ? _slots_39_io_uop_uopc : _GEN_582 ? _slots_38_io_uop_uopc : _GEN_597 ? _slots_37_io_uop_uopc : _GEN_557 ? _slots_36_io_uop_uopc : _GEN_543 ? _slots_35_io_uop_uopc : _GEN_526 ? _slots_34_io_uop_uopc : _GEN_512 ? _slots_33_io_uop_uopc : _GEN_531 ? _slots_32_io_uop_uopc : _GEN_487 ? _slots_31_io_uop_uopc : _GEN_473 ? _slots_30_io_uop_uopc : _GEN_456 ? _slots_29_io_uop_uopc : _GEN_442 ? _slots_28_io_uop_uopc : _GEN_461 ? _slots_27_io_uop_uopc : _GEN_417 ? _slots_26_io_uop_uopc : _GEN_403 ? _slots_25_io_uop_uopc : _GEN_386 ? _slots_24_io_uop_uopc : _GEN_372 ? _slots_23_io_uop_uopc : _GEN_391 ? _slots_22_io_uop_uopc : _GEN_347 ? _slots_21_io_uop_uopc : _GEN_333 ? _slots_20_io_uop_uopc : _GEN_316 ? _slots_19_io_uop_uopc : _GEN_302 ? _slots_18_io_uop_uopc : _GEN_321 ? _slots_17_io_uop_uopc : _GEN_277 ? _slots_16_io_uop_uopc : _GEN_263 ? _slots_15_io_uop_uopc : _GEN_246 ? _slots_14_io_uop_uopc : _GEN_232 ? _slots_13_io_uop_uopc : _GEN_251 ? _slots_12_io_uop_uopc : _GEN_207 ? _slots_11_io_uop_uopc : _GEN_193 ? _slots_10_io_uop_uopc : _GEN_176 ? _slots_9_io_uop_uopc : _GEN_162 ? _slots_8_io_uop_uopc : _GEN_181 ? _slots_7_io_uop_uopc : _GEN_137 ? _slots_6_io_uop_uopc : _GEN_123 ? _slots_5_io_uop_uopc : _GEN_106 ? _slots_4_io_uop_uopc : _GEN_86 ? _slots_3_io_uop_uopc : _GEN_111 ? _slots_2_io_uop_uopc : _GEN_36 ? _slots_1_io_uop_uopc : _GEN_13149 ? _slots_0_io_uop_uopc : 7'h0;
  assign io_iss_uops_3_is_rvc = _GEN_594 ? _slots_39_io_uop_is_rvc : _GEN_582 ? _slots_38_io_uop_is_rvc : _GEN_597 ? _slots_37_io_uop_is_rvc : _GEN_557 ? _slots_36_io_uop_is_rvc : _GEN_543 ? _slots_35_io_uop_is_rvc : _GEN_526 ? _slots_34_io_uop_is_rvc : _GEN_512 ? _slots_33_io_uop_is_rvc : _GEN_531 ? _slots_32_io_uop_is_rvc : _GEN_487 ? _slots_31_io_uop_is_rvc : _GEN_473 ? _slots_30_io_uop_is_rvc : _GEN_456 ? _slots_29_io_uop_is_rvc : _GEN_442 ? _slots_28_io_uop_is_rvc : _GEN_461 ? _slots_27_io_uop_is_rvc : _GEN_417 ? _slots_26_io_uop_is_rvc : _GEN_403 ? _slots_25_io_uop_is_rvc : _GEN_386 ? _slots_24_io_uop_is_rvc : _GEN_372 ? _slots_23_io_uop_is_rvc : _GEN_391 ? _slots_22_io_uop_is_rvc : _GEN_347 ? _slots_21_io_uop_is_rvc : _GEN_333 ? _slots_20_io_uop_is_rvc : _GEN_316 ? _slots_19_io_uop_is_rvc : _GEN_302 ? _slots_18_io_uop_is_rvc : _GEN_321 ? _slots_17_io_uop_is_rvc : _GEN_277 ? _slots_16_io_uop_is_rvc : _GEN_263 ? _slots_15_io_uop_is_rvc : _GEN_246 ? _slots_14_io_uop_is_rvc : _GEN_232 ? _slots_13_io_uop_is_rvc : _GEN_251 ? _slots_12_io_uop_is_rvc : _GEN_207 ? _slots_11_io_uop_is_rvc : _GEN_193 ? _slots_10_io_uop_is_rvc : _GEN_176 ? _slots_9_io_uop_is_rvc : _GEN_162 ? _slots_8_io_uop_is_rvc : _GEN_181 ? _slots_7_io_uop_is_rvc : _GEN_137 ? _slots_6_io_uop_is_rvc : _GEN_123 ? _slots_5_io_uop_is_rvc : _GEN_106 ? _slots_4_io_uop_is_rvc : _GEN_86 ? _slots_3_io_uop_is_rvc : _GEN_111 ? _slots_2_io_uop_is_rvc : _GEN_36 ? _slots_1_io_uop_is_rvc : _GEN_13149 & _slots_0_io_uop_is_rvc;
  assign io_iss_uops_3_fu_code = _GEN_594 ? _slots_39_io_uop_fu_code : _GEN_582 ? _slots_38_io_uop_fu_code : _GEN_597 ? _slots_37_io_uop_fu_code : _GEN_557 ? _slots_36_io_uop_fu_code : _GEN_543 ? _slots_35_io_uop_fu_code : _GEN_526 ? _slots_34_io_uop_fu_code : _GEN_512 ? _slots_33_io_uop_fu_code : _GEN_531 ? _slots_32_io_uop_fu_code : _GEN_487 ? _slots_31_io_uop_fu_code : _GEN_473 ? _slots_30_io_uop_fu_code : _GEN_456 ? _slots_29_io_uop_fu_code : _GEN_442 ? _slots_28_io_uop_fu_code : _GEN_461 ? _slots_27_io_uop_fu_code : _GEN_417 ? _slots_26_io_uop_fu_code : _GEN_403 ? _slots_25_io_uop_fu_code : _GEN_386 ? _slots_24_io_uop_fu_code : _GEN_372 ? _slots_23_io_uop_fu_code : _GEN_391 ? _slots_22_io_uop_fu_code : _GEN_347 ? _slots_21_io_uop_fu_code : _GEN_333 ? _slots_20_io_uop_fu_code : _GEN_316 ? _slots_19_io_uop_fu_code : _GEN_302 ? _slots_18_io_uop_fu_code : _GEN_321 ? _slots_17_io_uop_fu_code : _GEN_277 ? _slots_16_io_uop_fu_code : _GEN_263 ? _slots_15_io_uop_fu_code : _GEN_246 ? _slots_14_io_uop_fu_code : _GEN_232 ? _slots_13_io_uop_fu_code : _GEN_251 ? _slots_12_io_uop_fu_code : _GEN_207 ? _slots_11_io_uop_fu_code : _GEN_193 ? _slots_10_io_uop_fu_code : _GEN_176 ? _slots_9_io_uop_fu_code : _GEN_162 ? _slots_8_io_uop_fu_code : _GEN_181 ? _slots_7_io_uop_fu_code : _GEN_137 ? _slots_6_io_uop_fu_code : _GEN_123 ? _slots_5_io_uop_fu_code : _GEN_106 ? _slots_4_io_uop_fu_code : _GEN_86 ? _slots_3_io_uop_fu_code : _GEN_111 ? _slots_2_io_uop_fu_code : _GEN_36 ? _slots_1_io_uop_fu_code : _GEN_13149 ? _slots_0_io_uop_fu_code : 10'h0;
  assign io_iss_uops_3_iw_p1_poisoned = _GEN_594 ? _slots_39_io_uop_iw_p1_poisoned : _GEN_582 ? _slots_38_io_uop_iw_p1_poisoned : _GEN_597 ? _slots_37_io_uop_iw_p1_poisoned : _GEN_557 ? _slots_36_io_uop_iw_p1_poisoned : _GEN_543 ? _slots_35_io_uop_iw_p1_poisoned : _GEN_526 ? _slots_34_io_uop_iw_p1_poisoned : _GEN_512 ? _slots_33_io_uop_iw_p1_poisoned : _GEN_531 ? _slots_32_io_uop_iw_p1_poisoned : _GEN_487 ? _slots_31_io_uop_iw_p1_poisoned : _GEN_473 ? _slots_30_io_uop_iw_p1_poisoned : _GEN_456 ? _slots_29_io_uop_iw_p1_poisoned : _GEN_442 ? _slots_28_io_uop_iw_p1_poisoned : _GEN_461 ? _slots_27_io_uop_iw_p1_poisoned : _GEN_417 ? _slots_26_io_uop_iw_p1_poisoned : _GEN_403 ? _slots_25_io_uop_iw_p1_poisoned : _GEN_386 ? _slots_24_io_uop_iw_p1_poisoned : _GEN_372 ? _slots_23_io_uop_iw_p1_poisoned : _GEN_391 ? _slots_22_io_uop_iw_p1_poisoned : _GEN_347 ? _slots_21_io_uop_iw_p1_poisoned : _GEN_333 ? _slots_20_io_uop_iw_p1_poisoned : _GEN_316 ? _slots_19_io_uop_iw_p1_poisoned : _GEN_302 ? _slots_18_io_uop_iw_p1_poisoned : _GEN_321 ? _slots_17_io_uop_iw_p1_poisoned : _GEN_277 ? _slots_16_io_uop_iw_p1_poisoned : _GEN_263 ? _slots_15_io_uop_iw_p1_poisoned : _GEN_246 ? _slots_14_io_uop_iw_p1_poisoned : _GEN_232 ? _slots_13_io_uop_iw_p1_poisoned : _GEN_251 ? _slots_12_io_uop_iw_p1_poisoned : _GEN_207 ? _slots_11_io_uop_iw_p1_poisoned : _GEN_193 ? _slots_10_io_uop_iw_p1_poisoned : _GEN_176 ? _slots_9_io_uop_iw_p1_poisoned : _GEN_162 ? _slots_8_io_uop_iw_p1_poisoned : _GEN_181 ? _slots_7_io_uop_iw_p1_poisoned : _GEN_137 ? _slots_6_io_uop_iw_p1_poisoned : _GEN_123 ? _slots_5_io_uop_iw_p1_poisoned : _GEN_106 ? _slots_4_io_uop_iw_p1_poisoned : _GEN_86 ? _slots_3_io_uop_iw_p1_poisoned : _GEN_111 ? _slots_2_io_uop_iw_p1_poisoned : _GEN_36 ? _slots_1_io_uop_iw_p1_poisoned : _GEN_13149 & _slots_0_io_uop_iw_p1_poisoned;
  assign io_iss_uops_3_iw_p2_poisoned = _GEN_594 ? _slots_39_io_uop_iw_p2_poisoned : _GEN_582 ? _slots_38_io_uop_iw_p2_poisoned : _GEN_597 ? _slots_37_io_uop_iw_p2_poisoned : _GEN_557 ? _slots_36_io_uop_iw_p2_poisoned : _GEN_543 ? _slots_35_io_uop_iw_p2_poisoned : _GEN_526 ? _slots_34_io_uop_iw_p2_poisoned : _GEN_512 ? _slots_33_io_uop_iw_p2_poisoned : _GEN_531 ? _slots_32_io_uop_iw_p2_poisoned : _GEN_487 ? _slots_31_io_uop_iw_p2_poisoned : _GEN_473 ? _slots_30_io_uop_iw_p2_poisoned : _GEN_456 ? _slots_29_io_uop_iw_p2_poisoned : _GEN_442 ? _slots_28_io_uop_iw_p2_poisoned : _GEN_461 ? _slots_27_io_uop_iw_p2_poisoned : _GEN_417 ? _slots_26_io_uop_iw_p2_poisoned : _GEN_403 ? _slots_25_io_uop_iw_p2_poisoned : _GEN_386 ? _slots_24_io_uop_iw_p2_poisoned : _GEN_372 ? _slots_23_io_uop_iw_p2_poisoned : _GEN_391 ? _slots_22_io_uop_iw_p2_poisoned : _GEN_347 ? _slots_21_io_uop_iw_p2_poisoned : _GEN_333 ? _slots_20_io_uop_iw_p2_poisoned : _GEN_316 ? _slots_19_io_uop_iw_p2_poisoned : _GEN_302 ? _slots_18_io_uop_iw_p2_poisoned : _GEN_321 ? _slots_17_io_uop_iw_p2_poisoned : _GEN_277 ? _slots_16_io_uop_iw_p2_poisoned : _GEN_263 ? _slots_15_io_uop_iw_p2_poisoned : _GEN_246 ? _slots_14_io_uop_iw_p2_poisoned : _GEN_232 ? _slots_13_io_uop_iw_p2_poisoned : _GEN_251 ? _slots_12_io_uop_iw_p2_poisoned : _GEN_207 ? _slots_11_io_uop_iw_p2_poisoned : _GEN_193 ? _slots_10_io_uop_iw_p2_poisoned : _GEN_176 ? _slots_9_io_uop_iw_p2_poisoned : _GEN_162 ? _slots_8_io_uop_iw_p2_poisoned : _GEN_181 ? _slots_7_io_uop_iw_p2_poisoned : _GEN_137 ? _slots_6_io_uop_iw_p2_poisoned : _GEN_123 ? _slots_5_io_uop_iw_p2_poisoned : _GEN_106 ? _slots_4_io_uop_iw_p2_poisoned : _GEN_86 ? _slots_3_io_uop_iw_p2_poisoned : _GEN_111 ? _slots_2_io_uop_iw_p2_poisoned : _GEN_36 ? _slots_1_io_uop_iw_p2_poisoned : _GEN_13149 & _slots_0_io_uop_iw_p2_poisoned;
  assign io_iss_uops_3_is_br = _GEN_594 ? _slots_39_io_uop_is_br : _GEN_582 ? _slots_38_io_uop_is_br : _GEN_597 ? _slots_37_io_uop_is_br : _GEN_557 ? _slots_36_io_uop_is_br : _GEN_543 ? _slots_35_io_uop_is_br : _GEN_526 ? _slots_34_io_uop_is_br : _GEN_512 ? _slots_33_io_uop_is_br : _GEN_531 ? _slots_32_io_uop_is_br : _GEN_487 ? _slots_31_io_uop_is_br : _GEN_473 ? _slots_30_io_uop_is_br : _GEN_456 ? _slots_29_io_uop_is_br : _GEN_442 ? _slots_28_io_uop_is_br : _GEN_461 ? _slots_27_io_uop_is_br : _GEN_417 ? _slots_26_io_uop_is_br : _GEN_403 ? _slots_25_io_uop_is_br : _GEN_386 ? _slots_24_io_uop_is_br : _GEN_372 ? _slots_23_io_uop_is_br : _GEN_391 ? _slots_22_io_uop_is_br : _GEN_347 ? _slots_21_io_uop_is_br : _GEN_333 ? _slots_20_io_uop_is_br : _GEN_316 ? _slots_19_io_uop_is_br : _GEN_302 ? _slots_18_io_uop_is_br : _GEN_321 ? _slots_17_io_uop_is_br : _GEN_277 ? _slots_16_io_uop_is_br : _GEN_263 ? _slots_15_io_uop_is_br : _GEN_246 ? _slots_14_io_uop_is_br : _GEN_232 ? _slots_13_io_uop_is_br : _GEN_251 ? _slots_12_io_uop_is_br : _GEN_207 ? _slots_11_io_uop_is_br : _GEN_193 ? _slots_10_io_uop_is_br : _GEN_176 ? _slots_9_io_uop_is_br : _GEN_162 ? _slots_8_io_uop_is_br : _GEN_181 ? _slots_7_io_uop_is_br : _GEN_137 ? _slots_6_io_uop_is_br : _GEN_123 ? _slots_5_io_uop_is_br : _GEN_106 ? _slots_4_io_uop_is_br : _GEN_86 ? _slots_3_io_uop_is_br : _GEN_111 ? _slots_2_io_uop_is_br : _GEN_36 ? _slots_1_io_uop_is_br : _GEN_13149 & _slots_0_io_uop_is_br;
  assign io_iss_uops_3_is_jalr = _GEN_594 ? _slots_39_io_uop_is_jalr : _GEN_582 ? _slots_38_io_uop_is_jalr : _GEN_597 ? _slots_37_io_uop_is_jalr : _GEN_557 ? _slots_36_io_uop_is_jalr : _GEN_543 ? _slots_35_io_uop_is_jalr : _GEN_526 ? _slots_34_io_uop_is_jalr : _GEN_512 ? _slots_33_io_uop_is_jalr : _GEN_531 ? _slots_32_io_uop_is_jalr : _GEN_487 ? _slots_31_io_uop_is_jalr : _GEN_473 ? _slots_30_io_uop_is_jalr : _GEN_456 ? _slots_29_io_uop_is_jalr : _GEN_442 ? _slots_28_io_uop_is_jalr : _GEN_461 ? _slots_27_io_uop_is_jalr : _GEN_417 ? _slots_26_io_uop_is_jalr : _GEN_403 ? _slots_25_io_uop_is_jalr : _GEN_386 ? _slots_24_io_uop_is_jalr : _GEN_372 ? _slots_23_io_uop_is_jalr : _GEN_391 ? _slots_22_io_uop_is_jalr : _GEN_347 ? _slots_21_io_uop_is_jalr : _GEN_333 ? _slots_20_io_uop_is_jalr : _GEN_316 ? _slots_19_io_uop_is_jalr : _GEN_302 ? _slots_18_io_uop_is_jalr : _GEN_321 ? _slots_17_io_uop_is_jalr : _GEN_277 ? _slots_16_io_uop_is_jalr : _GEN_263 ? _slots_15_io_uop_is_jalr : _GEN_246 ? _slots_14_io_uop_is_jalr : _GEN_232 ? _slots_13_io_uop_is_jalr : _GEN_251 ? _slots_12_io_uop_is_jalr : _GEN_207 ? _slots_11_io_uop_is_jalr : _GEN_193 ? _slots_10_io_uop_is_jalr : _GEN_176 ? _slots_9_io_uop_is_jalr : _GEN_162 ? _slots_8_io_uop_is_jalr : _GEN_181 ? _slots_7_io_uop_is_jalr : _GEN_137 ? _slots_6_io_uop_is_jalr : _GEN_123 ? _slots_5_io_uop_is_jalr : _GEN_106 ? _slots_4_io_uop_is_jalr : _GEN_86 ? _slots_3_io_uop_is_jalr : _GEN_111 ? _slots_2_io_uop_is_jalr : _GEN_36 ? _slots_1_io_uop_is_jalr : _GEN_13149 & _slots_0_io_uop_is_jalr;
  assign io_iss_uops_3_is_jal = _GEN_594 ? _slots_39_io_uop_is_jal : _GEN_582 ? _slots_38_io_uop_is_jal : _GEN_597 ? _slots_37_io_uop_is_jal : _GEN_557 ? _slots_36_io_uop_is_jal : _GEN_543 ? _slots_35_io_uop_is_jal : _GEN_526 ? _slots_34_io_uop_is_jal : _GEN_512 ? _slots_33_io_uop_is_jal : _GEN_531 ? _slots_32_io_uop_is_jal : _GEN_487 ? _slots_31_io_uop_is_jal : _GEN_473 ? _slots_30_io_uop_is_jal : _GEN_456 ? _slots_29_io_uop_is_jal : _GEN_442 ? _slots_28_io_uop_is_jal : _GEN_461 ? _slots_27_io_uop_is_jal : _GEN_417 ? _slots_26_io_uop_is_jal : _GEN_403 ? _slots_25_io_uop_is_jal : _GEN_386 ? _slots_24_io_uop_is_jal : _GEN_372 ? _slots_23_io_uop_is_jal : _GEN_391 ? _slots_22_io_uop_is_jal : _GEN_347 ? _slots_21_io_uop_is_jal : _GEN_333 ? _slots_20_io_uop_is_jal : _GEN_316 ? _slots_19_io_uop_is_jal : _GEN_302 ? _slots_18_io_uop_is_jal : _GEN_321 ? _slots_17_io_uop_is_jal : _GEN_277 ? _slots_16_io_uop_is_jal : _GEN_263 ? _slots_15_io_uop_is_jal : _GEN_246 ? _slots_14_io_uop_is_jal : _GEN_232 ? _slots_13_io_uop_is_jal : _GEN_251 ? _slots_12_io_uop_is_jal : _GEN_207 ? _slots_11_io_uop_is_jal : _GEN_193 ? _slots_10_io_uop_is_jal : _GEN_176 ? _slots_9_io_uop_is_jal : _GEN_162 ? _slots_8_io_uop_is_jal : _GEN_181 ? _slots_7_io_uop_is_jal : _GEN_137 ? _slots_6_io_uop_is_jal : _GEN_123 ? _slots_5_io_uop_is_jal : _GEN_106 ? _slots_4_io_uop_is_jal : _GEN_86 ? _slots_3_io_uop_is_jal : _GEN_111 ? _slots_2_io_uop_is_jal : _GEN_36 ? _slots_1_io_uop_is_jal : _GEN_13149 & _slots_0_io_uop_is_jal;
  assign io_iss_uops_3_is_sfb = _GEN_594 ? _slots_39_io_uop_is_sfb : _GEN_582 ? _slots_38_io_uop_is_sfb : _GEN_597 ? _slots_37_io_uop_is_sfb : _GEN_557 ? _slots_36_io_uop_is_sfb : _GEN_543 ? _slots_35_io_uop_is_sfb : _GEN_526 ? _slots_34_io_uop_is_sfb : _GEN_512 ? _slots_33_io_uop_is_sfb : _GEN_531 ? _slots_32_io_uop_is_sfb : _GEN_487 ? _slots_31_io_uop_is_sfb : _GEN_473 ? _slots_30_io_uop_is_sfb : _GEN_456 ? _slots_29_io_uop_is_sfb : _GEN_442 ? _slots_28_io_uop_is_sfb : _GEN_461 ? _slots_27_io_uop_is_sfb : _GEN_417 ? _slots_26_io_uop_is_sfb : _GEN_403 ? _slots_25_io_uop_is_sfb : _GEN_386 ? _slots_24_io_uop_is_sfb : _GEN_372 ? _slots_23_io_uop_is_sfb : _GEN_391 ? _slots_22_io_uop_is_sfb : _GEN_347 ? _slots_21_io_uop_is_sfb : _GEN_333 ? _slots_20_io_uop_is_sfb : _GEN_316 ? _slots_19_io_uop_is_sfb : _GEN_302 ? _slots_18_io_uop_is_sfb : _GEN_321 ? _slots_17_io_uop_is_sfb : _GEN_277 ? _slots_16_io_uop_is_sfb : _GEN_263 ? _slots_15_io_uop_is_sfb : _GEN_246 ? _slots_14_io_uop_is_sfb : _GEN_232 ? _slots_13_io_uop_is_sfb : _GEN_251 ? _slots_12_io_uop_is_sfb : _GEN_207 ? _slots_11_io_uop_is_sfb : _GEN_193 ? _slots_10_io_uop_is_sfb : _GEN_176 ? _slots_9_io_uop_is_sfb : _GEN_162 ? _slots_8_io_uop_is_sfb : _GEN_181 ? _slots_7_io_uop_is_sfb : _GEN_137 ? _slots_6_io_uop_is_sfb : _GEN_123 ? _slots_5_io_uop_is_sfb : _GEN_106 ? _slots_4_io_uop_is_sfb : _GEN_86 ? _slots_3_io_uop_is_sfb : _GEN_111 ? _slots_2_io_uop_is_sfb : _GEN_36 ? _slots_1_io_uop_is_sfb : _GEN_13149 & _slots_0_io_uop_is_sfb;
  assign io_iss_uops_3_br_mask = _GEN_594 ? _slots_39_io_uop_br_mask : _GEN_582 ? _slots_38_io_uop_br_mask : _GEN_597 ? _slots_37_io_uop_br_mask : _GEN_557 ? _slots_36_io_uop_br_mask : _GEN_543 ? _slots_35_io_uop_br_mask : _GEN_526 ? _slots_34_io_uop_br_mask : _GEN_512 ? _slots_33_io_uop_br_mask : _GEN_531 ? _slots_32_io_uop_br_mask : _GEN_487 ? _slots_31_io_uop_br_mask : _GEN_473 ? _slots_30_io_uop_br_mask : _GEN_456 ? _slots_29_io_uop_br_mask : _GEN_442 ? _slots_28_io_uop_br_mask : _GEN_461 ? _slots_27_io_uop_br_mask : _GEN_417 ? _slots_26_io_uop_br_mask : _GEN_403 ? _slots_25_io_uop_br_mask : _GEN_386 ? _slots_24_io_uop_br_mask : _GEN_372 ? _slots_23_io_uop_br_mask : _GEN_391 ? _slots_22_io_uop_br_mask : _GEN_347 ? _slots_21_io_uop_br_mask : _GEN_333 ? _slots_20_io_uop_br_mask : _GEN_316 ? _slots_19_io_uop_br_mask : _GEN_302 ? _slots_18_io_uop_br_mask : _GEN_321 ? _slots_17_io_uop_br_mask : _GEN_277 ? _slots_16_io_uop_br_mask : _GEN_263 ? _slots_15_io_uop_br_mask : _GEN_246 ? _slots_14_io_uop_br_mask : _GEN_232 ? _slots_13_io_uop_br_mask : _GEN_251 ? _slots_12_io_uop_br_mask : _GEN_207 ? _slots_11_io_uop_br_mask : _GEN_193 ? _slots_10_io_uop_br_mask : _GEN_176 ? _slots_9_io_uop_br_mask : _GEN_162 ? _slots_8_io_uop_br_mask : _GEN_181 ? _slots_7_io_uop_br_mask : _GEN_137 ? _slots_6_io_uop_br_mask : _GEN_123 ? _slots_5_io_uop_br_mask : _GEN_106 ? _slots_4_io_uop_br_mask : _GEN_86 ? _slots_3_io_uop_br_mask : _GEN_111 ? _slots_2_io_uop_br_mask : _GEN_36 ? _slots_1_io_uop_br_mask : _GEN_13149 ? _slots_0_io_uop_br_mask : 20'h0;
  assign io_iss_uops_3_br_tag = _GEN_594 ? _slots_39_io_uop_br_tag : _GEN_582 ? _slots_38_io_uop_br_tag : _GEN_597 ? _slots_37_io_uop_br_tag : _GEN_557 ? _slots_36_io_uop_br_tag : _GEN_543 ? _slots_35_io_uop_br_tag : _GEN_526 ? _slots_34_io_uop_br_tag : _GEN_512 ? _slots_33_io_uop_br_tag : _GEN_531 ? _slots_32_io_uop_br_tag : _GEN_487 ? _slots_31_io_uop_br_tag : _GEN_473 ? _slots_30_io_uop_br_tag : _GEN_456 ? _slots_29_io_uop_br_tag : _GEN_442 ? _slots_28_io_uop_br_tag : _GEN_461 ? _slots_27_io_uop_br_tag : _GEN_417 ? _slots_26_io_uop_br_tag : _GEN_403 ? _slots_25_io_uop_br_tag : _GEN_386 ? _slots_24_io_uop_br_tag : _GEN_372 ? _slots_23_io_uop_br_tag : _GEN_391 ? _slots_22_io_uop_br_tag : _GEN_347 ? _slots_21_io_uop_br_tag : _GEN_333 ? _slots_20_io_uop_br_tag : _GEN_316 ? _slots_19_io_uop_br_tag : _GEN_302 ? _slots_18_io_uop_br_tag : _GEN_321 ? _slots_17_io_uop_br_tag : _GEN_277 ? _slots_16_io_uop_br_tag : _GEN_263 ? _slots_15_io_uop_br_tag : _GEN_246 ? _slots_14_io_uop_br_tag : _GEN_232 ? _slots_13_io_uop_br_tag : _GEN_251 ? _slots_12_io_uop_br_tag : _GEN_207 ? _slots_11_io_uop_br_tag : _GEN_193 ? _slots_10_io_uop_br_tag : _GEN_176 ? _slots_9_io_uop_br_tag : _GEN_162 ? _slots_8_io_uop_br_tag : _GEN_181 ? _slots_7_io_uop_br_tag : _GEN_137 ? _slots_6_io_uop_br_tag : _GEN_123 ? _slots_5_io_uop_br_tag : _GEN_106 ? _slots_4_io_uop_br_tag : _GEN_86 ? _slots_3_io_uop_br_tag : _GEN_111 ? _slots_2_io_uop_br_tag : _GEN_36 ? _slots_1_io_uop_br_tag : _GEN_13149 ? _slots_0_io_uop_br_tag : 5'h0;
  assign io_iss_uops_3_ftq_idx = _GEN_594 ? _slots_39_io_uop_ftq_idx : _GEN_582 ? _slots_38_io_uop_ftq_idx : _GEN_597 ? _slots_37_io_uop_ftq_idx : _GEN_557 ? _slots_36_io_uop_ftq_idx : _GEN_543 ? _slots_35_io_uop_ftq_idx : _GEN_526 ? _slots_34_io_uop_ftq_idx : _GEN_512 ? _slots_33_io_uop_ftq_idx : _GEN_531 ? _slots_32_io_uop_ftq_idx : _GEN_487 ? _slots_31_io_uop_ftq_idx : _GEN_473 ? _slots_30_io_uop_ftq_idx : _GEN_456 ? _slots_29_io_uop_ftq_idx : _GEN_442 ? _slots_28_io_uop_ftq_idx : _GEN_461 ? _slots_27_io_uop_ftq_idx : _GEN_417 ? _slots_26_io_uop_ftq_idx : _GEN_403 ? _slots_25_io_uop_ftq_idx : _GEN_386 ? _slots_24_io_uop_ftq_idx : _GEN_372 ? _slots_23_io_uop_ftq_idx : _GEN_391 ? _slots_22_io_uop_ftq_idx : _GEN_347 ? _slots_21_io_uop_ftq_idx : _GEN_333 ? _slots_20_io_uop_ftq_idx : _GEN_316 ? _slots_19_io_uop_ftq_idx : _GEN_302 ? _slots_18_io_uop_ftq_idx : _GEN_321 ? _slots_17_io_uop_ftq_idx : _GEN_277 ? _slots_16_io_uop_ftq_idx : _GEN_263 ? _slots_15_io_uop_ftq_idx : _GEN_246 ? _slots_14_io_uop_ftq_idx : _GEN_232 ? _slots_13_io_uop_ftq_idx : _GEN_251 ? _slots_12_io_uop_ftq_idx : _GEN_207 ? _slots_11_io_uop_ftq_idx : _GEN_193 ? _slots_10_io_uop_ftq_idx : _GEN_176 ? _slots_9_io_uop_ftq_idx : _GEN_162 ? _slots_8_io_uop_ftq_idx : _GEN_181 ? _slots_7_io_uop_ftq_idx : _GEN_137 ? _slots_6_io_uop_ftq_idx : _GEN_123 ? _slots_5_io_uop_ftq_idx : _GEN_106 ? _slots_4_io_uop_ftq_idx : _GEN_86 ? _slots_3_io_uop_ftq_idx : _GEN_111 ? _slots_2_io_uop_ftq_idx : _GEN_36 ? _slots_1_io_uop_ftq_idx : _GEN_13149 ? _slots_0_io_uop_ftq_idx : 6'h0;
  assign io_iss_uops_3_edge_inst = _GEN_594 ? _slots_39_io_uop_edge_inst : _GEN_582 ? _slots_38_io_uop_edge_inst : _GEN_597 ? _slots_37_io_uop_edge_inst : _GEN_557 ? _slots_36_io_uop_edge_inst : _GEN_543 ? _slots_35_io_uop_edge_inst : _GEN_526 ? _slots_34_io_uop_edge_inst : _GEN_512 ? _slots_33_io_uop_edge_inst : _GEN_531 ? _slots_32_io_uop_edge_inst : _GEN_487 ? _slots_31_io_uop_edge_inst : _GEN_473 ? _slots_30_io_uop_edge_inst : _GEN_456 ? _slots_29_io_uop_edge_inst : _GEN_442 ? _slots_28_io_uop_edge_inst : _GEN_461 ? _slots_27_io_uop_edge_inst : _GEN_417 ? _slots_26_io_uop_edge_inst : _GEN_403 ? _slots_25_io_uop_edge_inst : _GEN_386 ? _slots_24_io_uop_edge_inst : _GEN_372 ? _slots_23_io_uop_edge_inst : _GEN_391 ? _slots_22_io_uop_edge_inst : _GEN_347 ? _slots_21_io_uop_edge_inst : _GEN_333 ? _slots_20_io_uop_edge_inst : _GEN_316 ? _slots_19_io_uop_edge_inst : _GEN_302 ? _slots_18_io_uop_edge_inst : _GEN_321 ? _slots_17_io_uop_edge_inst : _GEN_277 ? _slots_16_io_uop_edge_inst : _GEN_263 ? _slots_15_io_uop_edge_inst : _GEN_246 ? _slots_14_io_uop_edge_inst : _GEN_232 ? _slots_13_io_uop_edge_inst : _GEN_251 ? _slots_12_io_uop_edge_inst : _GEN_207 ? _slots_11_io_uop_edge_inst : _GEN_193 ? _slots_10_io_uop_edge_inst : _GEN_176 ? _slots_9_io_uop_edge_inst : _GEN_162 ? _slots_8_io_uop_edge_inst : _GEN_181 ? _slots_7_io_uop_edge_inst : _GEN_137 ? _slots_6_io_uop_edge_inst : _GEN_123 ? _slots_5_io_uop_edge_inst : _GEN_106 ? _slots_4_io_uop_edge_inst : _GEN_86 ? _slots_3_io_uop_edge_inst : _GEN_111 ? _slots_2_io_uop_edge_inst : _GEN_36 ? _slots_1_io_uop_edge_inst : _GEN_13149 & _slots_0_io_uop_edge_inst;
  assign io_iss_uops_3_pc_lob = _GEN_594 ? _slots_39_io_uop_pc_lob : _GEN_582 ? _slots_38_io_uop_pc_lob : _GEN_597 ? _slots_37_io_uop_pc_lob : _GEN_557 ? _slots_36_io_uop_pc_lob : _GEN_543 ? _slots_35_io_uop_pc_lob : _GEN_526 ? _slots_34_io_uop_pc_lob : _GEN_512 ? _slots_33_io_uop_pc_lob : _GEN_531 ? _slots_32_io_uop_pc_lob : _GEN_487 ? _slots_31_io_uop_pc_lob : _GEN_473 ? _slots_30_io_uop_pc_lob : _GEN_456 ? _slots_29_io_uop_pc_lob : _GEN_442 ? _slots_28_io_uop_pc_lob : _GEN_461 ? _slots_27_io_uop_pc_lob : _GEN_417 ? _slots_26_io_uop_pc_lob : _GEN_403 ? _slots_25_io_uop_pc_lob : _GEN_386 ? _slots_24_io_uop_pc_lob : _GEN_372 ? _slots_23_io_uop_pc_lob : _GEN_391 ? _slots_22_io_uop_pc_lob : _GEN_347 ? _slots_21_io_uop_pc_lob : _GEN_333 ? _slots_20_io_uop_pc_lob : _GEN_316 ? _slots_19_io_uop_pc_lob : _GEN_302 ? _slots_18_io_uop_pc_lob : _GEN_321 ? _slots_17_io_uop_pc_lob : _GEN_277 ? _slots_16_io_uop_pc_lob : _GEN_263 ? _slots_15_io_uop_pc_lob : _GEN_246 ? _slots_14_io_uop_pc_lob : _GEN_232 ? _slots_13_io_uop_pc_lob : _GEN_251 ? _slots_12_io_uop_pc_lob : _GEN_207 ? _slots_11_io_uop_pc_lob : _GEN_193 ? _slots_10_io_uop_pc_lob : _GEN_176 ? _slots_9_io_uop_pc_lob : _GEN_162 ? _slots_8_io_uop_pc_lob : _GEN_181 ? _slots_7_io_uop_pc_lob : _GEN_137 ? _slots_6_io_uop_pc_lob : _GEN_123 ? _slots_5_io_uop_pc_lob : _GEN_106 ? _slots_4_io_uop_pc_lob : _GEN_86 ? _slots_3_io_uop_pc_lob : _GEN_111 ? _slots_2_io_uop_pc_lob : _GEN_36 ? _slots_1_io_uop_pc_lob : _GEN_13149 ? _slots_0_io_uop_pc_lob : 6'h0;
  assign io_iss_uops_3_taken = _GEN_594 ? _slots_39_io_uop_taken : _GEN_582 ? _slots_38_io_uop_taken : _GEN_597 ? _slots_37_io_uop_taken : _GEN_557 ? _slots_36_io_uop_taken : _GEN_543 ? _slots_35_io_uop_taken : _GEN_526 ? _slots_34_io_uop_taken : _GEN_512 ? _slots_33_io_uop_taken : _GEN_531 ? _slots_32_io_uop_taken : _GEN_487 ? _slots_31_io_uop_taken : _GEN_473 ? _slots_30_io_uop_taken : _GEN_456 ? _slots_29_io_uop_taken : _GEN_442 ? _slots_28_io_uop_taken : _GEN_461 ? _slots_27_io_uop_taken : _GEN_417 ? _slots_26_io_uop_taken : _GEN_403 ? _slots_25_io_uop_taken : _GEN_386 ? _slots_24_io_uop_taken : _GEN_372 ? _slots_23_io_uop_taken : _GEN_391 ? _slots_22_io_uop_taken : _GEN_347 ? _slots_21_io_uop_taken : _GEN_333 ? _slots_20_io_uop_taken : _GEN_316 ? _slots_19_io_uop_taken : _GEN_302 ? _slots_18_io_uop_taken : _GEN_321 ? _slots_17_io_uop_taken : _GEN_277 ? _slots_16_io_uop_taken : _GEN_263 ? _slots_15_io_uop_taken : _GEN_246 ? _slots_14_io_uop_taken : _GEN_232 ? _slots_13_io_uop_taken : _GEN_251 ? _slots_12_io_uop_taken : _GEN_207 ? _slots_11_io_uop_taken : _GEN_193 ? _slots_10_io_uop_taken : _GEN_176 ? _slots_9_io_uop_taken : _GEN_162 ? _slots_8_io_uop_taken : _GEN_181 ? _slots_7_io_uop_taken : _GEN_137 ? _slots_6_io_uop_taken : _GEN_123 ? _slots_5_io_uop_taken : _GEN_106 ? _slots_4_io_uop_taken : _GEN_86 ? _slots_3_io_uop_taken : _GEN_111 ? _slots_2_io_uop_taken : _GEN_36 ? _slots_1_io_uop_taken : _GEN_13149 & _slots_0_io_uop_taken;
  assign io_iss_uops_3_imm_packed = _GEN_594 ? _slots_39_io_uop_imm_packed : _GEN_582 ? _slots_38_io_uop_imm_packed : _GEN_597 ? _slots_37_io_uop_imm_packed : _GEN_557 ? _slots_36_io_uop_imm_packed : _GEN_543 ? _slots_35_io_uop_imm_packed : _GEN_526 ? _slots_34_io_uop_imm_packed : _GEN_512 ? _slots_33_io_uop_imm_packed : _GEN_531 ? _slots_32_io_uop_imm_packed : _GEN_487 ? _slots_31_io_uop_imm_packed : _GEN_473 ? _slots_30_io_uop_imm_packed : _GEN_456 ? _slots_29_io_uop_imm_packed : _GEN_442 ? _slots_28_io_uop_imm_packed : _GEN_461 ? _slots_27_io_uop_imm_packed : _GEN_417 ? _slots_26_io_uop_imm_packed : _GEN_403 ? _slots_25_io_uop_imm_packed : _GEN_386 ? _slots_24_io_uop_imm_packed : _GEN_372 ? _slots_23_io_uop_imm_packed : _GEN_391 ? _slots_22_io_uop_imm_packed : _GEN_347 ? _slots_21_io_uop_imm_packed : _GEN_333 ? _slots_20_io_uop_imm_packed : _GEN_316 ? _slots_19_io_uop_imm_packed : _GEN_302 ? _slots_18_io_uop_imm_packed : _GEN_321 ? _slots_17_io_uop_imm_packed : _GEN_277 ? _slots_16_io_uop_imm_packed : _GEN_263 ? _slots_15_io_uop_imm_packed : _GEN_246 ? _slots_14_io_uop_imm_packed : _GEN_232 ? _slots_13_io_uop_imm_packed : _GEN_251 ? _slots_12_io_uop_imm_packed : _GEN_207 ? _slots_11_io_uop_imm_packed : _GEN_193 ? _slots_10_io_uop_imm_packed : _GEN_176 ? _slots_9_io_uop_imm_packed : _GEN_162 ? _slots_8_io_uop_imm_packed : _GEN_181 ? _slots_7_io_uop_imm_packed : _GEN_137 ? _slots_6_io_uop_imm_packed : _GEN_123 ? _slots_5_io_uop_imm_packed : _GEN_106 ? _slots_4_io_uop_imm_packed : _GEN_86 ? _slots_3_io_uop_imm_packed : _GEN_111 ? _slots_2_io_uop_imm_packed : _GEN_36 ? _slots_1_io_uop_imm_packed : _GEN_13149 ? _slots_0_io_uop_imm_packed : 20'h0;
  assign io_iss_uops_3_rob_idx = _GEN_594 ? _slots_39_io_uop_rob_idx : _GEN_582 ? _slots_38_io_uop_rob_idx : _GEN_597 ? _slots_37_io_uop_rob_idx : _GEN_557 ? _slots_36_io_uop_rob_idx : _GEN_543 ? _slots_35_io_uop_rob_idx : _GEN_526 ? _slots_34_io_uop_rob_idx : _GEN_512 ? _slots_33_io_uop_rob_idx : _GEN_531 ? _slots_32_io_uop_rob_idx : _GEN_487 ? _slots_31_io_uop_rob_idx : _GEN_473 ? _slots_30_io_uop_rob_idx : _GEN_456 ? _slots_29_io_uop_rob_idx : _GEN_442 ? _slots_28_io_uop_rob_idx : _GEN_461 ? _slots_27_io_uop_rob_idx : _GEN_417 ? _slots_26_io_uop_rob_idx : _GEN_403 ? _slots_25_io_uop_rob_idx : _GEN_386 ? _slots_24_io_uop_rob_idx : _GEN_372 ? _slots_23_io_uop_rob_idx : _GEN_391 ? _slots_22_io_uop_rob_idx : _GEN_347 ? _slots_21_io_uop_rob_idx : _GEN_333 ? _slots_20_io_uop_rob_idx : _GEN_316 ? _slots_19_io_uop_rob_idx : _GEN_302 ? _slots_18_io_uop_rob_idx : _GEN_321 ? _slots_17_io_uop_rob_idx : _GEN_277 ? _slots_16_io_uop_rob_idx : _GEN_263 ? _slots_15_io_uop_rob_idx : _GEN_246 ? _slots_14_io_uop_rob_idx : _GEN_232 ? _slots_13_io_uop_rob_idx : _GEN_251 ? _slots_12_io_uop_rob_idx : _GEN_207 ? _slots_11_io_uop_rob_idx : _GEN_193 ? _slots_10_io_uop_rob_idx : _GEN_176 ? _slots_9_io_uop_rob_idx : _GEN_162 ? _slots_8_io_uop_rob_idx : _GEN_181 ? _slots_7_io_uop_rob_idx : _GEN_137 ? _slots_6_io_uop_rob_idx : _GEN_123 ? _slots_5_io_uop_rob_idx : _GEN_106 ? _slots_4_io_uop_rob_idx : _GEN_86 ? _slots_3_io_uop_rob_idx : _GEN_111 ? _slots_2_io_uop_rob_idx : _GEN_36 ? _slots_1_io_uop_rob_idx : _GEN_13149 ? _slots_0_io_uop_rob_idx : 7'h0;
  assign io_iss_uops_3_ldq_idx = _GEN_594 ? _slots_39_io_uop_ldq_idx : _GEN_582 ? _slots_38_io_uop_ldq_idx : _GEN_597 ? _slots_37_io_uop_ldq_idx : _GEN_557 ? _slots_36_io_uop_ldq_idx : _GEN_543 ? _slots_35_io_uop_ldq_idx : _GEN_526 ? _slots_34_io_uop_ldq_idx : _GEN_512 ? _slots_33_io_uop_ldq_idx : _GEN_531 ? _slots_32_io_uop_ldq_idx : _GEN_487 ? _slots_31_io_uop_ldq_idx : _GEN_473 ? _slots_30_io_uop_ldq_idx : _GEN_456 ? _slots_29_io_uop_ldq_idx : _GEN_442 ? _slots_28_io_uop_ldq_idx : _GEN_461 ? _slots_27_io_uop_ldq_idx : _GEN_417 ? _slots_26_io_uop_ldq_idx : _GEN_403 ? _slots_25_io_uop_ldq_idx : _GEN_386 ? _slots_24_io_uop_ldq_idx : _GEN_372 ? _slots_23_io_uop_ldq_idx : _GEN_391 ? _slots_22_io_uop_ldq_idx : _GEN_347 ? _slots_21_io_uop_ldq_idx : _GEN_333 ? _slots_20_io_uop_ldq_idx : _GEN_316 ? _slots_19_io_uop_ldq_idx : _GEN_302 ? _slots_18_io_uop_ldq_idx : _GEN_321 ? _slots_17_io_uop_ldq_idx : _GEN_277 ? _slots_16_io_uop_ldq_idx : _GEN_263 ? _slots_15_io_uop_ldq_idx : _GEN_246 ? _slots_14_io_uop_ldq_idx : _GEN_232 ? _slots_13_io_uop_ldq_idx : _GEN_251 ? _slots_12_io_uop_ldq_idx : _GEN_207 ? _slots_11_io_uop_ldq_idx : _GEN_193 ? _slots_10_io_uop_ldq_idx : _GEN_176 ? _slots_9_io_uop_ldq_idx : _GEN_162 ? _slots_8_io_uop_ldq_idx : _GEN_181 ? _slots_7_io_uop_ldq_idx : _GEN_137 ? _slots_6_io_uop_ldq_idx : _GEN_123 ? _slots_5_io_uop_ldq_idx : _GEN_106 ? _slots_4_io_uop_ldq_idx : _GEN_86 ? _slots_3_io_uop_ldq_idx : _GEN_111 ? _slots_2_io_uop_ldq_idx : _GEN_36 ? _slots_1_io_uop_ldq_idx : _GEN_13149 ? _slots_0_io_uop_ldq_idx : 5'h0;
  assign io_iss_uops_3_stq_idx = _GEN_594 ? _slots_39_io_uop_stq_idx : _GEN_582 ? _slots_38_io_uop_stq_idx : _GEN_597 ? _slots_37_io_uop_stq_idx : _GEN_557 ? _slots_36_io_uop_stq_idx : _GEN_543 ? _slots_35_io_uop_stq_idx : _GEN_526 ? _slots_34_io_uop_stq_idx : _GEN_512 ? _slots_33_io_uop_stq_idx : _GEN_531 ? _slots_32_io_uop_stq_idx : _GEN_487 ? _slots_31_io_uop_stq_idx : _GEN_473 ? _slots_30_io_uop_stq_idx : _GEN_456 ? _slots_29_io_uop_stq_idx : _GEN_442 ? _slots_28_io_uop_stq_idx : _GEN_461 ? _slots_27_io_uop_stq_idx : _GEN_417 ? _slots_26_io_uop_stq_idx : _GEN_403 ? _slots_25_io_uop_stq_idx : _GEN_386 ? _slots_24_io_uop_stq_idx : _GEN_372 ? _slots_23_io_uop_stq_idx : _GEN_391 ? _slots_22_io_uop_stq_idx : _GEN_347 ? _slots_21_io_uop_stq_idx : _GEN_333 ? _slots_20_io_uop_stq_idx : _GEN_316 ? _slots_19_io_uop_stq_idx : _GEN_302 ? _slots_18_io_uop_stq_idx : _GEN_321 ? _slots_17_io_uop_stq_idx : _GEN_277 ? _slots_16_io_uop_stq_idx : _GEN_263 ? _slots_15_io_uop_stq_idx : _GEN_246 ? _slots_14_io_uop_stq_idx : _GEN_232 ? _slots_13_io_uop_stq_idx : _GEN_251 ? _slots_12_io_uop_stq_idx : _GEN_207 ? _slots_11_io_uop_stq_idx : _GEN_193 ? _slots_10_io_uop_stq_idx : _GEN_176 ? _slots_9_io_uop_stq_idx : _GEN_162 ? _slots_8_io_uop_stq_idx : _GEN_181 ? _slots_7_io_uop_stq_idx : _GEN_137 ? _slots_6_io_uop_stq_idx : _GEN_123 ? _slots_5_io_uop_stq_idx : _GEN_106 ? _slots_4_io_uop_stq_idx : _GEN_86 ? _slots_3_io_uop_stq_idx : _GEN_111 ? _slots_2_io_uop_stq_idx : _GEN_36 ? _slots_1_io_uop_stq_idx : _GEN_13149 ? _slots_0_io_uop_stq_idx : 5'h0;
  assign io_iss_uops_3_pdst = _GEN_594 ? _slots_39_io_uop_pdst : _GEN_582 ? _slots_38_io_uop_pdst : _GEN_597 ? _slots_37_io_uop_pdst : _GEN_557 ? _slots_36_io_uop_pdst : _GEN_543 ? _slots_35_io_uop_pdst : _GEN_526 ? _slots_34_io_uop_pdst : _GEN_512 ? _slots_33_io_uop_pdst : _GEN_531 ? _slots_32_io_uop_pdst : _GEN_487 ? _slots_31_io_uop_pdst : _GEN_473 ? _slots_30_io_uop_pdst : _GEN_456 ? _slots_29_io_uop_pdst : _GEN_442 ? _slots_28_io_uop_pdst : _GEN_461 ? _slots_27_io_uop_pdst : _GEN_417 ? _slots_26_io_uop_pdst : _GEN_403 ? _slots_25_io_uop_pdst : _GEN_386 ? _slots_24_io_uop_pdst : _GEN_372 ? _slots_23_io_uop_pdst : _GEN_391 ? _slots_22_io_uop_pdst : _GEN_347 ? _slots_21_io_uop_pdst : _GEN_333 ? _slots_20_io_uop_pdst : _GEN_316 ? _slots_19_io_uop_pdst : _GEN_302 ? _slots_18_io_uop_pdst : _GEN_321 ? _slots_17_io_uop_pdst : _GEN_277 ? _slots_16_io_uop_pdst : _GEN_263 ? _slots_15_io_uop_pdst : _GEN_246 ? _slots_14_io_uop_pdst : _GEN_232 ? _slots_13_io_uop_pdst : _GEN_251 ? _slots_12_io_uop_pdst : _GEN_207 ? _slots_11_io_uop_pdst : _GEN_193 ? _slots_10_io_uop_pdst : _GEN_176 ? _slots_9_io_uop_pdst : _GEN_162 ? _slots_8_io_uop_pdst : _GEN_181 ? _slots_7_io_uop_pdst : _GEN_137 ? _slots_6_io_uop_pdst : _GEN_123 ? _slots_5_io_uop_pdst : _GEN_106 ? _slots_4_io_uop_pdst : _GEN_86 ? _slots_3_io_uop_pdst : _GEN_111 ? _slots_2_io_uop_pdst : _GEN_36 ? _slots_1_io_uop_pdst : _GEN_13149 ? _slots_0_io_uop_pdst : 7'h0;
  assign io_iss_uops_3_prs1 = _GEN_594 ? _slots_39_io_uop_prs1 : _GEN_582 ? _slots_38_io_uop_prs1 : _GEN_597 ? _slots_37_io_uop_prs1 : _GEN_557 ? _slots_36_io_uop_prs1 : _GEN_543 ? _slots_35_io_uop_prs1 : _GEN_526 ? _slots_34_io_uop_prs1 : _GEN_512 ? _slots_33_io_uop_prs1 : _GEN_531 ? _slots_32_io_uop_prs1 : _GEN_487 ? _slots_31_io_uop_prs1 : _GEN_473 ? _slots_30_io_uop_prs1 : _GEN_456 ? _slots_29_io_uop_prs1 : _GEN_442 ? _slots_28_io_uop_prs1 : _GEN_461 ? _slots_27_io_uop_prs1 : _GEN_417 ? _slots_26_io_uop_prs1 : _GEN_403 ? _slots_25_io_uop_prs1 : _GEN_386 ? _slots_24_io_uop_prs1 : _GEN_372 ? _slots_23_io_uop_prs1 : _GEN_391 ? _slots_22_io_uop_prs1 : _GEN_347 ? _slots_21_io_uop_prs1 : _GEN_333 ? _slots_20_io_uop_prs1 : _GEN_316 ? _slots_19_io_uop_prs1 : _GEN_302 ? _slots_18_io_uop_prs1 : _GEN_321 ? _slots_17_io_uop_prs1 : _GEN_277 ? _slots_16_io_uop_prs1 : _GEN_263 ? _slots_15_io_uop_prs1 : _GEN_246 ? _slots_14_io_uop_prs1 : _GEN_232 ? _slots_13_io_uop_prs1 : _GEN_251 ? _slots_12_io_uop_prs1 : _GEN_207 ? _slots_11_io_uop_prs1 : _GEN_193 ? _slots_10_io_uop_prs1 : _GEN_176 ? _slots_9_io_uop_prs1 : _GEN_162 ? _slots_8_io_uop_prs1 : _GEN_181 ? _slots_7_io_uop_prs1 : _GEN_137 ? _slots_6_io_uop_prs1 : _GEN_123 ? _slots_5_io_uop_prs1 : _GEN_106 ? _slots_4_io_uop_prs1 : _GEN_86 ? _slots_3_io_uop_prs1 : _GEN_111 ? _slots_2_io_uop_prs1 : _GEN_36 ? _slots_1_io_uop_prs1 : _GEN_13149 ? _slots_0_io_uop_prs1 : 7'h0;
  assign io_iss_uops_3_prs2 = _GEN_594 ? _slots_39_io_uop_prs2 : _GEN_582 ? _slots_38_io_uop_prs2 : _GEN_597 ? _slots_37_io_uop_prs2 : _GEN_557 ? _slots_36_io_uop_prs2 : _GEN_543 ? _slots_35_io_uop_prs2 : _GEN_526 ? _slots_34_io_uop_prs2 : _GEN_512 ? _slots_33_io_uop_prs2 : _GEN_531 ? _slots_32_io_uop_prs2 : _GEN_487 ? _slots_31_io_uop_prs2 : _GEN_473 ? _slots_30_io_uop_prs2 : _GEN_456 ? _slots_29_io_uop_prs2 : _GEN_442 ? _slots_28_io_uop_prs2 : _GEN_461 ? _slots_27_io_uop_prs2 : _GEN_417 ? _slots_26_io_uop_prs2 : _GEN_403 ? _slots_25_io_uop_prs2 : _GEN_386 ? _slots_24_io_uop_prs2 : _GEN_372 ? _slots_23_io_uop_prs2 : _GEN_391 ? _slots_22_io_uop_prs2 : _GEN_347 ? _slots_21_io_uop_prs2 : _GEN_333 ? _slots_20_io_uop_prs2 : _GEN_316 ? _slots_19_io_uop_prs2 : _GEN_302 ? _slots_18_io_uop_prs2 : _GEN_321 ? _slots_17_io_uop_prs2 : _GEN_277 ? _slots_16_io_uop_prs2 : _GEN_263 ? _slots_15_io_uop_prs2 : _GEN_246 ? _slots_14_io_uop_prs2 : _GEN_232 ? _slots_13_io_uop_prs2 : _GEN_251 ? _slots_12_io_uop_prs2 : _GEN_207 ? _slots_11_io_uop_prs2 : _GEN_193 ? _slots_10_io_uop_prs2 : _GEN_176 ? _slots_9_io_uop_prs2 : _GEN_162 ? _slots_8_io_uop_prs2 : _GEN_181 ? _slots_7_io_uop_prs2 : _GEN_137 ? _slots_6_io_uop_prs2 : _GEN_123 ? _slots_5_io_uop_prs2 : _GEN_106 ? _slots_4_io_uop_prs2 : _GEN_86 ? _slots_3_io_uop_prs2 : _GEN_111 ? _slots_2_io_uop_prs2 : _GEN_36 ? _slots_1_io_uop_prs2 : _GEN_13149 ? _slots_0_io_uop_prs2 : 7'h0;
  assign io_iss_uops_3_bypassable = _GEN_594 ? _slots_39_io_uop_bypassable : _GEN_582 ? _slots_38_io_uop_bypassable : _GEN_597 ? _slots_37_io_uop_bypassable : _GEN_557 ? _slots_36_io_uop_bypassable : _GEN_543 ? _slots_35_io_uop_bypassable : _GEN_526 ? _slots_34_io_uop_bypassable : _GEN_512 ? _slots_33_io_uop_bypassable : _GEN_531 ? _slots_32_io_uop_bypassable : _GEN_487 ? _slots_31_io_uop_bypassable : _GEN_473 ? _slots_30_io_uop_bypassable : _GEN_456 ? _slots_29_io_uop_bypassable : _GEN_442 ? _slots_28_io_uop_bypassable : _GEN_461 ? _slots_27_io_uop_bypassable : _GEN_417 ? _slots_26_io_uop_bypassable : _GEN_403 ? _slots_25_io_uop_bypassable : _GEN_386 ? _slots_24_io_uop_bypassable : _GEN_372 ? _slots_23_io_uop_bypassable : _GEN_391 ? _slots_22_io_uop_bypassable : _GEN_347 ? _slots_21_io_uop_bypassable : _GEN_333 ? _slots_20_io_uop_bypassable : _GEN_316 ? _slots_19_io_uop_bypassable : _GEN_302 ? _slots_18_io_uop_bypassable : _GEN_321 ? _slots_17_io_uop_bypassable : _GEN_277 ? _slots_16_io_uop_bypassable : _GEN_263 ? _slots_15_io_uop_bypassable : _GEN_246 ? _slots_14_io_uop_bypassable : _GEN_232 ? _slots_13_io_uop_bypassable : _GEN_251 ? _slots_12_io_uop_bypassable : _GEN_207 ? _slots_11_io_uop_bypassable : _GEN_193 ? _slots_10_io_uop_bypassable : _GEN_176 ? _slots_9_io_uop_bypassable : _GEN_162 ? _slots_8_io_uop_bypassable : _GEN_181 ? _slots_7_io_uop_bypassable : _GEN_137 ? _slots_6_io_uop_bypassable : _GEN_123 ? _slots_5_io_uop_bypassable : _GEN_106 ? _slots_4_io_uop_bypassable : _GEN_86 ? _slots_3_io_uop_bypassable : _GEN_111 ? _slots_2_io_uop_bypassable : _GEN_36 ? _slots_1_io_uop_bypassable : _GEN_13149 & _slots_0_io_uop_bypassable;
  assign io_iss_uops_3_mem_cmd = _GEN_594 ? _slots_39_io_uop_mem_cmd : _GEN_582 ? _slots_38_io_uop_mem_cmd : _GEN_597 ? _slots_37_io_uop_mem_cmd : _GEN_557 ? _slots_36_io_uop_mem_cmd : _GEN_543 ? _slots_35_io_uop_mem_cmd : _GEN_526 ? _slots_34_io_uop_mem_cmd : _GEN_512 ? _slots_33_io_uop_mem_cmd : _GEN_531 ? _slots_32_io_uop_mem_cmd : _GEN_487 ? _slots_31_io_uop_mem_cmd : _GEN_473 ? _slots_30_io_uop_mem_cmd : _GEN_456 ? _slots_29_io_uop_mem_cmd : _GEN_442 ? _slots_28_io_uop_mem_cmd : _GEN_461 ? _slots_27_io_uop_mem_cmd : _GEN_417 ? _slots_26_io_uop_mem_cmd : _GEN_403 ? _slots_25_io_uop_mem_cmd : _GEN_386 ? _slots_24_io_uop_mem_cmd : _GEN_372 ? _slots_23_io_uop_mem_cmd : _GEN_391 ? _slots_22_io_uop_mem_cmd : _GEN_347 ? _slots_21_io_uop_mem_cmd : _GEN_333 ? _slots_20_io_uop_mem_cmd : _GEN_316 ? _slots_19_io_uop_mem_cmd : _GEN_302 ? _slots_18_io_uop_mem_cmd : _GEN_321 ? _slots_17_io_uop_mem_cmd : _GEN_277 ? _slots_16_io_uop_mem_cmd : _GEN_263 ? _slots_15_io_uop_mem_cmd : _GEN_246 ? _slots_14_io_uop_mem_cmd : _GEN_232 ? _slots_13_io_uop_mem_cmd : _GEN_251 ? _slots_12_io_uop_mem_cmd : _GEN_207 ? _slots_11_io_uop_mem_cmd : _GEN_193 ? _slots_10_io_uop_mem_cmd : _GEN_176 ? _slots_9_io_uop_mem_cmd : _GEN_162 ? _slots_8_io_uop_mem_cmd : _GEN_181 ? _slots_7_io_uop_mem_cmd : _GEN_137 ? _slots_6_io_uop_mem_cmd : _GEN_123 ? _slots_5_io_uop_mem_cmd : _GEN_106 ? _slots_4_io_uop_mem_cmd : _GEN_86 ? _slots_3_io_uop_mem_cmd : _GEN_111 ? _slots_2_io_uop_mem_cmd : _GEN_36 ? _slots_1_io_uop_mem_cmd : _GEN_13149 ? _slots_0_io_uop_mem_cmd : 5'h0;
  assign io_iss_uops_3_is_amo = _GEN_594 ? _slots_39_io_uop_is_amo : _GEN_582 ? _slots_38_io_uop_is_amo : _GEN_597 ? _slots_37_io_uop_is_amo : _GEN_557 ? _slots_36_io_uop_is_amo : _GEN_543 ? _slots_35_io_uop_is_amo : _GEN_526 ? _slots_34_io_uop_is_amo : _GEN_512 ? _slots_33_io_uop_is_amo : _GEN_531 ? _slots_32_io_uop_is_amo : _GEN_487 ? _slots_31_io_uop_is_amo : _GEN_473 ? _slots_30_io_uop_is_amo : _GEN_456 ? _slots_29_io_uop_is_amo : _GEN_442 ? _slots_28_io_uop_is_amo : _GEN_461 ? _slots_27_io_uop_is_amo : _GEN_417 ? _slots_26_io_uop_is_amo : _GEN_403 ? _slots_25_io_uop_is_amo : _GEN_386 ? _slots_24_io_uop_is_amo : _GEN_372 ? _slots_23_io_uop_is_amo : _GEN_391 ? _slots_22_io_uop_is_amo : _GEN_347 ? _slots_21_io_uop_is_amo : _GEN_333 ? _slots_20_io_uop_is_amo : _GEN_316 ? _slots_19_io_uop_is_amo : _GEN_302 ? _slots_18_io_uop_is_amo : _GEN_321 ? _slots_17_io_uop_is_amo : _GEN_277 ? _slots_16_io_uop_is_amo : _GEN_263 ? _slots_15_io_uop_is_amo : _GEN_246 ? _slots_14_io_uop_is_amo : _GEN_232 ? _slots_13_io_uop_is_amo : _GEN_251 ? _slots_12_io_uop_is_amo : _GEN_207 ? _slots_11_io_uop_is_amo : _GEN_193 ? _slots_10_io_uop_is_amo : _GEN_176 ? _slots_9_io_uop_is_amo : _GEN_162 ? _slots_8_io_uop_is_amo : _GEN_181 ? _slots_7_io_uop_is_amo : _GEN_137 ? _slots_6_io_uop_is_amo : _GEN_123 ? _slots_5_io_uop_is_amo : _GEN_106 ? _slots_4_io_uop_is_amo : _GEN_86 ? _slots_3_io_uop_is_amo : _GEN_111 ? _slots_2_io_uop_is_amo : _GEN_36 ? _slots_1_io_uop_is_amo : _GEN_13149 & _slots_0_io_uop_is_amo;
  assign io_iss_uops_3_uses_stq = _GEN_594 ? _slots_39_io_uop_uses_stq : _GEN_582 ? _slots_38_io_uop_uses_stq : _GEN_597 ? _slots_37_io_uop_uses_stq : _GEN_557 ? _slots_36_io_uop_uses_stq : _GEN_543 ? _slots_35_io_uop_uses_stq : _GEN_526 ? _slots_34_io_uop_uses_stq : _GEN_512 ? _slots_33_io_uop_uses_stq : _GEN_531 ? _slots_32_io_uop_uses_stq : _GEN_487 ? _slots_31_io_uop_uses_stq : _GEN_473 ? _slots_30_io_uop_uses_stq : _GEN_456 ? _slots_29_io_uop_uses_stq : _GEN_442 ? _slots_28_io_uop_uses_stq : _GEN_461 ? _slots_27_io_uop_uses_stq : _GEN_417 ? _slots_26_io_uop_uses_stq : _GEN_403 ? _slots_25_io_uop_uses_stq : _GEN_386 ? _slots_24_io_uop_uses_stq : _GEN_372 ? _slots_23_io_uop_uses_stq : _GEN_391 ? _slots_22_io_uop_uses_stq : _GEN_347 ? _slots_21_io_uop_uses_stq : _GEN_333 ? _slots_20_io_uop_uses_stq : _GEN_316 ? _slots_19_io_uop_uses_stq : _GEN_302 ? _slots_18_io_uop_uses_stq : _GEN_321 ? _slots_17_io_uop_uses_stq : _GEN_277 ? _slots_16_io_uop_uses_stq : _GEN_263 ? _slots_15_io_uop_uses_stq : _GEN_246 ? _slots_14_io_uop_uses_stq : _GEN_232 ? _slots_13_io_uop_uses_stq : _GEN_251 ? _slots_12_io_uop_uses_stq : _GEN_207 ? _slots_11_io_uop_uses_stq : _GEN_193 ? _slots_10_io_uop_uses_stq : _GEN_176 ? _slots_9_io_uop_uses_stq : _GEN_162 ? _slots_8_io_uop_uses_stq : _GEN_181 ? _slots_7_io_uop_uses_stq : _GEN_137 ? _slots_6_io_uop_uses_stq : _GEN_123 ? _slots_5_io_uop_uses_stq : _GEN_106 ? _slots_4_io_uop_uses_stq : _GEN_86 ? _slots_3_io_uop_uses_stq : _GEN_111 ? _slots_2_io_uop_uses_stq : _GEN_36 ? _slots_1_io_uop_uses_stq : _GEN_13149 & _slots_0_io_uop_uses_stq;
  assign io_iss_uops_3_ldst_val = _GEN_594 ? _slots_39_io_uop_ldst_val : _GEN_582 ? _slots_38_io_uop_ldst_val : _GEN_597 ? _slots_37_io_uop_ldst_val : _GEN_557 ? _slots_36_io_uop_ldst_val : _GEN_543 ? _slots_35_io_uop_ldst_val : _GEN_526 ? _slots_34_io_uop_ldst_val : _GEN_512 ? _slots_33_io_uop_ldst_val : _GEN_531 ? _slots_32_io_uop_ldst_val : _GEN_487 ? _slots_31_io_uop_ldst_val : _GEN_473 ? _slots_30_io_uop_ldst_val : _GEN_456 ? _slots_29_io_uop_ldst_val : _GEN_442 ? _slots_28_io_uop_ldst_val : _GEN_461 ? _slots_27_io_uop_ldst_val : _GEN_417 ? _slots_26_io_uop_ldst_val : _GEN_403 ? _slots_25_io_uop_ldst_val : _GEN_386 ? _slots_24_io_uop_ldst_val : _GEN_372 ? _slots_23_io_uop_ldst_val : _GEN_391 ? _slots_22_io_uop_ldst_val : _GEN_347 ? _slots_21_io_uop_ldst_val : _GEN_333 ? _slots_20_io_uop_ldst_val : _GEN_316 ? _slots_19_io_uop_ldst_val : _GEN_302 ? _slots_18_io_uop_ldst_val : _GEN_321 ? _slots_17_io_uop_ldst_val : _GEN_277 ? _slots_16_io_uop_ldst_val : _GEN_263 ? _slots_15_io_uop_ldst_val : _GEN_246 ? _slots_14_io_uop_ldst_val : _GEN_232 ? _slots_13_io_uop_ldst_val : _GEN_251 ? _slots_12_io_uop_ldst_val : _GEN_207 ? _slots_11_io_uop_ldst_val : _GEN_193 ? _slots_10_io_uop_ldst_val : _GEN_176 ? _slots_9_io_uop_ldst_val : _GEN_162 ? _slots_8_io_uop_ldst_val : _GEN_181 ? _slots_7_io_uop_ldst_val : _GEN_137 ? _slots_6_io_uop_ldst_val : _GEN_123 ? _slots_5_io_uop_ldst_val : _GEN_106 ? _slots_4_io_uop_ldst_val : _GEN_86 ? _slots_3_io_uop_ldst_val : _GEN_111 ? _slots_2_io_uop_ldst_val : _GEN_36 ? _slots_1_io_uop_ldst_val : _GEN_13149 & _slots_0_io_uop_ldst_val;
  assign io_iss_uops_3_dst_rtype = _GEN_594 ? _slots_39_io_uop_dst_rtype : _GEN_582 ? _slots_38_io_uop_dst_rtype : _GEN_597 ? _slots_37_io_uop_dst_rtype : _GEN_557 ? _slots_36_io_uop_dst_rtype : _GEN_543 ? _slots_35_io_uop_dst_rtype : _GEN_526 ? _slots_34_io_uop_dst_rtype : _GEN_512 ? _slots_33_io_uop_dst_rtype : _GEN_531 ? _slots_32_io_uop_dst_rtype : _GEN_487 ? _slots_31_io_uop_dst_rtype : _GEN_473 ? _slots_30_io_uop_dst_rtype : _GEN_456 ? _slots_29_io_uop_dst_rtype : _GEN_442 ? _slots_28_io_uop_dst_rtype : _GEN_461 ? _slots_27_io_uop_dst_rtype : _GEN_417 ? _slots_26_io_uop_dst_rtype : _GEN_403 ? _slots_25_io_uop_dst_rtype : _GEN_386 ? _slots_24_io_uop_dst_rtype : _GEN_372 ? _slots_23_io_uop_dst_rtype : _GEN_391 ? _slots_22_io_uop_dst_rtype : _GEN_347 ? _slots_21_io_uop_dst_rtype : _GEN_333 ? _slots_20_io_uop_dst_rtype : _GEN_316 ? _slots_19_io_uop_dst_rtype : _GEN_302 ? _slots_18_io_uop_dst_rtype : _GEN_321 ? _slots_17_io_uop_dst_rtype : _GEN_277 ? _slots_16_io_uop_dst_rtype : _GEN_263 ? _slots_15_io_uop_dst_rtype : _GEN_246 ? _slots_14_io_uop_dst_rtype : _GEN_232 ? _slots_13_io_uop_dst_rtype : _GEN_251 ? _slots_12_io_uop_dst_rtype : _GEN_207 ? _slots_11_io_uop_dst_rtype : _GEN_193 ? _slots_10_io_uop_dst_rtype : _GEN_176 ? _slots_9_io_uop_dst_rtype : _GEN_162 ? _slots_8_io_uop_dst_rtype : _GEN_181 ? _slots_7_io_uop_dst_rtype : _GEN_137 ? _slots_6_io_uop_dst_rtype : _GEN_123 ? _slots_5_io_uop_dst_rtype : _GEN_106 ? _slots_4_io_uop_dst_rtype : _GEN_86 ? _slots_3_io_uop_dst_rtype : _GEN_111 ? _slots_2_io_uop_dst_rtype : _GEN_36 ? _slots_1_io_uop_dst_rtype : _GEN_13149 ? _slots_0_io_uop_dst_rtype : 2'h2;
  assign io_iss_uops_3_lrs1_rtype = _GEN_594 ? _slots_39_io_uop_lrs1_rtype : _GEN_582 ? _slots_38_io_uop_lrs1_rtype : _GEN_597 ? _slots_37_io_uop_lrs1_rtype : _GEN_557 ? _slots_36_io_uop_lrs1_rtype : _GEN_543 ? _slots_35_io_uop_lrs1_rtype : _GEN_526 ? _slots_34_io_uop_lrs1_rtype : _GEN_512 ? _slots_33_io_uop_lrs1_rtype : _GEN_531 ? _slots_32_io_uop_lrs1_rtype : _GEN_487 ? _slots_31_io_uop_lrs1_rtype : _GEN_473 ? _slots_30_io_uop_lrs1_rtype : _GEN_456 ? _slots_29_io_uop_lrs1_rtype : _GEN_442 ? _slots_28_io_uop_lrs1_rtype : _GEN_461 ? _slots_27_io_uop_lrs1_rtype : _GEN_417 ? _slots_26_io_uop_lrs1_rtype : _GEN_403 ? _slots_25_io_uop_lrs1_rtype : _GEN_386 ? _slots_24_io_uop_lrs1_rtype : _GEN_372 ? _slots_23_io_uop_lrs1_rtype : _GEN_391 ? _slots_22_io_uop_lrs1_rtype : _GEN_347 ? _slots_21_io_uop_lrs1_rtype : _GEN_333 ? _slots_20_io_uop_lrs1_rtype : _GEN_316 ? _slots_19_io_uop_lrs1_rtype : _GEN_302 ? _slots_18_io_uop_lrs1_rtype : _GEN_321 ? _slots_17_io_uop_lrs1_rtype : _GEN_277 ? _slots_16_io_uop_lrs1_rtype : _GEN_263 ? _slots_15_io_uop_lrs1_rtype : _GEN_246 ? _slots_14_io_uop_lrs1_rtype : _GEN_232 ? _slots_13_io_uop_lrs1_rtype : _GEN_251 ? _slots_12_io_uop_lrs1_rtype : _GEN_207 ? _slots_11_io_uop_lrs1_rtype : _GEN_193 ? _slots_10_io_uop_lrs1_rtype : _GEN_176 ? _slots_9_io_uop_lrs1_rtype : _GEN_162 ? _slots_8_io_uop_lrs1_rtype : _GEN_181 ? _slots_7_io_uop_lrs1_rtype : _GEN_137 ? _slots_6_io_uop_lrs1_rtype : _GEN_123 ? _slots_5_io_uop_lrs1_rtype : _GEN_106 ? _slots_4_io_uop_lrs1_rtype : _GEN_86 ? _slots_3_io_uop_lrs1_rtype : _GEN_111 ? _slots_2_io_uop_lrs1_rtype : _GEN_36 ? _slots_1_io_uop_lrs1_rtype : _GEN_13149 ? _slots_0_io_uop_lrs1_rtype : 2'h2;
  assign io_iss_uops_3_lrs2_rtype = _GEN_594 ? _slots_39_io_uop_lrs2_rtype : _GEN_582 ? _slots_38_io_uop_lrs2_rtype : _GEN_597 ? _slots_37_io_uop_lrs2_rtype : _GEN_557 ? _slots_36_io_uop_lrs2_rtype : _GEN_543 ? _slots_35_io_uop_lrs2_rtype : _GEN_526 ? _slots_34_io_uop_lrs2_rtype : _GEN_512 ? _slots_33_io_uop_lrs2_rtype : _GEN_531 ? _slots_32_io_uop_lrs2_rtype : _GEN_487 ? _slots_31_io_uop_lrs2_rtype : _GEN_473 ? _slots_30_io_uop_lrs2_rtype : _GEN_456 ? _slots_29_io_uop_lrs2_rtype : _GEN_442 ? _slots_28_io_uop_lrs2_rtype : _GEN_461 ? _slots_27_io_uop_lrs2_rtype : _GEN_417 ? _slots_26_io_uop_lrs2_rtype : _GEN_403 ? _slots_25_io_uop_lrs2_rtype : _GEN_386 ? _slots_24_io_uop_lrs2_rtype : _GEN_372 ? _slots_23_io_uop_lrs2_rtype : _GEN_391 ? _slots_22_io_uop_lrs2_rtype : _GEN_347 ? _slots_21_io_uop_lrs2_rtype : _GEN_333 ? _slots_20_io_uop_lrs2_rtype : _GEN_316 ? _slots_19_io_uop_lrs2_rtype : _GEN_302 ? _slots_18_io_uop_lrs2_rtype : _GEN_321 ? _slots_17_io_uop_lrs2_rtype : _GEN_277 ? _slots_16_io_uop_lrs2_rtype : _GEN_263 ? _slots_15_io_uop_lrs2_rtype : _GEN_246 ? _slots_14_io_uop_lrs2_rtype : _GEN_232 ? _slots_13_io_uop_lrs2_rtype : _GEN_251 ? _slots_12_io_uop_lrs2_rtype : _GEN_207 ? _slots_11_io_uop_lrs2_rtype : _GEN_193 ? _slots_10_io_uop_lrs2_rtype : _GEN_176 ? _slots_9_io_uop_lrs2_rtype : _GEN_162 ? _slots_8_io_uop_lrs2_rtype : _GEN_181 ? _slots_7_io_uop_lrs2_rtype : _GEN_137 ? _slots_6_io_uop_lrs2_rtype : _GEN_123 ? _slots_5_io_uop_lrs2_rtype : _GEN_106 ? _slots_4_io_uop_lrs2_rtype : _GEN_86 ? _slots_3_io_uop_lrs2_rtype : _GEN_111 ? _slots_2_io_uop_lrs2_rtype : _GEN_36 ? _slots_1_io_uop_lrs2_rtype : _GEN_13149 ? _slots_0_io_uop_lrs2_rtype : 2'h2;
endmodule

