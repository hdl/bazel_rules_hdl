// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// VCS coverage exclude_file
module Rob_assert(
  input [4:0] rob_tail,
  input       rob_val__31,
              rob_val__30,
              rob_val__29,
              rob_val__28,
              rob_val__27,
              rob_val__26,
              rob_val__25,
              rob_val__24,
              rob_val__23,
              rob_val__22,
              rob_val__21,
              rob_val__20,
              rob_val__19,
              rob_val__18,
              rob_val__17,
              rob_val__16,
              rob_val__15,
              rob_val__14,
              rob_val__13,
              rob_val__12,
              rob_val__11,
              rob_val__10,
              rob_val__9,
              rob_val__8,
              rob_val__7,
              rob_val__6,
              rob_val__5,
              rob_val__4,
              rob_val__3,
              rob_val__2,
              rob_val__1,
              rob_val__0,
  input [6:0] io_enq_uops_0_rob_idx,
  input [4:0] _GEN,
  input       rob_bsy__31,
              rob_bsy__30,
              rob_bsy__29,
              rob_bsy__28,
              rob_bsy__27,
              rob_bsy__26,
              rob_bsy__25,
              rob_bsy__24,
              rob_bsy__23,
              rob_bsy__22,
              rob_bsy__21,
              rob_bsy__20,
              rob_bsy__19,
              rob_bsy__18,
              rob_bsy__17,
              rob_bsy__16,
              rob_bsy__15,
              rob_bsy__14,
              rob_bsy__13,
              rob_bsy__12,
              rob_bsy__11,
              rob_bsy__10,
              rob_bsy__9,
              rob_bsy__8,
              rob_bsy__7,
              rob_bsy__6,
              rob_bsy__5,
              rob_bsy__4,
              rob_bsy__3,
              rob_bsy__2,
              rob_bsy__1,
              rob_bsy__0,
  input [4:0] _GEN_0,
              _GEN_1,
              _GEN_2,
  input       clock,
              _GEN_3,
              _GEN_4,
              _GEN_5,
              _GEN_6,
              _GEN_7,
              _GEN_8,
              _GEN_9,
              io_enq_uops_0_uses_ldq,
              io_enq_uops_0_is_br,
              io_enq_uops_0_is_jalr,
              io_enq_uops_0_uses_stq,
              io_enq_uops_0_is_fence,
              _GEN_10,
              _GEN_11,
              _GEN_12,
              _GEN_13,
              _GEN_14,
              _GEN_15,
              _GEN_16,
              _GEN_17,
              _GEN_18,
              _GEN_19,
              _GEN_20,
              _GEN_21,
              _GEN_22,
              _GEN_23,
              _GEN_24,
              _GEN_25,
              _GEN_26,
              _GEN_27,
              _GEN_28,
              _GEN_29,
              _GEN_30,
              _GEN_31,
              _GEN_32,
              _GEN_33,
              _GEN_34,
              _GEN_35,
              _GEN_36,
              _GEN_37,
              _GEN_38,
              _GEN_39,
              _GEN_40,
              _GEN_41,
              _GEN_42,
              _GEN_43,
              _GEN_44,
              _GEN_45,
              _GEN_46,
              _GEN_47,
              _GEN_48,
              _GEN_49,
              _GEN_50,
              _GEN_51,
              _GEN_52,
              _GEN_53,
              _GEN_54,
              _GEN_55,
              _GEN_56,
              _GEN_57,
              _GEN_58,
              _GEN_59,
              _GEN_60,
              _GEN_61,
              _GEN_62,
              _GEN_63,
              _GEN_64,
              _GEN_65,
              _GEN_66,
              _GEN_67,
              _GEN_68,
              _GEN_69,
              _GEN_70,
              _GEN_71,
              _GEN_72,
              _GEN_73,
              _GEN_74,
              _GEN_75,
              _GEN_76,
              _GEN_77,
              _GEN_78,
              _GEN_79,
              _GEN_80,
              _GEN_81,
              _GEN_82,
              _GEN_83,
              _GEN_84,
              _GEN_85,
              _GEN_86,
              _GEN_87,
              _GEN_88,
              _GEN_89,
              _GEN_90,
              _GEN_91,
              _GEN_92,
              _GEN_93,
              _GEN_94,
              _GEN_95,
              _GEN_96,
              _GEN_97,
              _GEN_98,
              _GEN_99,
              _GEN_100,
              _GEN_101,
              _GEN_102,
              _GEN_103,
              _GEN_104,
              _GEN_105,
              _GEN_106,
              _GEN_107,
              _GEN_108,
              _GEN_109,
              _GEN_110,
              _GEN_111,
              _GEN_112,
              _GEN_113,
              _GEN_114,
              _GEN_115,
              _GEN_116,
              _GEN_117,
              _GEN_118,
              _GEN_119,
              _GEN_120,
              _GEN_121,
              _GEN_122,
              _GEN_123,
              _GEN_124,
              _GEN_125,
              _GEN_126,
              _GEN_127,
              _GEN_128,
              _GEN_129,
              _GEN_130,
              _GEN_131,
              _GEN_132,
              _GEN_133,
              _GEN_134,
              _GEN_135,
              _GEN_136,
              _GEN_137,
              _GEN_138,
              _GEN_139,
              _GEN_140,
              _GEN_141,
              _GEN_142,
              _GEN_143,
              _GEN_144,
              _GEN_145,
              _GEN_146,
              _GEN_147,
              _GEN_148,
              _GEN_149,
              _GEN_150,
              _GEN_151,
              _GEN_152,
              _GEN_153,
              _GEN_154,
              _GEN_155,
              _GEN_156,
              _GEN_157,
              _GEN_158,
              _GEN_159,
              _GEN_160,
              _GEN_161,
              _GEN_162,
              _GEN_163,
              _GEN_164,
              _GEN_165,
              _GEN_166,
              _GEN_167,
              _GEN_168,
              _GEN_169,
              _GEN_170,
              _GEN_171,
              _GEN_172,
              _GEN_173,
              _GEN_174,
              _GEN_175,
              _GEN_176,
              _GEN_177,
              _GEN_178,
              _GEN_179,
              _GEN_180,
              _GEN_181,
              _GEN_182,
              _GEN_183,
              _GEN_184,
              _GEN_185,
              _GEN_186,
              _GEN_187,
              _GEN_188,
              _GEN_189,
              _GEN_190,
              _GEN_191,
              _GEN_192,
              _GEN_193,
              _GEN_194,
              _GEN_195,
              _GEN_196,
              _GEN_197,
              _GEN_198,
              _GEN_199,
              _GEN_200,
              _GEN_201,
              _GEN_202,
              _GEN_203,
              _GEN_204,
              _GEN_205,
              _GEN_206,
              _GEN_207,
              _GEN_208,
              _GEN_209,
              _GEN_210,
              _GEN_211,
              _GEN_212,
              _GEN_213,
              _GEN_214,
              _GEN_215,
              _GEN_216,
              _GEN_217,
              _GEN_218,
              _GEN_219,
              _GEN_220,
              _GEN_221,
              _GEN_222,
              _GEN_223,
              _GEN_224,
              _GEN_225,
              _GEN_226,
              _GEN_227,
              _GEN_228,
              _GEN_229,
              _GEN_230,
              _GEN_231,
              _GEN_232,
              _GEN_233,
              _GEN_234,
              _GEN_235,
              _GEN_236,
              _GEN_237,
              _GEN_238,
              _GEN_239,
              _GEN_240,
              _GEN_241,
              _GEN_242,
              _GEN_243,
              _GEN_244,
              _GEN_245,
              _GEN_246,
              _GEN_247,
              _GEN_248,
              _GEN_249,
              _GEN_250,
              _GEN_251,
              _GEN_252,
              _GEN_253,
              _GEN_254,
              _GEN_255,
              _GEN_256,
              _GEN_257,
              _GEN_258,
              _GEN_259,
              _GEN_260,
              _GEN_261,
              _GEN_262,
              _GEN_263,
              _GEN_264,
              _GEN_265,
              _GEN_266,
              _GEN_267,
              _GEN_268,
              _GEN_269,
              _GEN_270,
              _GEN_271,
              _GEN_272,
              _GEN_273,
              _GEN_274,
              _GEN_275,
              _GEN_276,
              _GEN_277,
              _GEN_278,
              _GEN_279,
              _GEN_280,
              _GEN_281,
              _GEN_282,
              _GEN_283,
              _GEN_284,
              _GEN_285,
              _GEN_286,
              _GEN_287,
              _GEN_288,
              _GEN_289,
              _GEN_290,
              _GEN_291,
              _GEN_292,
              _GEN_293,
              _GEN_294,
              _GEN_295,
              _GEN_296,
              _GEN_297,
              _GEN_298,
              _GEN_299,
              _GEN_300,
              _GEN_301,
              _GEN_302,
              _GEN_303,
              _GEN_304,
              _GEN_305,
              _GEN_306,
              _GEN_307,
              _GEN_308,
              _GEN_309,
              _GEN_310,
              _GEN_311,
              _GEN_312,
              _GEN_313,
              _GEN_314,
              _GEN_315,
              _GEN_316,
              _GEN_317,
              _GEN_318,
              _GEN_319,
              _GEN_320,
              _GEN_321,
              _GEN_322,
              _GEN_323,
              _GEN_324,
              _GEN_325,
              _GEN_326,
              _GEN_327,
              _GEN_328,
              _GEN_329,
              _GEN_330,
              _GEN_331,
              _GEN_332,
              _GEN_333,
              _GEN_334,
              _GEN_335,
              _GEN_336,
              _GEN_337,
              _GEN_338,
              _GEN_339,
              _GEN_340,
              _GEN_341,
              _GEN_342,
              _GEN_343,
              _GEN_344,
              _GEN_345,
              _GEN_346,
              _GEN_347,
              _GEN_348,
              _GEN_349,
              _GEN_350,
              _GEN_351,
              _GEN_352,
              _GEN_353,
              _GEN_354,
              _GEN_355,
              _GEN_356,
              _GEN_357,
              _GEN_358,
              _GEN_359,
              _GEN_360,
              _GEN_361,
              _GEN_362,
              _GEN_363,
              _GEN_364,
              _GEN_365,
              _GEN_366,
              _GEN_367,
              _GEN_368,
              _GEN_369,
              _GEN_370,
              _GEN_371,
              _GEN_372,
              _GEN_373,
              _GEN_374,
              _GEN_375,
              _GEN_376,
              _GEN_377,
              _GEN_378,
              _GEN_379,
              _GEN_380,
              _GEN_381,
              _GEN_382,
              _GEN_383,
              _GEN_384,
              _GEN_385,
              _GEN_386,
              _GEN_387,
              _GEN_388,
              _GEN_389,
              _GEN_390,
              _GEN_391,
              _GEN_392,
              _GEN_393,
              _GEN_394,
              _GEN_395,
              _GEN_396,
              _GEN_397,
              _GEN_398,
              _GEN_399,
              _GEN_400,
              _GEN_401,
              _GEN_402,
              _GEN_403,
              _GEN_404,
              _GEN_405,
              _GEN_406,
              _GEN_407,
              _GEN_408,
              _GEN_409,
              _GEN_410,
              _GEN_411,
              _GEN_412,
              _GEN_413,
              _GEN_414,
              _GEN_415,
              _GEN_416,
              _GEN_417,
              _GEN_418,
              _GEN_419,
              _GEN_420,
              _GEN_421,
              _GEN_422,
              _GEN_423,
              _GEN_424,
              _GEN_425,
              _GEN_426,
              _GEN_427,
              _GEN_428,
              _GEN_429,
              _GEN_430,
              _GEN_431,
              _GEN_432,
              _GEN_433,
              _GEN_434,
              _GEN_435,
              _GEN_436,
              _GEN_437,
              _GEN_438,
              _GEN_439,
              _GEN_440,
              _GEN_441,
              _GEN_442,
              _GEN_443,
              _GEN_444,
              _GEN_445,
              _GEN_446,
              _GEN_447,
              _GEN_448,
              _GEN_449,
              _GEN_450,
              _GEN_451,
              _GEN_452,
              _GEN_453,
              _GEN_454,
              _GEN_455,
              _GEN_456,
              _io_commit_rbk_valids_0_output,
              _io_commit_rbk_valids_1_output,
              _io_commit_rbk_valids_2_output,
              _io_commit_rbk_valids_3_output,
              _io_commit_valids_0_output,
              _io_commit_valids_1_output,
              _io_commit_valids_2_output,
              _io_commit_valids_3_output,
              _GEN_457,
  input [4:0] _temp_uop_T_61,
  input [6:0] io_wb_resps_0_bits_uop_pdst,
              rob_uop__31_pdst,
              rob_uop__30_pdst,
              rob_uop__29_pdst,
              rob_uop__28_pdst,
              rob_uop__27_pdst,
              rob_uop__26_pdst,
              rob_uop__25_pdst,
              rob_uop__24_pdst,
              rob_uop__23_pdst,
              rob_uop__22_pdst,
              rob_uop__21_pdst,
              rob_uop__20_pdst,
              rob_uop__19_pdst,
              rob_uop__18_pdst,
              rob_uop__17_pdst,
              rob_uop__16_pdst,
              rob_uop__15_pdst,
              rob_uop__14_pdst,
              rob_uop__13_pdst,
              rob_uop__12_pdst,
              rob_uop__11_pdst,
              rob_uop__10_pdst,
              rob_uop__9_pdst,
              rob_uop__8_pdst,
              rob_uop__7_pdst,
              rob_uop__6_pdst,
              rob_uop__5_pdst,
              rob_uop__4_pdst,
              rob_uop__3_pdst,
              rob_uop__2_pdst,
              rob_uop__1_pdst,
              rob_uop__0_pdst,
  input       rob_uop__31_ldst_val,
              rob_uop__30_ldst_val,
              rob_uop__29_ldst_val,
              rob_uop__28_ldst_val,
              rob_uop__27_ldst_val,
              rob_uop__26_ldst_val,
              rob_uop__25_ldst_val,
              rob_uop__24_ldst_val,
              rob_uop__23_ldst_val,
              rob_uop__22_ldst_val,
              rob_uop__21_ldst_val,
              rob_uop__20_ldst_val,
              rob_uop__19_ldst_val,
              rob_uop__18_ldst_val,
              rob_uop__17_ldst_val,
              rob_uop__16_ldst_val,
              rob_uop__15_ldst_val,
              rob_uop__14_ldst_val,
              rob_uop__13_ldst_val,
              rob_uop__12_ldst_val,
              rob_uop__11_ldst_val,
              rob_uop__10_ldst_val,
              rob_uop__9_ldst_val,
              rob_uop__8_ldst_val,
              rob_uop__7_ldst_val,
              rob_uop__6_ldst_val,
              rob_uop__5_ldst_val,
              rob_uop__4_ldst_val,
              rob_uop__3_ldst_val,
              rob_uop__2_ldst_val,
              rob_uop__1_ldst_val,
              rob_uop__0_ldst_val,
  input [4:0] _temp_uop_T_63,
  input [6:0] io_wb_resps_1_bits_uop_pdst,
  input       _GEN_458,
  input [4:0] _temp_uop_T_65,
  input [6:0] io_wb_resps_2_bits_uop_pdst,
  input [4:0] _temp_uop_T_67,
  input [6:0] io_wb_resps_3_bits_uop_pdst,
  input       _GEN_459,
  input [4:0] _temp_uop_T_69,
  input [6:0] io_wb_resps_4_bits_uop_pdst,
  input [4:0] _temp_uop_T_71,
  input [6:0] io_wb_resps_5_bits_uop_pdst,
  input       _GEN_460,
  input [4:0] _temp_uop_T_73,
  input [6:0] io_wb_resps_6_bits_uop_pdst,
  input [4:0] _temp_uop_T_75,
  input [6:0] io_wb_resps_7_bits_uop_pdst,
  input       _GEN_461,
  input [4:0] _temp_uop_T_77,
  input [6:0] io_wb_resps_8_bits_uop_pdst,
  input [4:0] _temp_uop_T_79,
  input [6:0] io_wb_resps_9_bits_uop_pdst,
  input       rob_val_1_31,
              rob_val_1_30,
              rob_val_1_29,
              rob_val_1_28,
              rob_val_1_27,
              rob_val_1_26,
              rob_val_1_25,
              rob_val_1_24,
              rob_val_1_23,
              rob_val_1_22,
              rob_val_1_21,
              rob_val_1_20,
              rob_val_1_19,
              rob_val_1_18,
              rob_val_1_17,
              rob_val_1_16,
              rob_val_1_15,
              rob_val_1_14,
              rob_val_1_13,
              rob_val_1_12,
              rob_val_1_11,
              rob_val_1_10,
              rob_val_1_9,
              rob_val_1_8,
              rob_val_1_7,
              rob_val_1_6,
              rob_val_1_5,
              rob_val_1_4,
              rob_val_1_3,
              rob_val_1_2,
              rob_val_1_1,
              rob_val_1_0,
  input [6:0] io_enq_uops_1_rob_idx,
  input       rob_bsy_1_31,
              rob_bsy_1_30,
              rob_bsy_1_29,
              rob_bsy_1_28,
              rob_bsy_1_27,
              rob_bsy_1_26,
              rob_bsy_1_25,
              rob_bsy_1_24,
              rob_bsy_1_23,
              rob_bsy_1_22,
              rob_bsy_1_21,
              rob_bsy_1_20,
              rob_bsy_1_19,
              rob_bsy_1_18,
              rob_bsy_1_17,
              rob_bsy_1_16,
              rob_bsy_1_15,
              rob_bsy_1_14,
              rob_bsy_1_13,
              rob_bsy_1_12,
              rob_bsy_1_11,
              rob_bsy_1_10,
              rob_bsy_1_9,
              rob_bsy_1_8,
              rob_bsy_1_7,
              rob_bsy_1_6,
              rob_bsy_1_5,
              rob_bsy_1_4,
              rob_bsy_1_3,
              rob_bsy_1_2,
              rob_bsy_1_1,
              rob_bsy_1_0,
              _GEN_462,
              _GEN_463,
              _GEN_464,
              _GEN_465,
              _GEN_466,
              _GEN_467,
              _GEN_468,
              io_enq_uops_1_uses_ldq,
              io_enq_uops_1_is_br,
              io_enq_uops_1_is_jalr,
              io_enq_uops_1_uses_stq,
              io_enq_uops_1_is_fence,
              _GEN_469,
              _GEN_470,
              _GEN_471,
              _GEN_472,
              _GEN_473,
              _GEN_474,
              _GEN_475,
              _GEN_476,
              _GEN_477,
              _GEN_478,
              _GEN_479,
              _GEN_480,
              _GEN_481,
              _GEN_482,
              _GEN_483,
              _GEN_484,
              _GEN_485,
              _GEN_486,
              _GEN_487,
              _GEN_488,
              _GEN_489,
              _GEN_490,
              _GEN_491,
              _GEN_492,
              _GEN_493,
              _GEN_494,
              _GEN_495,
              _GEN_496,
              _GEN_497,
              _GEN_498,
              _GEN_499,
              _GEN_500,
              _GEN_501,
              _GEN_502,
              _GEN_503,
              _GEN_504,
              _GEN_505,
              _GEN_506,
              _GEN_507,
              _GEN_508,
              _GEN_509,
              _GEN_510,
              _GEN_511,
              _GEN_512,
              _GEN_513,
              _GEN_514,
              _GEN_515,
              _GEN_516,
              _GEN_517,
              _GEN_518,
              _GEN_519,
              _GEN_520,
              _GEN_521,
              _GEN_522,
              _GEN_523,
              _GEN_524,
              _GEN_525,
              _GEN_526,
              _GEN_527,
              _GEN_528,
              _GEN_529,
              _GEN_530,
              _GEN_531,
              _GEN_532,
              _GEN_533,
              _GEN_534,
              _GEN_535,
              _GEN_536,
              _GEN_537,
              _GEN_538,
              _GEN_539,
              _GEN_540,
              _GEN_541,
              _GEN_542,
              _GEN_543,
              _GEN_544,
              _GEN_545,
              _GEN_546,
              _GEN_547,
              _GEN_548,
              _GEN_549,
              _GEN_550,
              _GEN_551,
              _GEN_552,
              _GEN_553,
              _GEN_554,
              _GEN_555,
              _GEN_556,
              _GEN_557,
              _GEN_558,
              _GEN_559,
              _GEN_560,
              _GEN_561,
              _GEN_562,
              _GEN_563,
              _GEN_564,
              _GEN_565,
              _GEN_566,
              _GEN_567,
              _GEN_568,
              _GEN_569,
              _GEN_570,
              _GEN_571,
              _GEN_572,
              _GEN_573,
              _GEN_574,
              _GEN_575,
              _GEN_576,
              _GEN_577,
              _GEN_578,
              _GEN_579,
              _GEN_580,
              _GEN_581,
              _GEN_582,
              _GEN_583,
              _GEN_584,
              _GEN_585,
              _GEN_586,
              _GEN_587,
              _GEN_588,
              _GEN_589,
              _GEN_590,
              _GEN_591,
              _GEN_592,
              _GEN_593,
              _GEN_594,
              _GEN_595,
              _GEN_596,
              _GEN_597,
              _GEN_598,
              _GEN_599,
              _GEN_600,
              _GEN_601,
              _GEN_602,
              _GEN_603,
              _GEN_604,
              _GEN_605,
              _GEN_606,
              _GEN_607,
              _GEN_608,
              _GEN_609,
              _GEN_610,
              _GEN_611,
              _GEN_612,
              _GEN_613,
              _GEN_614,
              _GEN_615,
              _GEN_616,
              _GEN_617,
              _GEN_618,
              _GEN_619,
              _GEN_620,
              _GEN_621,
              _GEN_622,
              _GEN_623,
              _GEN_624,
              _GEN_625,
              _GEN_626,
              _GEN_627,
              _GEN_628,
              _GEN_629,
              _GEN_630,
              _GEN_631,
              _GEN_632,
              _GEN_633,
              _GEN_634,
              _GEN_635,
              _GEN_636,
              _GEN_637,
              _GEN_638,
              _GEN_639,
              _GEN_640,
              _GEN_641,
              _GEN_642,
              _GEN_643,
              _GEN_644,
              _GEN_645,
              _GEN_646,
              _GEN_647,
              _GEN_648,
              _GEN_649,
              _GEN_650,
              _GEN_651,
              _GEN_652,
              _GEN_653,
              _GEN_654,
              _GEN_655,
              _GEN_656,
              _GEN_657,
              _GEN_658,
              _GEN_659,
              _GEN_660,
              _GEN_661,
              _GEN_662,
              _GEN_663,
              _GEN_664,
              _GEN_665,
              _GEN_666,
              _GEN_667,
              _GEN_668,
              _GEN_669,
              _GEN_670,
              _GEN_671,
              _GEN_672,
              _GEN_673,
              _GEN_674,
              _GEN_675,
              _GEN_676,
              _GEN_677,
              _GEN_678,
              _GEN_679,
              _GEN_680,
              _GEN_681,
              _GEN_682,
              _GEN_683,
              _GEN_684,
              _GEN_685,
              _GEN_686,
              _GEN_687,
              _GEN_688,
              _GEN_689,
              _GEN_690,
              _GEN_691,
              _GEN_692,
              _GEN_693,
              _GEN_694,
              _GEN_695,
              _GEN_696,
              _GEN_697,
              _GEN_698,
              _GEN_699,
              _GEN_700,
              _GEN_701,
              _GEN_702,
              _GEN_703,
              _GEN_704,
              _GEN_705,
              _GEN_706,
              _GEN_707,
              _GEN_708,
              _GEN_709,
              _GEN_710,
              _GEN_711,
              _GEN_712,
              _GEN_713,
              _GEN_714,
              _GEN_715,
              _GEN_716,
              _GEN_717,
              _GEN_718,
              _GEN_719,
              _GEN_720,
              _GEN_721,
              _GEN_722,
              _GEN_723,
              _GEN_724,
              _GEN_725,
              _GEN_726,
              _GEN_727,
              _GEN_728,
              _GEN_729,
              _GEN_730,
              _GEN_731,
              _GEN_732,
              _GEN_733,
              _GEN_734,
              _GEN_735,
              _GEN_736,
              _GEN_737,
              _GEN_738,
              _GEN_739,
              _GEN_740,
              _GEN_741,
              _GEN_742,
              _GEN_743,
              _GEN_744,
              _GEN_745,
              _GEN_746,
              _GEN_747,
              _GEN_748,
              _GEN_749,
              _GEN_750,
              _GEN_751,
              _GEN_752,
              _GEN_753,
              _GEN_754,
              _GEN_755,
              _GEN_756,
              _GEN_757,
              _GEN_758,
              _GEN_759,
              _GEN_760,
              _GEN_761,
              _GEN_762,
              _GEN_763,
              _GEN_764,
              _GEN_765,
              _GEN_766,
              _GEN_767,
              _GEN_768,
              _GEN_769,
              _GEN_770,
              _GEN_771,
              _GEN_772,
              _GEN_773,
              _GEN_774,
              _GEN_775,
              _GEN_776,
              _GEN_777,
              _GEN_778,
              _GEN_779,
              _GEN_780,
              _GEN_781,
              _GEN_782,
              _GEN_783,
              _GEN_784,
              _GEN_785,
              _GEN_786,
              _GEN_787,
              _GEN_788,
              _GEN_789,
              _GEN_790,
              _GEN_791,
              _GEN_792,
              _GEN_793,
              _GEN_794,
              _GEN_795,
              _GEN_796,
              _GEN_797,
              _GEN_798,
              _GEN_799,
              _GEN_800,
              _GEN_801,
              _GEN_802,
              _GEN_803,
              _GEN_804,
              _GEN_805,
              _GEN_806,
              _GEN_807,
              _GEN_808,
              _GEN_809,
              _GEN_810,
              _GEN_811,
              _GEN_812,
              _GEN_813,
              _GEN_814,
              _GEN_815,
              _GEN_816,
              _GEN_817,
              _GEN_818,
              _GEN_819,
              _GEN_820,
              _GEN_821,
              _GEN_822,
              _GEN_823,
              _GEN_824,
              _GEN_825,
              _GEN_826,
              _GEN_827,
              _GEN_828,
              _GEN_829,
              _GEN_830,
              _GEN_831,
              _GEN_832,
              _GEN_833,
              _GEN_834,
              _GEN_835,
              _GEN_836,
              _GEN_837,
              _GEN_838,
              _GEN_839,
              _GEN_840,
              _GEN_841,
              _GEN_842,
              _GEN_843,
              _GEN_844,
              _GEN_845,
              _GEN_846,
              _GEN_847,
              _GEN_848,
              _GEN_849,
              _GEN_850,
              _GEN_851,
              _GEN_852,
              _GEN_853,
              _GEN_854,
              _GEN_855,
              _GEN_856,
              _GEN_857,
              _GEN_858,
              _GEN_859,
              _GEN_860,
              _GEN_861,
              _GEN_862,
              _GEN_863,
              _GEN_864,
              _GEN_865,
              _GEN_866,
              _GEN_867,
              _GEN_868,
              _GEN_869,
              _GEN_870,
              _GEN_871,
              _GEN_872,
              _GEN_873,
              _GEN_874,
              _GEN_875,
              _GEN_876,
              _GEN_877,
              _GEN_878,
              _GEN_879,
              _GEN_880,
              _GEN_881,
              _GEN_882,
              _GEN_883,
              _GEN_884,
              _GEN_885,
              _GEN_886,
              _GEN_887,
              _GEN_888,
              _GEN_889,
              _GEN_890,
              _GEN_891,
              _GEN_892,
              _GEN_893,
              _GEN_894,
              _GEN_895,
              _GEN_896,
              _GEN_897,
              _GEN_898,
              _GEN_899,
              _GEN_900,
              _GEN_901,
              _GEN_902,
              _GEN_903,
              _GEN_904,
              _GEN_905,
              _GEN_906,
              _GEN_907,
              _GEN_908,
              _GEN_909,
              _GEN_910,
              _GEN_911,
              _GEN_912,
              _GEN_913,
              _GEN_914,
              _GEN_915,
              _GEN_916,
  input [6:0] rob_uop_1_31_pdst,
              rob_uop_1_30_pdst,
              rob_uop_1_29_pdst,
              rob_uop_1_28_pdst,
              rob_uop_1_27_pdst,
              rob_uop_1_26_pdst,
              rob_uop_1_25_pdst,
              rob_uop_1_24_pdst,
              rob_uop_1_23_pdst,
              rob_uop_1_22_pdst,
              rob_uop_1_21_pdst,
              rob_uop_1_20_pdst,
              rob_uop_1_19_pdst,
              rob_uop_1_18_pdst,
              rob_uop_1_17_pdst,
              rob_uop_1_16_pdst,
              rob_uop_1_15_pdst,
              rob_uop_1_14_pdst,
              rob_uop_1_13_pdst,
              rob_uop_1_12_pdst,
              rob_uop_1_11_pdst,
              rob_uop_1_10_pdst,
              rob_uop_1_9_pdst,
              rob_uop_1_8_pdst,
              rob_uop_1_7_pdst,
              rob_uop_1_6_pdst,
              rob_uop_1_5_pdst,
              rob_uop_1_4_pdst,
              rob_uop_1_3_pdst,
              rob_uop_1_2_pdst,
              rob_uop_1_1_pdst,
              rob_uop_1_0_pdst,
  input       rob_uop_1_31_ldst_val,
              rob_uop_1_30_ldst_val,
              rob_uop_1_29_ldst_val,
              rob_uop_1_28_ldst_val,
              rob_uop_1_27_ldst_val,
              rob_uop_1_26_ldst_val,
              rob_uop_1_25_ldst_val,
              rob_uop_1_24_ldst_val,
              rob_uop_1_23_ldst_val,
              rob_uop_1_22_ldst_val,
              rob_uop_1_21_ldst_val,
              rob_uop_1_20_ldst_val,
              rob_uop_1_19_ldst_val,
              rob_uop_1_18_ldst_val,
              rob_uop_1_17_ldst_val,
              rob_uop_1_16_ldst_val,
              rob_uop_1_15_ldst_val,
              rob_uop_1_14_ldst_val,
              rob_uop_1_13_ldst_val,
              rob_uop_1_12_ldst_val,
              rob_uop_1_11_ldst_val,
              rob_uop_1_10_ldst_val,
              rob_uop_1_9_ldst_val,
              rob_uop_1_8_ldst_val,
              rob_uop_1_7_ldst_val,
              rob_uop_1_6_ldst_val,
              rob_uop_1_5_ldst_val,
              rob_uop_1_4_ldst_val,
              rob_uop_1_3_ldst_val,
              rob_uop_1_2_ldst_val,
              rob_uop_1_1_ldst_val,
              rob_uop_1_0_ldst_val,
              _GEN_917,
              _GEN_918,
              _GEN_919,
              _GEN_920,
              rob_val_2_31,
              rob_val_2_30,
              rob_val_2_29,
              rob_val_2_28,
              rob_val_2_27,
              rob_val_2_26,
              rob_val_2_25,
              rob_val_2_24,
              rob_val_2_23,
              rob_val_2_22,
              rob_val_2_21,
              rob_val_2_20,
              rob_val_2_19,
              rob_val_2_18,
              rob_val_2_17,
              rob_val_2_16,
              rob_val_2_15,
              rob_val_2_14,
              rob_val_2_13,
              rob_val_2_12,
              rob_val_2_11,
              rob_val_2_10,
              rob_val_2_9,
              rob_val_2_8,
              rob_val_2_7,
              rob_val_2_6,
              rob_val_2_5,
              rob_val_2_4,
              rob_val_2_3,
              rob_val_2_2,
              rob_val_2_1,
              rob_val_2_0,
  input [6:0] io_enq_uops_2_rob_idx,
  input       rob_bsy_2_31,
              rob_bsy_2_30,
              rob_bsy_2_29,
              rob_bsy_2_28,
              rob_bsy_2_27,
              rob_bsy_2_26,
              rob_bsy_2_25,
              rob_bsy_2_24,
              rob_bsy_2_23,
              rob_bsy_2_22,
              rob_bsy_2_21,
              rob_bsy_2_20,
              rob_bsy_2_19,
              rob_bsy_2_18,
              rob_bsy_2_17,
              rob_bsy_2_16,
              rob_bsy_2_15,
              rob_bsy_2_14,
              rob_bsy_2_13,
              rob_bsy_2_12,
              rob_bsy_2_11,
              rob_bsy_2_10,
              rob_bsy_2_9,
              rob_bsy_2_8,
              rob_bsy_2_7,
              rob_bsy_2_6,
              rob_bsy_2_5,
              rob_bsy_2_4,
              rob_bsy_2_3,
              rob_bsy_2_2,
              rob_bsy_2_1,
              rob_bsy_2_0,
              _GEN_921,
              _GEN_922,
              _GEN_923,
              _GEN_924,
              _GEN_925,
              _GEN_926,
              _GEN_927,
              io_enq_uops_2_uses_ldq,
              io_enq_uops_2_is_br,
              io_enq_uops_2_is_jalr,
              io_enq_uops_2_uses_stq,
              io_enq_uops_2_is_fence,
              _GEN_928,
              _GEN_929,
              _GEN_930,
              _GEN_931,
              _GEN_932,
              _GEN_933,
              _GEN_934,
              _GEN_935,
              _GEN_936,
              _GEN_937,
              _GEN_938,
              _GEN_939,
              _GEN_940,
              _GEN_941,
              _GEN_942,
              _GEN_943,
              _GEN_944,
              _GEN_945,
              _GEN_946,
              _GEN_947,
              _GEN_948,
              _GEN_949,
              _GEN_950,
              _GEN_951,
              _GEN_952,
              _GEN_953,
              _GEN_954,
              _GEN_955,
              _GEN_956,
              _GEN_957,
              _GEN_958,
              _GEN_959,
              _GEN_960,
              _GEN_961,
              _GEN_962,
              _GEN_963,
              _GEN_964,
              _GEN_965,
              _GEN_966,
              _GEN_967,
              _GEN_968,
              _GEN_969,
              _GEN_970,
              _GEN_971,
              _GEN_972,
              _GEN_973,
              _GEN_974,
              _GEN_975,
              _GEN_976,
              _GEN_977,
              _GEN_978,
              _GEN_979,
              _GEN_980,
              _GEN_981,
              _GEN_982,
              _GEN_983,
              _GEN_984,
              _GEN_985,
              _GEN_986,
              _GEN_987,
              _GEN_988,
              _GEN_989,
              _GEN_990,
              _GEN_991,
              _GEN_992,
              _GEN_993,
              _GEN_994,
              _GEN_995,
              _GEN_996,
              _GEN_997,
              _GEN_998,
              _GEN_999,
              _GEN_1000,
              _GEN_1001,
              _GEN_1002,
              _GEN_1003,
              _GEN_1004,
              _GEN_1005,
              _GEN_1006,
              _GEN_1007,
              _GEN_1008,
              _GEN_1009,
              _GEN_1010,
              _GEN_1011,
              _GEN_1012,
              _GEN_1013,
              _GEN_1014,
              _GEN_1015,
              _GEN_1016,
              _GEN_1017,
              _GEN_1018,
              _GEN_1019,
              _GEN_1020,
              _GEN_1021,
              _GEN_1022,
              _GEN_1023,
              _GEN_1024,
              _GEN_1025,
              _GEN_1026,
              _GEN_1027,
              _GEN_1028,
              _GEN_1029,
              _GEN_1030,
              _GEN_1031,
              _GEN_1032,
              _GEN_1033,
              _GEN_1034,
              _GEN_1035,
              _GEN_1036,
              _GEN_1037,
              _GEN_1038,
              _GEN_1039,
              _GEN_1040,
              _GEN_1041,
              _GEN_1042,
              _GEN_1043,
              _GEN_1044,
              _GEN_1045,
              _GEN_1046,
              _GEN_1047,
              _GEN_1048,
              _GEN_1049,
              _GEN_1050,
              _GEN_1051,
              _GEN_1052,
              _GEN_1053,
              _GEN_1054,
              _GEN_1055,
              _GEN_1056,
              _GEN_1057,
              _GEN_1058,
              _GEN_1059,
              _GEN_1060,
              _GEN_1061,
              _GEN_1062,
              _GEN_1063,
              _GEN_1064,
              _GEN_1065,
              _GEN_1066,
              _GEN_1067,
              _GEN_1068,
              _GEN_1069,
              _GEN_1070,
              _GEN_1071,
              _GEN_1072,
              _GEN_1073,
              _GEN_1074,
              _GEN_1075,
              _GEN_1076,
              _GEN_1077,
              _GEN_1078,
              _GEN_1079,
              _GEN_1080,
              _GEN_1081,
              _GEN_1082,
              _GEN_1083,
              _GEN_1084,
              _GEN_1085,
              _GEN_1086,
              _GEN_1087,
              _GEN_1088,
              _GEN_1089,
              _GEN_1090,
              _GEN_1091,
              _GEN_1092,
              _GEN_1093,
              _GEN_1094,
              _GEN_1095,
              _GEN_1096,
              _GEN_1097,
              _GEN_1098,
              _GEN_1099,
              _GEN_1100,
              _GEN_1101,
              _GEN_1102,
              _GEN_1103,
              _GEN_1104,
              _GEN_1105,
              _GEN_1106,
              _GEN_1107,
              _GEN_1108,
              _GEN_1109,
              _GEN_1110,
              _GEN_1111,
              _GEN_1112,
              _GEN_1113,
              _GEN_1114,
              _GEN_1115,
              _GEN_1116,
              _GEN_1117,
              _GEN_1118,
              _GEN_1119,
              _GEN_1120,
              _GEN_1121,
              _GEN_1122,
              _GEN_1123,
              _GEN_1124,
              _GEN_1125,
              _GEN_1126,
              _GEN_1127,
              _GEN_1128,
              _GEN_1129,
              _GEN_1130,
              _GEN_1131,
              _GEN_1132,
              _GEN_1133,
              _GEN_1134,
              _GEN_1135,
              _GEN_1136,
              _GEN_1137,
              _GEN_1138,
              _GEN_1139,
              _GEN_1140,
              _GEN_1141,
              _GEN_1142,
              _GEN_1143,
              _GEN_1144,
              _GEN_1145,
              _GEN_1146,
              _GEN_1147,
              _GEN_1148,
              _GEN_1149,
              _GEN_1150,
              _GEN_1151,
              _GEN_1152,
              _GEN_1153,
              _GEN_1154,
              _GEN_1155,
              _GEN_1156,
              _GEN_1157,
              _GEN_1158,
              _GEN_1159,
              _GEN_1160,
              _GEN_1161,
              _GEN_1162,
              _GEN_1163,
              _GEN_1164,
              _GEN_1165,
              _GEN_1166,
              _GEN_1167,
              _GEN_1168,
              _GEN_1169,
              _GEN_1170,
              _GEN_1171,
              _GEN_1172,
              _GEN_1173,
              _GEN_1174,
              _GEN_1175,
              _GEN_1176,
              _GEN_1177,
              _GEN_1178,
              _GEN_1179,
              _GEN_1180,
              _GEN_1181,
              _GEN_1182,
              _GEN_1183,
              _GEN_1184,
              _GEN_1185,
              _GEN_1186,
              _GEN_1187,
              _GEN_1188,
              _GEN_1189,
              _GEN_1190,
              _GEN_1191,
              _GEN_1192,
              _GEN_1193,
              _GEN_1194,
              _GEN_1195,
              _GEN_1196,
              _GEN_1197,
              _GEN_1198,
              _GEN_1199,
              _GEN_1200,
              _GEN_1201,
              _GEN_1202,
              _GEN_1203,
              _GEN_1204,
              _GEN_1205,
              _GEN_1206,
              _GEN_1207,
              _GEN_1208,
              _GEN_1209,
              _GEN_1210,
              _GEN_1211,
              _GEN_1212,
              _GEN_1213,
              _GEN_1214,
              _GEN_1215,
              _GEN_1216,
              _GEN_1217,
              _GEN_1218,
              _GEN_1219,
              _GEN_1220,
              _GEN_1221,
              _GEN_1222,
              _GEN_1223,
              _GEN_1224,
              _GEN_1225,
              _GEN_1226,
              _GEN_1227,
              _GEN_1228,
              _GEN_1229,
              _GEN_1230,
              _GEN_1231,
              _GEN_1232,
              _GEN_1233,
              _GEN_1234,
              _GEN_1235,
              _GEN_1236,
              _GEN_1237,
              _GEN_1238,
              _GEN_1239,
              _GEN_1240,
              _GEN_1241,
              _GEN_1242,
              _GEN_1243,
              _GEN_1244,
              _GEN_1245,
              _GEN_1246,
              _GEN_1247,
              _GEN_1248,
              _GEN_1249,
              _GEN_1250,
              _GEN_1251,
              _GEN_1252,
              _GEN_1253,
              _GEN_1254,
              _GEN_1255,
              _GEN_1256,
              _GEN_1257,
              _GEN_1258,
              _GEN_1259,
              _GEN_1260,
              _GEN_1261,
              _GEN_1262,
              _GEN_1263,
              _GEN_1264,
              _GEN_1265,
              _GEN_1266,
              _GEN_1267,
              _GEN_1268,
              _GEN_1269,
              _GEN_1270,
              _GEN_1271,
              _GEN_1272,
              _GEN_1273,
              _GEN_1274,
              _GEN_1275,
              _GEN_1276,
              _GEN_1277,
              _GEN_1278,
              _GEN_1279,
              _GEN_1280,
              _GEN_1281,
              _GEN_1282,
              _GEN_1283,
              _GEN_1284,
              _GEN_1285,
              _GEN_1286,
              _GEN_1287,
              _GEN_1288,
              _GEN_1289,
              _GEN_1290,
              _GEN_1291,
              _GEN_1292,
              _GEN_1293,
              _GEN_1294,
              _GEN_1295,
              _GEN_1296,
              _GEN_1297,
              _GEN_1298,
              _GEN_1299,
              _GEN_1300,
              _GEN_1301,
              _GEN_1302,
              _GEN_1303,
              _GEN_1304,
              _GEN_1305,
              _GEN_1306,
              _GEN_1307,
              _GEN_1308,
              _GEN_1309,
              _GEN_1310,
              _GEN_1311,
              _GEN_1312,
              _GEN_1313,
              _GEN_1314,
              _GEN_1315,
              _GEN_1316,
              _GEN_1317,
              _GEN_1318,
              _GEN_1319,
              _GEN_1320,
              _GEN_1321,
              _GEN_1322,
              _GEN_1323,
              _GEN_1324,
              _GEN_1325,
              _GEN_1326,
              _GEN_1327,
              _GEN_1328,
              _GEN_1329,
              _GEN_1330,
              _GEN_1331,
              _GEN_1332,
              _GEN_1333,
              _GEN_1334,
              _GEN_1335,
              _GEN_1336,
              _GEN_1337,
              _GEN_1338,
              _GEN_1339,
              _GEN_1340,
              _GEN_1341,
              _GEN_1342,
              _GEN_1343,
              _GEN_1344,
              _GEN_1345,
              _GEN_1346,
              _GEN_1347,
              _GEN_1348,
              _GEN_1349,
              _GEN_1350,
              _GEN_1351,
              _GEN_1352,
              _GEN_1353,
              _GEN_1354,
              _GEN_1355,
              _GEN_1356,
              _GEN_1357,
              _GEN_1358,
              _GEN_1359,
              _GEN_1360,
              _GEN_1361,
              _GEN_1362,
              _GEN_1363,
              _GEN_1364,
              _GEN_1365,
              _GEN_1366,
              _GEN_1367,
              _GEN_1368,
              _GEN_1369,
              _GEN_1370,
              _GEN_1371,
              _GEN_1372,
              _GEN_1373,
              _GEN_1374,
              _GEN_1375,
  input [6:0] rob_uop_2_31_pdst,
              rob_uop_2_30_pdst,
              rob_uop_2_29_pdst,
              rob_uop_2_28_pdst,
              rob_uop_2_27_pdst,
              rob_uop_2_26_pdst,
              rob_uop_2_25_pdst,
              rob_uop_2_24_pdst,
              rob_uop_2_23_pdst,
              rob_uop_2_22_pdst,
              rob_uop_2_21_pdst,
              rob_uop_2_20_pdst,
              rob_uop_2_19_pdst,
              rob_uop_2_18_pdst,
              rob_uop_2_17_pdst,
              rob_uop_2_16_pdst,
              rob_uop_2_15_pdst,
              rob_uop_2_14_pdst,
              rob_uop_2_13_pdst,
              rob_uop_2_12_pdst,
              rob_uop_2_11_pdst,
              rob_uop_2_10_pdst,
              rob_uop_2_9_pdst,
              rob_uop_2_8_pdst,
              rob_uop_2_7_pdst,
              rob_uop_2_6_pdst,
              rob_uop_2_5_pdst,
              rob_uop_2_4_pdst,
              rob_uop_2_3_pdst,
              rob_uop_2_2_pdst,
              rob_uop_2_1_pdst,
              rob_uop_2_0_pdst,
  input       rob_uop_2_31_ldst_val,
              rob_uop_2_30_ldst_val,
              rob_uop_2_29_ldst_val,
              rob_uop_2_28_ldst_val,
              rob_uop_2_27_ldst_val,
              rob_uop_2_26_ldst_val,
              rob_uop_2_25_ldst_val,
              rob_uop_2_24_ldst_val,
              rob_uop_2_23_ldst_val,
              rob_uop_2_22_ldst_val,
              rob_uop_2_21_ldst_val,
              rob_uop_2_20_ldst_val,
              rob_uop_2_19_ldst_val,
              rob_uop_2_18_ldst_val,
              rob_uop_2_17_ldst_val,
              rob_uop_2_16_ldst_val,
              rob_uop_2_15_ldst_val,
              rob_uop_2_14_ldst_val,
              rob_uop_2_13_ldst_val,
              rob_uop_2_12_ldst_val,
              rob_uop_2_11_ldst_val,
              rob_uop_2_10_ldst_val,
              rob_uop_2_9_ldst_val,
              rob_uop_2_8_ldst_val,
              rob_uop_2_7_ldst_val,
              rob_uop_2_6_ldst_val,
              rob_uop_2_5_ldst_val,
              rob_uop_2_4_ldst_val,
              rob_uop_2_3_ldst_val,
              rob_uop_2_2_ldst_val,
              rob_uop_2_1_ldst_val,
              rob_uop_2_0_ldst_val,
              _GEN_1376,
              _GEN_1377,
              _GEN_1378,
              _GEN_1379,
              rob_val_3_31,
              rob_val_3_30,
              rob_val_3_29,
              rob_val_3_28,
              rob_val_3_27,
              rob_val_3_26,
              rob_val_3_25,
              rob_val_3_24,
              rob_val_3_23,
              rob_val_3_22,
              rob_val_3_21,
              rob_val_3_20,
              rob_val_3_19,
              rob_val_3_18,
              rob_val_3_17,
              rob_val_3_16,
              rob_val_3_15,
              rob_val_3_14,
              rob_val_3_13,
              rob_val_3_12,
              rob_val_3_11,
              rob_val_3_10,
              rob_val_3_9,
              rob_val_3_8,
              rob_val_3_7,
              rob_val_3_6,
              rob_val_3_5,
              rob_val_3_4,
              rob_val_3_3,
              rob_val_3_2,
              rob_val_3_1,
              rob_val_3_0,
  input [6:0] io_enq_uops_3_rob_idx,
  input       rob_bsy_3_31,
              rob_bsy_3_30,
              rob_bsy_3_29,
              rob_bsy_3_28,
              rob_bsy_3_27,
              rob_bsy_3_26,
              rob_bsy_3_25,
              rob_bsy_3_24,
              rob_bsy_3_23,
              rob_bsy_3_22,
              rob_bsy_3_21,
              rob_bsy_3_20,
              rob_bsy_3_19,
              rob_bsy_3_18,
              rob_bsy_3_17,
              rob_bsy_3_16,
              rob_bsy_3_15,
              rob_bsy_3_14,
              rob_bsy_3_13,
              rob_bsy_3_12,
              rob_bsy_3_11,
              rob_bsy_3_10,
              rob_bsy_3_9,
              rob_bsy_3_8,
              rob_bsy_3_7,
              rob_bsy_3_6,
              rob_bsy_3_5,
              rob_bsy_3_4,
              rob_bsy_3_3,
              rob_bsy_3_2,
              rob_bsy_3_1,
              rob_bsy_3_0,
              _GEN_1380,
              _GEN_1381,
              _GEN_1382,
              _GEN_1383,
              _GEN_1384,
              _GEN_1385,
              _GEN_1386,
              io_enq_uops_3_uses_ldq,
              io_enq_uops_3_is_br,
              io_enq_uops_3_is_jalr,
              io_enq_uops_3_uses_stq,
              io_enq_uops_3_is_fence,
              _GEN_1387,
              _GEN_1388,
              _GEN_1389,
              _GEN_1390,
              _GEN_1391,
              _GEN_1392,
              _GEN_1393,
              _GEN_1394,
              _GEN_1395,
              _GEN_1396,
              _GEN_1397,
              _GEN_1398,
              _GEN_1399,
              _GEN_1400,
              _GEN_1401,
              _GEN_1402,
              _GEN_1403,
              _GEN_1404,
              _GEN_1405,
              _GEN_1406,
              _GEN_1407,
              _GEN_1408,
              _GEN_1409,
              _GEN_1410,
              _GEN_1411,
              _GEN_1412,
              _GEN_1413,
              _GEN_1414,
              _GEN_1415,
              _GEN_1416,
              _GEN_1417,
              _GEN_1418,
              _GEN_1419,
              _GEN_1420,
              _GEN_1421,
              _GEN_1422,
              _GEN_1423,
              _GEN_1424,
              _GEN_1425,
              _GEN_1426,
              _GEN_1427,
              _GEN_1428,
              _GEN_1429,
              _GEN_1430,
              _GEN_1431,
              _GEN_1432,
              _GEN_1433,
              _GEN_1434,
              _GEN_1435,
              _GEN_1436,
              _GEN_1437,
              _GEN_1438,
              _GEN_1439,
              _GEN_1440,
              _GEN_1441,
              _GEN_1442,
              _GEN_1443,
              _GEN_1444,
              _GEN_1445,
              _GEN_1446,
              _GEN_1447,
              _GEN_1448,
              _GEN_1449,
              _GEN_1450,
              _GEN_1451,
              _GEN_1452,
              _GEN_1453,
              _GEN_1454,
              _GEN_1455,
              _GEN_1456,
              _GEN_1457,
              _GEN_1458,
              _GEN_1459,
              _GEN_1460,
              _GEN_1461,
              _GEN_1462,
              _GEN_1463,
              _GEN_1464,
              _GEN_1465,
              _GEN_1466,
              _GEN_1467,
              _GEN_1468,
              _GEN_1469,
              _GEN_1470,
              _GEN_1471,
              _GEN_1472,
              _GEN_1473,
              _GEN_1474,
              _GEN_1475,
              _GEN_1476,
              _GEN_1477,
              _GEN_1478,
              _GEN_1479,
              _GEN_1480,
              _GEN_1481,
              _GEN_1482,
              _GEN_1483,
              _GEN_1484,
              _GEN_1485,
              _GEN_1486,
              _GEN_1487,
              _GEN_1488,
              _GEN_1489,
              _GEN_1490,
              _GEN_1491,
              _GEN_1492,
              _GEN_1493,
              _GEN_1494,
              _GEN_1495,
              _GEN_1496,
              _GEN_1497,
              _GEN_1498,
              _GEN_1499,
              _GEN_1500,
              _GEN_1501,
              _GEN_1502,
              _GEN_1503,
              _GEN_1504,
              _GEN_1505,
              _GEN_1506,
              _GEN_1507,
              _GEN_1508,
              _GEN_1509,
              _GEN_1510,
              _GEN_1511,
              _GEN_1512,
              _GEN_1513,
              _GEN_1514,
              _GEN_1515,
              _GEN_1516,
              _GEN_1517,
              _GEN_1518,
              _GEN_1519,
              _GEN_1520,
              _GEN_1521,
              _GEN_1522,
              _GEN_1523,
              _GEN_1524,
              _GEN_1525,
              _GEN_1526,
              _GEN_1527,
              _GEN_1528,
              _GEN_1529,
              _GEN_1530,
              _GEN_1531,
              _GEN_1532,
              _GEN_1533,
              _GEN_1534,
              _GEN_1535,
              _GEN_1536,
              _GEN_1537,
              _GEN_1538,
              _GEN_1539,
              _GEN_1540,
              _GEN_1541,
              _GEN_1542,
              _GEN_1543,
              _GEN_1544,
              _GEN_1545,
              _GEN_1546,
              _GEN_1547,
              _GEN_1548,
              _GEN_1549,
              _GEN_1550,
              _GEN_1551,
              _GEN_1552,
              _GEN_1553,
              _GEN_1554,
              _GEN_1555,
              _GEN_1556,
              _GEN_1557,
              _GEN_1558,
              _GEN_1559,
              _GEN_1560,
              _GEN_1561,
              _GEN_1562,
              _GEN_1563,
              _GEN_1564,
              _GEN_1565,
              _GEN_1566,
              _GEN_1567,
              _GEN_1568,
              _GEN_1569,
              _GEN_1570,
              _GEN_1571,
              _GEN_1572,
              _GEN_1573,
              _GEN_1574,
              _GEN_1575,
              _GEN_1576,
              _GEN_1577,
              _GEN_1578,
              _GEN_1579,
              _GEN_1580,
              _GEN_1581,
              _GEN_1582,
              _GEN_1583,
              _GEN_1584,
              _GEN_1585,
              _GEN_1586,
              _GEN_1587,
              _GEN_1588,
              _GEN_1589,
              _GEN_1590,
              _GEN_1591,
              _GEN_1592,
              _GEN_1593,
              _GEN_1594,
              _GEN_1595,
              _GEN_1596,
              _GEN_1597,
              _GEN_1598,
              _GEN_1599,
              _GEN_1600,
              _GEN_1601,
              _GEN_1602,
              _GEN_1603,
              _GEN_1604,
              _GEN_1605,
              _GEN_1606,
              _GEN_1607,
              _GEN_1608,
              _GEN_1609,
              _GEN_1610,
              _GEN_1611,
              _GEN_1612,
              _GEN_1613,
              _GEN_1614,
              _GEN_1615,
              _GEN_1616,
              _GEN_1617,
              _GEN_1618,
              _GEN_1619,
              _GEN_1620,
              _GEN_1621,
              _GEN_1622,
              _GEN_1623,
              _GEN_1624,
              _GEN_1625,
              _GEN_1626,
              _GEN_1627,
              _GEN_1628,
              _GEN_1629,
              _GEN_1630,
              _GEN_1631,
              _GEN_1632,
              _GEN_1633,
              _GEN_1634,
              _GEN_1635,
              _GEN_1636,
              _GEN_1637,
              _GEN_1638,
              _GEN_1639,
              _GEN_1640,
              _GEN_1641,
              _GEN_1642,
              _GEN_1643,
              _GEN_1644,
              _GEN_1645,
              _GEN_1646,
              _GEN_1647,
              _GEN_1648,
              _GEN_1649,
              _GEN_1650,
              _GEN_1651,
              _GEN_1652,
              _GEN_1653,
              _GEN_1654,
              _GEN_1655,
              _GEN_1656,
              _GEN_1657,
              _GEN_1658,
              _GEN_1659,
              _GEN_1660,
              _GEN_1661,
              _GEN_1662,
              _GEN_1663,
              _GEN_1664,
              _GEN_1665,
              _GEN_1666,
              _GEN_1667,
              _GEN_1668,
              _GEN_1669,
              _GEN_1670,
              _GEN_1671,
              _GEN_1672,
              _GEN_1673,
              _GEN_1674,
              _GEN_1675,
              _GEN_1676,
              _GEN_1677,
              _GEN_1678,
              _GEN_1679,
              _GEN_1680,
              _GEN_1681,
              _GEN_1682,
              _GEN_1683,
              _GEN_1684,
              _GEN_1685,
              _GEN_1686,
              _GEN_1687,
              _GEN_1688,
              _GEN_1689,
              _GEN_1690,
              _GEN_1691,
              _GEN_1692,
              _GEN_1693,
              _GEN_1694,
              _GEN_1695,
              _GEN_1696,
              _GEN_1697,
              _GEN_1698,
              _GEN_1699,
              _GEN_1700,
              _GEN_1701,
              _GEN_1702,
              _GEN_1703,
              _GEN_1704,
              _GEN_1705,
              _GEN_1706,
              _GEN_1707,
              _GEN_1708,
              _GEN_1709,
              _GEN_1710,
              _GEN_1711,
              _GEN_1712,
              _GEN_1713,
              _GEN_1714,
              _GEN_1715,
              _GEN_1716,
              _GEN_1717,
              _GEN_1718,
              _GEN_1719,
              _GEN_1720,
              _GEN_1721,
              _GEN_1722,
              _GEN_1723,
              _GEN_1724,
              _GEN_1725,
              _GEN_1726,
              _GEN_1727,
              _GEN_1728,
              _GEN_1729,
              _GEN_1730,
              _GEN_1731,
              _GEN_1732,
              _GEN_1733,
              _GEN_1734,
              _GEN_1735,
              _GEN_1736,
              _GEN_1737,
              _GEN_1738,
              _GEN_1739,
              _GEN_1740,
              _GEN_1741,
              _GEN_1742,
              _GEN_1743,
              _GEN_1744,
              _GEN_1745,
              _GEN_1746,
              _GEN_1747,
              _GEN_1748,
              _GEN_1749,
              _GEN_1750,
              _GEN_1751,
              _GEN_1752,
              _GEN_1753,
              _GEN_1754,
              _GEN_1755,
              _GEN_1756,
              _GEN_1757,
              _GEN_1758,
              _GEN_1759,
              _GEN_1760,
              _GEN_1761,
              _GEN_1762,
              _GEN_1763,
              _GEN_1764,
              _GEN_1765,
              _GEN_1766,
              _GEN_1767,
              _GEN_1768,
              _GEN_1769,
              _GEN_1770,
              _GEN_1771,
              _GEN_1772,
              _GEN_1773,
              _GEN_1774,
              _GEN_1775,
              _GEN_1776,
              _GEN_1777,
              _GEN_1778,
              _GEN_1779,
              _GEN_1780,
              _GEN_1781,
              _GEN_1782,
              _GEN_1783,
              _GEN_1784,
              _GEN_1785,
              _GEN_1786,
              _GEN_1787,
              _GEN_1788,
              _GEN_1789,
              _GEN_1790,
              _GEN_1791,
              _GEN_1792,
              _GEN_1793,
              _GEN_1794,
              _GEN_1795,
              _GEN_1796,
              _GEN_1797,
              _GEN_1798,
              _GEN_1799,
              _GEN_1800,
              _GEN_1801,
              _GEN_1802,
              _GEN_1803,
              _GEN_1804,
              _GEN_1805,
              _GEN_1806,
              _GEN_1807,
              _GEN_1808,
              _GEN_1809,
              _GEN_1810,
              _GEN_1811,
              _GEN_1812,
              _GEN_1813,
              _GEN_1814,
              _GEN_1815,
              _GEN_1816,
              _GEN_1817,
              _GEN_1818,
              _GEN_1819,
              _GEN_1820,
              _GEN_1821,
              _GEN_1822,
              _GEN_1823,
              _GEN_1824,
              _GEN_1825,
              _GEN_1826,
              _GEN_1827,
              _GEN_1828,
              _GEN_1829,
              _GEN_1830,
              _GEN_1831,
              _GEN_1832,
              _GEN_1833,
              _GEN_1834,
  input [6:0] rob_uop_3_31_pdst,
              rob_uop_3_30_pdst,
              rob_uop_3_29_pdst,
              rob_uop_3_28_pdst,
              rob_uop_3_27_pdst,
              rob_uop_3_26_pdst,
              rob_uop_3_25_pdst,
              rob_uop_3_24_pdst,
              rob_uop_3_23_pdst,
              rob_uop_3_22_pdst,
              rob_uop_3_21_pdst,
              rob_uop_3_20_pdst,
              rob_uop_3_19_pdst,
              rob_uop_3_18_pdst,
              rob_uop_3_17_pdst,
              rob_uop_3_16_pdst,
              rob_uop_3_15_pdst,
              rob_uop_3_14_pdst,
              rob_uop_3_13_pdst,
              rob_uop_3_12_pdst,
              rob_uop_3_11_pdst,
              rob_uop_3_10_pdst,
              rob_uop_3_9_pdst,
              rob_uop_3_8_pdst,
              rob_uop_3_7_pdst,
              rob_uop_3_6_pdst,
              rob_uop_3_5_pdst,
              rob_uop_3_4_pdst,
              rob_uop_3_3_pdst,
              rob_uop_3_2_pdst,
              rob_uop_3_1_pdst,
              rob_uop_3_0_pdst,
  input       rob_uop_3_31_ldst_val,
              rob_uop_3_30_ldst_val,
              rob_uop_3_29_ldst_val,
              rob_uop_3_28_ldst_val,
              rob_uop_3_27_ldst_val,
              rob_uop_3_26_ldst_val,
              rob_uop_3_25_ldst_val,
              rob_uop_3_24_ldst_val,
              rob_uop_3_23_ldst_val,
              rob_uop_3_22_ldst_val,
              rob_uop_3_21_ldst_val,
              rob_uop_3_20_ldst_val,
              rob_uop_3_19_ldst_val,
              rob_uop_3_18_ldst_val,
              rob_uop_3_17_ldst_val,
              rob_uop_3_16_ldst_val,
              rob_uop_3_15_ldst_val,
              rob_uop_3_14_ldst_val,
              rob_uop_3_13_ldst_val,
              rob_uop_3_12_ldst_val,
              rob_uop_3_11_ldst_val,
              rob_uop_3_10_ldst_val,
              rob_uop_3_9_ldst_val,
              rob_uop_3_8_ldst_val,
              rob_uop_3_7_ldst_val,
              rob_uop_3_6_ldst_val,
              rob_uop_3_5_ldst_val,
              rob_uop_3_4_ldst_val,
              rob_uop_3_3_ldst_val,
              rob_uop_3_2_ldst_val,
              rob_uop_3_1_ldst_val,
              rob_uop_3_0_ldst_val,
              _GEN_1835,
              _GEN_1836,
              _GEN_1837,
              _GEN_1838,
              flush_commit_mask_3,
              flush_commit_mask_2,
              flush_commit_mask_1,
              flush_commit_mask_0,
  input [4:0] rob_head_fflags_0,
  input       _rob_uop_com_idx_fp_val,
              _fflags_val_0_T,
              _io_commit_uops_0_uses_ldq_output,
              _io_commit_uops_0_uses_stq_output,
  input [4:0] rob_head_fflags_1,
  input       _rob_uop_1_com_idx_fp_val,
              _fflags_val_1_T,
              _io_commit_uops_1_uses_ldq_output,
              _io_commit_uops_1_uses_stq_output,
  input [4:0] rob_head_fflags_2,
  input       _rob_uop_2_com_idx_fp_val,
              _fflags_val_2_T,
              _io_commit_uops_2_uses_ldq_output,
              _io_commit_uops_2_uses_stq_output,
  input [4:0] rob_head_fflags_3,
  input       _rob_uop_3_com_idx_fp_val,
              _fflags_val_3_T,
              _io_commit_uops_3_uses_ldq_output,
              _io_commit_uops_3_uses_stq_output,
              exception_thrown,
              _io_ready_T_3,
              empty,
              r_xcpt_val,
  input [4:0] rob_head,
  input [6:0] r_xcpt_uop_rob_idx,
              rob_tail_idx,
  input       reset,
              full,
              _maybe_full_T,
              _io_ready_T,
  input [1:0] rob_state,
  input       _GEN_1839,
              rob_exception_3_31,
              rob_exception_3_30,
              rob_exception_3_29,
              rob_exception_3_28,
              rob_exception_3_27,
              rob_exception_3_26,
              rob_exception_3_25,
              rob_exception_3_24,
              rob_exception_3_23,
              rob_exception_3_22,
              rob_exception_3_21,
              rob_exception_3_20,
              rob_exception_3_19,
              rob_exception_3_18,
              rob_exception_3_17,
              rob_exception_3_16,
              rob_exception_3_15,
              rob_exception_3_14,
              rob_exception_3_13,
              rob_exception_3_12,
              rob_exception_3_11,
              rob_exception_3_10,
              rob_exception_3_9,
              rob_exception_3_8,
              rob_exception_3_7,
              rob_exception_3_6,
              rob_exception_3_5,
              rob_exception_3_4,
              rob_exception_3_3,
              rob_exception_3_2,
              rob_exception_3_1,
              rob_exception_3_0,
              rob_exception_2_31,
              rob_exception_2_30,
              rob_exception_2_29,
              rob_exception_2_28,
              rob_exception_2_27,
              rob_exception_2_26,
              rob_exception_2_25,
              rob_exception_2_24,
              rob_exception_2_23,
              rob_exception_2_22,
              rob_exception_2_21,
              rob_exception_2_20,
              rob_exception_2_19,
              rob_exception_2_18,
              rob_exception_2_17,
              rob_exception_2_16,
              rob_exception_2_15,
              rob_exception_2_14,
              rob_exception_2_13,
              rob_exception_2_12,
              rob_exception_2_11,
              rob_exception_2_10,
              rob_exception_2_9,
              rob_exception_2_8,
              rob_exception_2_7,
              rob_exception_2_6,
              rob_exception_2_5,
              rob_exception_2_4,
              rob_exception_2_3,
              rob_exception_2_2,
              rob_exception_2_1,
              rob_exception_2_0,
              rob_exception_1_31,
              rob_exception_1_30,
              rob_exception_1_29,
              rob_exception_1_28,
              rob_exception_1_27,
              rob_exception_1_26,
              rob_exception_1_25,
              rob_exception_1_24,
              rob_exception_1_23,
              rob_exception_1_22,
              rob_exception_1_21,
              rob_exception_1_20,
              rob_exception_1_19,
              rob_exception_1_18,
              rob_exception_1_17,
              rob_exception_1_16,
              rob_exception_1_15,
              rob_exception_1_14,
              rob_exception_1_13,
              rob_exception_1_12,
              rob_exception_1_11,
              rob_exception_1_10,
              rob_exception_1_9,
              rob_exception_1_8,
              rob_exception_1_7,
              rob_exception_1_6,
              rob_exception_1_5,
              rob_exception_1_4,
              rob_exception_1_3,
              rob_exception_1_2,
              rob_exception_1_1,
              rob_exception_1_0,
              rob_exception__31,
              rob_exception__30,
              rob_exception__29,
              rob_exception__28,
              rob_exception__27,
              rob_exception__26,
              rob_exception__25,
              rob_exception__24,
              rob_exception__23,
              rob_exception__22,
              rob_exception__21,
              rob_exception__20,
              rob_exception__19,
              rob_exception__18,
              rob_exception__17,
              rob_exception__16,
              rob_exception__15,
              rob_exception__14,
              rob_exception__13,
              rob_exception__12,
              rob_exception__11,
              rob_exception__10,
              rob_exception__9,
              rob_exception__8,
              rob_exception__7,
              rob_exception__6,
              rob_exception__5,
              rob_exception__4,
              rob_exception__3,
              rob_exception__2,
              rob_exception__1,
              rob_exception__0,
              _io_ready_T_1,
              io_enq_valids_0,
              io_enq_valids_1,
              io_enq_valids_2,
  input [6:0] rob_head_idx,
  input       _GEN_1840,
              _GEN_1841,
              _GEN_1842,
  input [4:0] io_lxcpt_bits_cause,
  input       _GEN_1843,
              _GEN_1844,
              _GEN_1845,
              _GEN_1846,
              _GEN_1847,
              _GEN_1848,
              io_enq_valids_3,
              _GEN_1849,
              _GEN_1850,
              _GEN_1851
);

  reg        casez_tmp;
  reg        casez_tmp_0;
  reg        casez_tmp_1;
  reg        casez_tmp_2;
  reg        casez_tmp_3;
  reg        casez_tmp_4;
  reg        casez_tmp_5;
  reg        casez_tmp_6;
  reg        casez_tmp_7;
  reg        casez_tmp_8;
  reg        casez_tmp_9;
  reg        casez_tmp_10;
  reg        casez_tmp_11;
  reg        casez_tmp_12;
  reg  [6:0] casez_tmp_13;
  reg        casez_tmp_14;
  reg        casez_tmp_15;
  reg        casez_tmp_16;
  reg  [6:0] casez_tmp_17;
  reg        casez_tmp_18;
  reg        casez_tmp_19;
  reg        casez_tmp_20;
  reg  [6:0] casez_tmp_21;
  reg        casez_tmp_22;
  reg        casez_tmp_23;
  reg        casez_tmp_24;
  reg  [6:0] casez_tmp_25;
  reg        casez_tmp_26;
  reg        casez_tmp_27;
  reg        casez_tmp_28;
  reg  [6:0] casez_tmp_29;
  reg        casez_tmp_30;
  reg        casez_tmp_31;
  reg        casez_tmp_32;
  reg  [6:0] casez_tmp_33;
  reg        casez_tmp_34;
  reg        casez_tmp_35;
  reg        casez_tmp_36;
  reg  [6:0] casez_tmp_37;
  reg        casez_tmp_38;
  reg        casez_tmp_39;
  reg        casez_tmp_40;
  reg  [6:0] casez_tmp_41;
  reg        casez_tmp_42;
  reg        casez_tmp_43;
  reg        casez_tmp_44;
  reg  [6:0] casez_tmp_45;
  reg        casez_tmp_46;
  reg        casez_tmp_47;
  reg        casez_tmp_48;
  reg  [6:0] casez_tmp_49;
  reg        casez_tmp_50;
  reg        casez_tmp_51;
  reg        casez_tmp_52;
  reg        casez_tmp_53;
  reg        casez_tmp_54;
  reg        casez_tmp_55;
  reg        casez_tmp_56;
  reg        casez_tmp_57;
  reg        casez_tmp_58;
  reg        casez_tmp_59;
  reg        casez_tmp_60;
  reg        casez_tmp_61;
  reg        casez_tmp_62;
  reg        casez_tmp_63;
  reg  [6:0] casez_tmp_64;
  reg        casez_tmp_65;
  reg        casez_tmp_66;
  reg        casez_tmp_67;
  reg  [6:0] casez_tmp_68;
  reg        casez_tmp_69;
  reg        casez_tmp_70;
  reg        casez_tmp_71;
  reg  [6:0] casez_tmp_72;
  reg        casez_tmp_73;
  reg        casez_tmp_74;
  reg        casez_tmp_75;
  reg  [6:0] casez_tmp_76;
  reg        casez_tmp_77;
  reg        casez_tmp_78;
  reg        casez_tmp_79;
  reg  [6:0] casez_tmp_80;
  reg        casez_tmp_81;
  reg        casez_tmp_82;
  reg        casez_tmp_83;
  reg  [6:0] casez_tmp_84;
  reg        casez_tmp_85;
  reg        casez_tmp_86;
  reg        casez_tmp_87;
  reg  [6:0] casez_tmp_88;
  reg        casez_tmp_89;
  reg        casez_tmp_90;
  reg        casez_tmp_91;
  reg  [6:0] casez_tmp_92;
  reg        casez_tmp_93;
  reg        casez_tmp_94;
  reg        casez_tmp_95;
  reg  [6:0] casez_tmp_96;
  reg        casez_tmp_97;
  reg        casez_tmp_98;
  reg        casez_tmp_99;
  reg  [6:0] casez_tmp_100;
  reg        casez_tmp_101;
  reg        casez_tmp_102;
  reg        casez_tmp_103;
  reg        casez_tmp_104;
  reg        casez_tmp_105;
  reg        casez_tmp_106;
  reg        casez_tmp_107;
  reg        casez_tmp_108;
  reg        casez_tmp_109;
  reg        casez_tmp_110;
  reg        casez_tmp_111;
  reg        casez_tmp_112;
  reg        casez_tmp_113;
  reg        casez_tmp_114;
  reg  [6:0] casez_tmp_115;
  reg        casez_tmp_116;
  reg        casez_tmp_117;
  reg        casez_tmp_118;
  reg  [6:0] casez_tmp_119;
  reg        casez_tmp_120;
  reg        casez_tmp_121;
  reg        casez_tmp_122;
  reg  [6:0] casez_tmp_123;
  reg        casez_tmp_124;
  reg        casez_tmp_125;
  reg        casez_tmp_126;
  reg  [6:0] casez_tmp_127;
  reg        casez_tmp_128;
  reg        casez_tmp_129;
  reg        casez_tmp_130;
  reg  [6:0] casez_tmp_131;
  reg        casez_tmp_132;
  reg        casez_tmp_133;
  reg        casez_tmp_134;
  reg  [6:0] casez_tmp_135;
  reg        casez_tmp_136;
  reg        casez_tmp_137;
  reg        casez_tmp_138;
  reg  [6:0] casez_tmp_139;
  reg        casez_tmp_140;
  reg        casez_tmp_141;
  reg        casez_tmp_142;
  reg  [6:0] casez_tmp_143;
  reg        casez_tmp_144;
  reg        casez_tmp_145;
  reg        casez_tmp_146;
  reg  [6:0] casez_tmp_147;
  reg        casez_tmp_148;
  reg        casez_tmp_149;
  reg        casez_tmp_150;
  reg  [6:0] casez_tmp_151;
  reg        casez_tmp_152;
  reg        casez_tmp_153;
  reg        casez_tmp_154;
  reg        casez_tmp_155;
  reg        casez_tmp_156;
  reg        casez_tmp_157;
  reg        casez_tmp_158;
  reg        casez_tmp_159;
  reg        casez_tmp_160;
  reg        casez_tmp_161;
  reg        casez_tmp_162;
  reg        casez_tmp_163;
  reg        casez_tmp_164;
  reg        casez_tmp_165;
  reg  [6:0] casez_tmp_166;
  reg        casez_tmp_167;
  reg        casez_tmp_168;
  reg        casez_tmp_169;
  reg  [6:0] casez_tmp_170;
  reg        casez_tmp_171;
  reg        casez_tmp_172;
  reg        casez_tmp_173;
  reg  [6:0] casez_tmp_174;
  reg        casez_tmp_175;
  reg        casez_tmp_176;
  reg        casez_tmp_177;
  reg  [6:0] casez_tmp_178;
  reg        casez_tmp_179;
  reg        casez_tmp_180;
  reg        casez_tmp_181;
  reg  [6:0] casez_tmp_182;
  reg        casez_tmp_183;
  reg        casez_tmp_184;
  reg        casez_tmp_185;
  reg  [6:0] casez_tmp_186;
  reg        casez_tmp_187;
  reg        casez_tmp_188;
  reg        casez_tmp_189;
  reg  [6:0] casez_tmp_190;
  reg        casez_tmp_191;
  reg        casez_tmp_192;
  reg        casez_tmp_193;
  reg  [6:0] casez_tmp_194;
  reg        casez_tmp_195;
  reg        casez_tmp_196;
  reg        casez_tmp_197;
  reg  [6:0] casez_tmp_198;
  reg        casez_tmp_199;
  reg        casez_tmp_200;
  reg        casez_tmp_201;
  reg  [6:0] casez_tmp_202;
  reg  [4:0] rob_pnr;
  reg  [1:0] rob_pnr_lsb;
  wire [6:0] rob_pnr_idx = {rob_pnr, rob_pnr_lsb};
  reg        rob_unsafe__0;
  reg        rob_unsafe__1;
  reg        rob_unsafe__2;
  reg        rob_unsafe__3;
  reg        rob_unsafe__4;
  reg        rob_unsafe__5;
  reg        rob_unsafe__6;
  reg        rob_unsafe__7;
  reg        rob_unsafe__8;
  reg        rob_unsafe__9;
  reg        rob_unsafe__10;
  reg        rob_unsafe__11;
  reg        rob_unsafe__12;
  reg        rob_unsafe__13;
  reg        rob_unsafe__14;
  reg        rob_unsafe__15;
  reg        rob_unsafe__16;
  reg        rob_unsafe__17;
  reg        rob_unsafe__18;
  reg        rob_unsafe__19;
  reg        rob_unsafe__20;
  reg        rob_unsafe__21;
  reg        rob_unsafe__22;
  reg        rob_unsafe__23;
  reg        rob_unsafe__24;
  reg        rob_unsafe__25;
  reg        rob_unsafe__26;
  reg        rob_unsafe__27;
  reg        rob_unsafe__28;
  reg        rob_unsafe__29;
  reg        rob_unsafe__30;
  reg        rob_unsafe__31;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp = rob_val__0;
      5'b00001:
        casez_tmp = rob_val__1;
      5'b00010:
        casez_tmp = rob_val__2;
      5'b00011:
        casez_tmp = rob_val__3;
      5'b00100:
        casez_tmp = rob_val__4;
      5'b00101:
        casez_tmp = rob_val__5;
      5'b00110:
        casez_tmp = rob_val__6;
      5'b00111:
        casez_tmp = rob_val__7;
      5'b01000:
        casez_tmp = rob_val__8;
      5'b01001:
        casez_tmp = rob_val__9;
      5'b01010:
        casez_tmp = rob_val__10;
      5'b01011:
        casez_tmp = rob_val__11;
      5'b01100:
        casez_tmp = rob_val__12;
      5'b01101:
        casez_tmp = rob_val__13;
      5'b01110:
        casez_tmp = rob_val__14;
      5'b01111:
        casez_tmp = rob_val__15;
      5'b10000:
        casez_tmp = rob_val__16;
      5'b10001:
        casez_tmp = rob_val__17;
      5'b10010:
        casez_tmp = rob_val__18;
      5'b10011:
        casez_tmp = rob_val__19;
      5'b10100:
        casez_tmp = rob_val__20;
      5'b10101:
        casez_tmp = rob_val__21;
      5'b10110:
        casez_tmp = rob_val__22;
      5'b10111:
        casez_tmp = rob_val__23;
      5'b11000:
        casez_tmp = rob_val__24;
      5'b11001:
        casez_tmp = rob_val__25;
      5'b11010:
        casez_tmp = rob_val__26;
      5'b11011:
        casez_tmp = rob_val__27;
      5'b11100:
        casez_tmp = rob_val__28;
      5'b11101:
        casez_tmp = rob_val__29;
      5'b11110:
        casez_tmp = rob_val__30;
      default:
        casez_tmp = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1852 = io_enq_uops_0_rob_idx[6:2] == rob_tail;
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_0 = rob_val__0;
      5'b00001:
        casez_tmp_0 = rob_val__1;
      5'b00010:
        casez_tmp_0 = rob_val__2;
      5'b00011:
        casez_tmp_0 = rob_val__3;
      5'b00100:
        casez_tmp_0 = rob_val__4;
      5'b00101:
        casez_tmp_0 = rob_val__5;
      5'b00110:
        casez_tmp_0 = rob_val__6;
      5'b00111:
        casez_tmp_0 = rob_val__7;
      5'b01000:
        casez_tmp_0 = rob_val__8;
      5'b01001:
        casez_tmp_0 = rob_val__9;
      5'b01010:
        casez_tmp_0 = rob_val__10;
      5'b01011:
        casez_tmp_0 = rob_val__11;
      5'b01100:
        casez_tmp_0 = rob_val__12;
      5'b01101:
        casez_tmp_0 = rob_val__13;
      5'b01110:
        casez_tmp_0 = rob_val__14;
      5'b01111:
        casez_tmp_0 = rob_val__15;
      5'b10000:
        casez_tmp_0 = rob_val__16;
      5'b10001:
        casez_tmp_0 = rob_val__17;
      5'b10010:
        casez_tmp_0 = rob_val__18;
      5'b10011:
        casez_tmp_0 = rob_val__19;
      5'b10100:
        casez_tmp_0 = rob_val__20;
      5'b10101:
        casez_tmp_0 = rob_val__21;
      5'b10110:
        casez_tmp_0 = rob_val__22;
      5'b10111:
        casez_tmp_0 = rob_val__23;
      5'b11000:
        casez_tmp_0 = rob_val__24;
      5'b11001:
        casez_tmp_0 = rob_val__25;
      5'b11010:
        casez_tmp_0 = rob_val__26;
      5'b11011:
        casez_tmp_0 = rob_val__27;
      5'b11100:
        casez_tmp_0 = rob_val__28;
      5'b11101:
        casez_tmp_0 = rob_val__29;
      5'b11110:
        casez_tmp_0 = rob_val__30;
      default:
        casez_tmp_0 = rob_val__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_1 = rob_bsy__0;
      5'b00001:
        casez_tmp_1 = rob_bsy__1;
      5'b00010:
        casez_tmp_1 = rob_bsy__2;
      5'b00011:
        casez_tmp_1 = rob_bsy__3;
      5'b00100:
        casez_tmp_1 = rob_bsy__4;
      5'b00101:
        casez_tmp_1 = rob_bsy__5;
      5'b00110:
        casez_tmp_1 = rob_bsy__6;
      5'b00111:
        casez_tmp_1 = rob_bsy__7;
      5'b01000:
        casez_tmp_1 = rob_bsy__8;
      5'b01001:
        casez_tmp_1 = rob_bsy__9;
      5'b01010:
        casez_tmp_1 = rob_bsy__10;
      5'b01011:
        casez_tmp_1 = rob_bsy__11;
      5'b01100:
        casez_tmp_1 = rob_bsy__12;
      5'b01101:
        casez_tmp_1 = rob_bsy__13;
      5'b01110:
        casez_tmp_1 = rob_bsy__14;
      5'b01111:
        casez_tmp_1 = rob_bsy__15;
      5'b10000:
        casez_tmp_1 = rob_bsy__16;
      5'b10001:
        casez_tmp_1 = rob_bsy__17;
      5'b10010:
        casez_tmp_1 = rob_bsy__18;
      5'b10011:
        casez_tmp_1 = rob_bsy__19;
      5'b10100:
        casez_tmp_1 = rob_bsy__20;
      5'b10101:
        casez_tmp_1 = rob_bsy__21;
      5'b10110:
        casez_tmp_1 = rob_bsy__22;
      5'b10111:
        casez_tmp_1 = rob_bsy__23;
      5'b11000:
        casez_tmp_1 = rob_bsy__24;
      5'b11001:
        casez_tmp_1 = rob_bsy__25;
      5'b11010:
        casez_tmp_1 = rob_bsy__26;
      5'b11011:
        casez_tmp_1 = rob_bsy__27;
      5'b11100:
        casez_tmp_1 = rob_bsy__28;
      5'b11101:
        casez_tmp_1 = rob_bsy__29;
      5'b11110:
        casez_tmp_1 = rob_bsy__30;
      default:
        casez_tmp_1 = rob_bsy__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_2 = rob_val__0;
      5'b00001:
        casez_tmp_2 = rob_val__1;
      5'b00010:
        casez_tmp_2 = rob_val__2;
      5'b00011:
        casez_tmp_2 = rob_val__3;
      5'b00100:
        casez_tmp_2 = rob_val__4;
      5'b00101:
        casez_tmp_2 = rob_val__5;
      5'b00110:
        casez_tmp_2 = rob_val__6;
      5'b00111:
        casez_tmp_2 = rob_val__7;
      5'b01000:
        casez_tmp_2 = rob_val__8;
      5'b01001:
        casez_tmp_2 = rob_val__9;
      5'b01010:
        casez_tmp_2 = rob_val__10;
      5'b01011:
        casez_tmp_2 = rob_val__11;
      5'b01100:
        casez_tmp_2 = rob_val__12;
      5'b01101:
        casez_tmp_2 = rob_val__13;
      5'b01110:
        casez_tmp_2 = rob_val__14;
      5'b01111:
        casez_tmp_2 = rob_val__15;
      5'b10000:
        casez_tmp_2 = rob_val__16;
      5'b10001:
        casez_tmp_2 = rob_val__17;
      5'b10010:
        casez_tmp_2 = rob_val__18;
      5'b10011:
        casez_tmp_2 = rob_val__19;
      5'b10100:
        casez_tmp_2 = rob_val__20;
      5'b10101:
        casez_tmp_2 = rob_val__21;
      5'b10110:
        casez_tmp_2 = rob_val__22;
      5'b10111:
        casez_tmp_2 = rob_val__23;
      5'b11000:
        casez_tmp_2 = rob_val__24;
      5'b11001:
        casez_tmp_2 = rob_val__25;
      5'b11010:
        casez_tmp_2 = rob_val__26;
      5'b11011:
        casez_tmp_2 = rob_val__27;
      5'b11100:
        casez_tmp_2 = rob_val__28;
      5'b11101:
        casez_tmp_2 = rob_val__29;
      5'b11110:
        casez_tmp_2 = rob_val__30;
      default:
        casez_tmp_2 = rob_val__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_3 = rob_bsy__0;
      5'b00001:
        casez_tmp_3 = rob_bsy__1;
      5'b00010:
        casez_tmp_3 = rob_bsy__2;
      5'b00011:
        casez_tmp_3 = rob_bsy__3;
      5'b00100:
        casez_tmp_3 = rob_bsy__4;
      5'b00101:
        casez_tmp_3 = rob_bsy__5;
      5'b00110:
        casez_tmp_3 = rob_bsy__6;
      5'b00111:
        casez_tmp_3 = rob_bsy__7;
      5'b01000:
        casez_tmp_3 = rob_bsy__8;
      5'b01001:
        casez_tmp_3 = rob_bsy__9;
      5'b01010:
        casez_tmp_3 = rob_bsy__10;
      5'b01011:
        casez_tmp_3 = rob_bsy__11;
      5'b01100:
        casez_tmp_3 = rob_bsy__12;
      5'b01101:
        casez_tmp_3 = rob_bsy__13;
      5'b01110:
        casez_tmp_3 = rob_bsy__14;
      5'b01111:
        casez_tmp_3 = rob_bsy__15;
      5'b10000:
        casez_tmp_3 = rob_bsy__16;
      5'b10001:
        casez_tmp_3 = rob_bsy__17;
      5'b10010:
        casez_tmp_3 = rob_bsy__18;
      5'b10011:
        casez_tmp_3 = rob_bsy__19;
      5'b10100:
        casez_tmp_3 = rob_bsy__20;
      5'b10101:
        casez_tmp_3 = rob_bsy__21;
      5'b10110:
        casez_tmp_3 = rob_bsy__22;
      5'b10111:
        casez_tmp_3 = rob_bsy__23;
      5'b11000:
        casez_tmp_3 = rob_bsy__24;
      5'b11001:
        casez_tmp_3 = rob_bsy__25;
      5'b11010:
        casez_tmp_3 = rob_bsy__26;
      5'b11011:
        casez_tmp_3 = rob_bsy__27;
      5'b11100:
        casez_tmp_3 = rob_bsy__28;
      5'b11101:
        casez_tmp_3 = rob_bsy__29;
      5'b11110:
        casez_tmp_3 = rob_bsy__30;
      default:
        casez_tmp_3 = rob_bsy__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_4 = rob_val__0;
      5'b00001:
        casez_tmp_4 = rob_val__1;
      5'b00010:
        casez_tmp_4 = rob_val__2;
      5'b00011:
        casez_tmp_4 = rob_val__3;
      5'b00100:
        casez_tmp_4 = rob_val__4;
      5'b00101:
        casez_tmp_4 = rob_val__5;
      5'b00110:
        casez_tmp_4 = rob_val__6;
      5'b00111:
        casez_tmp_4 = rob_val__7;
      5'b01000:
        casez_tmp_4 = rob_val__8;
      5'b01001:
        casez_tmp_4 = rob_val__9;
      5'b01010:
        casez_tmp_4 = rob_val__10;
      5'b01011:
        casez_tmp_4 = rob_val__11;
      5'b01100:
        casez_tmp_4 = rob_val__12;
      5'b01101:
        casez_tmp_4 = rob_val__13;
      5'b01110:
        casez_tmp_4 = rob_val__14;
      5'b01111:
        casez_tmp_4 = rob_val__15;
      5'b10000:
        casez_tmp_4 = rob_val__16;
      5'b10001:
        casez_tmp_4 = rob_val__17;
      5'b10010:
        casez_tmp_4 = rob_val__18;
      5'b10011:
        casez_tmp_4 = rob_val__19;
      5'b10100:
        casez_tmp_4 = rob_val__20;
      5'b10101:
        casez_tmp_4 = rob_val__21;
      5'b10110:
        casez_tmp_4 = rob_val__22;
      5'b10111:
        casez_tmp_4 = rob_val__23;
      5'b11000:
        casez_tmp_4 = rob_val__24;
      5'b11001:
        casez_tmp_4 = rob_val__25;
      5'b11010:
        casez_tmp_4 = rob_val__26;
      5'b11011:
        casez_tmp_4 = rob_val__27;
      5'b11100:
        casez_tmp_4 = rob_val__28;
      5'b11101:
        casez_tmp_4 = rob_val__29;
      5'b11110:
        casez_tmp_4 = rob_val__30;
      default:
        casez_tmp_4 = rob_val__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_5 = rob_bsy__0;
      5'b00001:
        casez_tmp_5 = rob_bsy__1;
      5'b00010:
        casez_tmp_5 = rob_bsy__2;
      5'b00011:
        casez_tmp_5 = rob_bsy__3;
      5'b00100:
        casez_tmp_5 = rob_bsy__4;
      5'b00101:
        casez_tmp_5 = rob_bsy__5;
      5'b00110:
        casez_tmp_5 = rob_bsy__6;
      5'b00111:
        casez_tmp_5 = rob_bsy__7;
      5'b01000:
        casez_tmp_5 = rob_bsy__8;
      5'b01001:
        casez_tmp_5 = rob_bsy__9;
      5'b01010:
        casez_tmp_5 = rob_bsy__10;
      5'b01011:
        casez_tmp_5 = rob_bsy__11;
      5'b01100:
        casez_tmp_5 = rob_bsy__12;
      5'b01101:
        casez_tmp_5 = rob_bsy__13;
      5'b01110:
        casez_tmp_5 = rob_bsy__14;
      5'b01111:
        casez_tmp_5 = rob_bsy__15;
      5'b10000:
        casez_tmp_5 = rob_bsy__16;
      5'b10001:
        casez_tmp_5 = rob_bsy__17;
      5'b10010:
        casez_tmp_5 = rob_bsy__18;
      5'b10011:
        casez_tmp_5 = rob_bsy__19;
      5'b10100:
        casez_tmp_5 = rob_bsy__20;
      5'b10101:
        casez_tmp_5 = rob_bsy__21;
      5'b10110:
        casez_tmp_5 = rob_bsy__22;
      5'b10111:
        casez_tmp_5 = rob_bsy__23;
      5'b11000:
        casez_tmp_5 = rob_bsy__24;
      5'b11001:
        casez_tmp_5 = rob_bsy__25;
      5'b11010:
        casez_tmp_5 = rob_bsy__26;
      5'b11011:
        casez_tmp_5 = rob_bsy__27;
      5'b11100:
        casez_tmp_5 = rob_bsy__28;
      5'b11101:
        casez_tmp_5 = rob_bsy__29;
      5'b11110:
        casez_tmp_5 = rob_bsy__30;
      default:
        casez_tmp_5 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1853 = io_lxcpt_bits_cause != 5'h10;
  always @(*) begin
    casez (_GEN_2)
      5'b00000:
        casez_tmp_6 = rob_unsafe__0;
      5'b00001:
        casez_tmp_6 = rob_unsafe__1;
      5'b00010:
        casez_tmp_6 = rob_unsafe__2;
      5'b00011:
        casez_tmp_6 = rob_unsafe__3;
      5'b00100:
        casez_tmp_6 = rob_unsafe__4;
      5'b00101:
        casez_tmp_6 = rob_unsafe__5;
      5'b00110:
        casez_tmp_6 = rob_unsafe__6;
      5'b00111:
        casez_tmp_6 = rob_unsafe__7;
      5'b01000:
        casez_tmp_6 = rob_unsafe__8;
      5'b01001:
        casez_tmp_6 = rob_unsafe__9;
      5'b01010:
        casez_tmp_6 = rob_unsafe__10;
      5'b01011:
        casez_tmp_6 = rob_unsafe__11;
      5'b01100:
        casez_tmp_6 = rob_unsafe__12;
      5'b01101:
        casez_tmp_6 = rob_unsafe__13;
      5'b01110:
        casez_tmp_6 = rob_unsafe__14;
      5'b01111:
        casez_tmp_6 = rob_unsafe__15;
      5'b10000:
        casez_tmp_6 = rob_unsafe__16;
      5'b10001:
        casez_tmp_6 = rob_unsafe__17;
      5'b10010:
        casez_tmp_6 = rob_unsafe__18;
      5'b10011:
        casez_tmp_6 = rob_unsafe__19;
      5'b10100:
        casez_tmp_6 = rob_unsafe__20;
      5'b10101:
        casez_tmp_6 = rob_unsafe__21;
      5'b10110:
        casez_tmp_6 = rob_unsafe__22;
      5'b10111:
        casez_tmp_6 = rob_unsafe__23;
      5'b11000:
        casez_tmp_6 = rob_unsafe__24;
      5'b11001:
        casez_tmp_6 = rob_unsafe__25;
      5'b11010:
        casez_tmp_6 = rob_unsafe__26;
      5'b11011:
        casez_tmp_6 = rob_unsafe__27;
      5'b11100:
        casez_tmp_6 = rob_unsafe__28;
      5'b11101:
        casez_tmp_6 = rob_unsafe__29;
      5'b11110:
        casez_tmp_6 = rob_unsafe__30;
      default:
        casez_tmp_6 = rob_unsafe__31;
    endcase
  end // always @(*)
  wire       _GEN_1854 = (_io_commit_valids_0_output | _io_commit_valids_1_output | _io_commit_valids_2_output | _io_commit_valids_3_output) & (_io_commit_rbk_valids_0_output | _io_commit_rbk_valids_1_output | _io_commit_rbk_valids_2_output | _io_commit_rbk_valids_3_output);
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_7 = rob_unsafe__0;
      5'b00001:
        casez_tmp_7 = rob_unsafe__1;
      5'b00010:
        casez_tmp_7 = rob_unsafe__2;
      5'b00011:
        casez_tmp_7 = rob_unsafe__3;
      5'b00100:
        casez_tmp_7 = rob_unsafe__4;
      5'b00101:
        casez_tmp_7 = rob_unsafe__5;
      5'b00110:
        casez_tmp_7 = rob_unsafe__6;
      5'b00111:
        casez_tmp_7 = rob_unsafe__7;
      5'b01000:
        casez_tmp_7 = rob_unsafe__8;
      5'b01001:
        casez_tmp_7 = rob_unsafe__9;
      5'b01010:
        casez_tmp_7 = rob_unsafe__10;
      5'b01011:
        casez_tmp_7 = rob_unsafe__11;
      5'b01100:
        casez_tmp_7 = rob_unsafe__12;
      5'b01101:
        casez_tmp_7 = rob_unsafe__13;
      5'b01110:
        casez_tmp_7 = rob_unsafe__14;
      5'b01111:
        casez_tmp_7 = rob_unsafe__15;
      5'b10000:
        casez_tmp_7 = rob_unsafe__16;
      5'b10001:
        casez_tmp_7 = rob_unsafe__17;
      5'b10010:
        casez_tmp_7 = rob_unsafe__18;
      5'b10011:
        casez_tmp_7 = rob_unsafe__19;
      5'b10100:
        casez_tmp_7 = rob_unsafe__20;
      5'b10101:
        casez_tmp_7 = rob_unsafe__21;
      5'b10110:
        casez_tmp_7 = rob_unsafe__22;
      5'b10111:
        casez_tmp_7 = rob_unsafe__23;
      5'b11000:
        casez_tmp_7 = rob_unsafe__24;
      5'b11001:
        casez_tmp_7 = rob_unsafe__25;
      5'b11010:
        casez_tmp_7 = rob_unsafe__26;
      5'b11011:
        casez_tmp_7 = rob_unsafe__27;
      5'b11100:
        casez_tmp_7 = rob_unsafe__28;
      5'b11101:
        casez_tmp_7 = rob_unsafe__29;
      5'b11110:
        casez_tmp_7 = rob_unsafe__30;
      default:
        casez_tmp_7 = rob_unsafe__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_8 = rob_exception__0;
      5'b00001:
        casez_tmp_8 = rob_exception__1;
      5'b00010:
        casez_tmp_8 = rob_exception__2;
      5'b00011:
        casez_tmp_8 = rob_exception__3;
      5'b00100:
        casez_tmp_8 = rob_exception__4;
      5'b00101:
        casez_tmp_8 = rob_exception__5;
      5'b00110:
        casez_tmp_8 = rob_exception__6;
      5'b00111:
        casez_tmp_8 = rob_exception__7;
      5'b01000:
        casez_tmp_8 = rob_exception__8;
      5'b01001:
        casez_tmp_8 = rob_exception__9;
      5'b01010:
        casez_tmp_8 = rob_exception__10;
      5'b01011:
        casez_tmp_8 = rob_exception__11;
      5'b01100:
        casez_tmp_8 = rob_exception__12;
      5'b01101:
        casez_tmp_8 = rob_exception__13;
      5'b01110:
        casez_tmp_8 = rob_exception__14;
      5'b01111:
        casez_tmp_8 = rob_exception__15;
      5'b10000:
        casez_tmp_8 = rob_exception__16;
      5'b10001:
        casez_tmp_8 = rob_exception__17;
      5'b10010:
        casez_tmp_8 = rob_exception__18;
      5'b10011:
        casez_tmp_8 = rob_exception__19;
      5'b10100:
        casez_tmp_8 = rob_exception__20;
      5'b10101:
        casez_tmp_8 = rob_exception__21;
      5'b10110:
        casez_tmp_8 = rob_exception__22;
      5'b10111:
        casez_tmp_8 = rob_exception__23;
      5'b11000:
        casez_tmp_8 = rob_exception__24;
      5'b11001:
        casez_tmp_8 = rob_exception__25;
      5'b11010:
        casez_tmp_8 = rob_exception__26;
      5'b11011:
        casez_tmp_8 = rob_exception__27;
      5'b11100:
        casez_tmp_8 = rob_exception__28;
      5'b11101:
        casez_tmp_8 = rob_exception__29;
      5'b11110:
        casez_tmp_8 = rob_exception__30;
      default:
        casez_tmp_8 = rob_exception__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_9 = rob_val__0;
      5'b00001:
        casez_tmp_9 = rob_val__1;
      5'b00010:
        casez_tmp_9 = rob_val__2;
      5'b00011:
        casez_tmp_9 = rob_val__3;
      5'b00100:
        casez_tmp_9 = rob_val__4;
      5'b00101:
        casez_tmp_9 = rob_val__5;
      5'b00110:
        casez_tmp_9 = rob_val__6;
      5'b00111:
        casez_tmp_9 = rob_val__7;
      5'b01000:
        casez_tmp_9 = rob_val__8;
      5'b01001:
        casez_tmp_9 = rob_val__9;
      5'b01010:
        casez_tmp_9 = rob_val__10;
      5'b01011:
        casez_tmp_9 = rob_val__11;
      5'b01100:
        casez_tmp_9 = rob_val__12;
      5'b01101:
        casez_tmp_9 = rob_val__13;
      5'b01110:
        casez_tmp_9 = rob_val__14;
      5'b01111:
        casez_tmp_9 = rob_val__15;
      5'b10000:
        casez_tmp_9 = rob_val__16;
      5'b10001:
        casez_tmp_9 = rob_val__17;
      5'b10010:
        casez_tmp_9 = rob_val__18;
      5'b10011:
        casez_tmp_9 = rob_val__19;
      5'b10100:
        casez_tmp_9 = rob_val__20;
      5'b10101:
        casez_tmp_9 = rob_val__21;
      5'b10110:
        casez_tmp_9 = rob_val__22;
      5'b10111:
        casez_tmp_9 = rob_val__23;
      5'b11000:
        casez_tmp_9 = rob_val__24;
      5'b11001:
        casez_tmp_9 = rob_val__25;
      5'b11010:
        casez_tmp_9 = rob_val__26;
      5'b11011:
        casez_tmp_9 = rob_val__27;
      5'b11100:
        casez_tmp_9 = rob_val__28;
      5'b11101:
        casez_tmp_9 = rob_val__29;
      5'b11110:
        casez_tmp_9 = rob_val__30;
      default:
        casez_tmp_9 = rob_val__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_10 = rob_val__0;
      5'b00001:
        casez_tmp_10 = rob_val__1;
      5'b00010:
        casez_tmp_10 = rob_val__2;
      5'b00011:
        casez_tmp_10 = rob_val__3;
      5'b00100:
        casez_tmp_10 = rob_val__4;
      5'b00101:
        casez_tmp_10 = rob_val__5;
      5'b00110:
        casez_tmp_10 = rob_val__6;
      5'b00111:
        casez_tmp_10 = rob_val__7;
      5'b01000:
        casez_tmp_10 = rob_val__8;
      5'b01001:
        casez_tmp_10 = rob_val__9;
      5'b01010:
        casez_tmp_10 = rob_val__10;
      5'b01011:
        casez_tmp_10 = rob_val__11;
      5'b01100:
        casez_tmp_10 = rob_val__12;
      5'b01101:
        casez_tmp_10 = rob_val__13;
      5'b01110:
        casez_tmp_10 = rob_val__14;
      5'b01111:
        casez_tmp_10 = rob_val__15;
      5'b10000:
        casez_tmp_10 = rob_val__16;
      5'b10001:
        casez_tmp_10 = rob_val__17;
      5'b10010:
        casez_tmp_10 = rob_val__18;
      5'b10011:
        casez_tmp_10 = rob_val__19;
      5'b10100:
        casez_tmp_10 = rob_val__20;
      5'b10101:
        casez_tmp_10 = rob_val__21;
      5'b10110:
        casez_tmp_10 = rob_val__22;
      5'b10111:
        casez_tmp_10 = rob_val__23;
      5'b11000:
        casez_tmp_10 = rob_val__24;
      5'b11001:
        casez_tmp_10 = rob_val__25;
      5'b11010:
        casez_tmp_10 = rob_val__26;
      5'b11011:
        casez_tmp_10 = rob_val__27;
      5'b11100:
        casez_tmp_10 = rob_val__28;
      5'b11101:
        casez_tmp_10 = rob_val__29;
      5'b11110:
        casez_tmp_10 = rob_val__30;
      default:
        casez_tmp_10 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1855 = _GEN_457 & ~casez_tmp_10;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_11 = rob_bsy__0;
      5'b00001:
        casez_tmp_11 = rob_bsy__1;
      5'b00010:
        casez_tmp_11 = rob_bsy__2;
      5'b00011:
        casez_tmp_11 = rob_bsy__3;
      5'b00100:
        casez_tmp_11 = rob_bsy__4;
      5'b00101:
        casez_tmp_11 = rob_bsy__5;
      5'b00110:
        casez_tmp_11 = rob_bsy__6;
      5'b00111:
        casez_tmp_11 = rob_bsy__7;
      5'b01000:
        casez_tmp_11 = rob_bsy__8;
      5'b01001:
        casez_tmp_11 = rob_bsy__9;
      5'b01010:
        casez_tmp_11 = rob_bsy__10;
      5'b01011:
        casez_tmp_11 = rob_bsy__11;
      5'b01100:
        casez_tmp_11 = rob_bsy__12;
      5'b01101:
        casez_tmp_11 = rob_bsy__13;
      5'b01110:
        casez_tmp_11 = rob_bsy__14;
      5'b01111:
        casez_tmp_11 = rob_bsy__15;
      5'b10000:
        casez_tmp_11 = rob_bsy__16;
      5'b10001:
        casez_tmp_11 = rob_bsy__17;
      5'b10010:
        casez_tmp_11 = rob_bsy__18;
      5'b10011:
        casez_tmp_11 = rob_bsy__19;
      5'b10100:
        casez_tmp_11 = rob_bsy__20;
      5'b10101:
        casez_tmp_11 = rob_bsy__21;
      5'b10110:
        casez_tmp_11 = rob_bsy__22;
      5'b10111:
        casez_tmp_11 = rob_bsy__23;
      5'b11000:
        casez_tmp_11 = rob_bsy__24;
      5'b11001:
        casez_tmp_11 = rob_bsy__25;
      5'b11010:
        casez_tmp_11 = rob_bsy__26;
      5'b11011:
        casez_tmp_11 = rob_bsy__27;
      5'b11100:
        casez_tmp_11 = rob_bsy__28;
      5'b11101:
        casez_tmp_11 = rob_bsy__29;
      5'b11110:
        casez_tmp_11 = rob_bsy__30;
      default:
        casez_tmp_11 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1856 = _GEN_457 & ~casez_tmp_11;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_12 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_12 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_12 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_12 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_12 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_12 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_12 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_12 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_12 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_12 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_12 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_12 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_12 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_12 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_12 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_12 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_12 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_12 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_12 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_12 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_12 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_12 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_12 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_12 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_12 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_12 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_12 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_12 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_12 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_12 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_12 = rob_uop__30_ldst_val;
      default:
        casez_tmp_12 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_13 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_13 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_13 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_13 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_13 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_13 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_13 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_13 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_13 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_13 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_13 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_13 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_13 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_13 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_13 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_13 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_13 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_13 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_13 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_13 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_13 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_13 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_13 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_13 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_13 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_13 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_13 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_13 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_13 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_13 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_13 = rob_uop__30_pdst;
      default:
        casez_tmp_13 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1857 = _GEN_457 & casez_tmp_12 & casez_tmp_13 != io_wb_resps_0_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_14 = rob_val__0;
      5'b00001:
        casez_tmp_14 = rob_val__1;
      5'b00010:
        casez_tmp_14 = rob_val__2;
      5'b00011:
        casez_tmp_14 = rob_val__3;
      5'b00100:
        casez_tmp_14 = rob_val__4;
      5'b00101:
        casez_tmp_14 = rob_val__5;
      5'b00110:
        casez_tmp_14 = rob_val__6;
      5'b00111:
        casez_tmp_14 = rob_val__7;
      5'b01000:
        casez_tmp_14 = rob_val__8;
      5'b01001:
        casez_tmp_14 = rob_val__9;
      5'b01010:
        casez_tmp_14 = rob_val__10;
      5'b01011:
        casez_tmp_14 = rob_val__11;
      5'b01100:
        casez_tmp_14 = rob_val__12;
      5'b01101:
        casez_tmp_14 = rob_val__13;
      5'b01110:
        casez_tmp_14 = rob_val__14;
      5'b01111:
        casez_tmp_14 = rob_val__15;
      5'b10000:
        casez_tmp_14 = rob_val__16;
      5'b10001:
        casez_tmp_14 = rob_val__17;
      5'b10010:
        casez_tmp_14 = rob_val__18;
      5'b10011:
        casez_tmp_14 = rob_val__19;
      5'b10100:
        casez_tmp_14 = rob_val__20;
      5'b10101:
        casez_tmp_14 = rob_val__21;
      5'b10110:
        casez_tmp_14 = rob_val__22;
      5'b10111:
        casez_tmp_14 = rob_val__23;
      5'b11000:
        casez_tmp_14 = rob_val__24;
      5'b11001:
        casez_tmp_14 = rob_val__25;
      5'b11010:
        casez_tmp_14 = rob_val__26;
      5'b11011:
        casez_tmp_14 = rob_val__27;
      5'b11100:
        casez_tmp_14 = rob_val__28;
      5'b11101:
        casez_tmp_14 = rob_val__29;
      5'b11110:
        casez_tmp_14 = rob_val__30;
      default:
        casez_tmp_14 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1858 = _GEN_8 & ~casez_tmp_14;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_15 = rob_bsy__0;
      5'b00001:
        casez_tmp_15 = rob_bsy__1;
      5'b00010:
        casez_tmp_15 = rob_bsy__2;
      5'b00011:
        casez_tmp_15 = rob_bsy__3;
      5'b00100:
        casez_tmp_15 = rob_bsy__4;
      5'b00101:
        casez_tmp_15 = rob_bsy__5;
      5'b00110:
        casez_tmp_15 = rob_bsy__6;
      5'b00111:
        casez_tmp_15 = rob_bsy__7;
      5'b01000:
        casez_tmp_15 = rob_bsy__8;
      5'b01001:
        casez_tmp_15 = rob_bsy__9;
      5'b01010:
        casez_tmp_15 = rob_bsy__10;
      5'b01011:
        casez_tmp_15 = rob_bsy__11;
      5'b01100:
        casez_tmp_15 = rob_bsy__12;
      5'b01101:
        casez_tmp_15 = rob_bsy__13;
      5'b01110:
        casez_tmp_15 = rob_bsy__14;
      5'b01111:
        casez_tmp_15 = rob_bsy__15;
      5'b10000:
        casez_tmp_15 = rob_bsy__16;
      5'b10001:
        casez_tmp_15 = rob_bsy__17;
      5'b10010:
        casez_tmp_15 = rob_bsy__18;
      5'b10011:
        casez_tmp_15 = rob_bsy__19;
      5'b10100:
        casez_tmp_15 = rob_bsy__20;
      5'b10101:
        casez_tmp_15 = rob_bsy__21;
      5'b10110:
        casez_tmp_15 = rob_bsy__22;
      5'b10111:
        casez_tmp_15 = rob_bsy__23;
      5'b11000:
        casez_tmp_15 = rob_bsy__24;
      5'b11001:
        casez_tmp_15 = rob_bsy__25;
      5'b11010:
        casez_tmp_15 = rob_bsy__26;
      5'b11011:
        casez_tmp_15 = rob_bsy__27;
      5'b11100:
        casez_tmp_15 = rob_bsy__28;
      5'b11101:
        casez_tmp_15 = rob_bsy__29;
      5'b11110:
        casez_tmp_15 = rob_bsy__30;
      default:
        casez_tmp_15 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1859 = _GEN_8 & ~casez_tmp_15;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_16 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_16 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_16 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_16 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_16 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_16 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_16 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_16 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_16 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_16 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_16 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_16 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_16 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_16 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_16 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_16 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_16 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_16 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_16 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_16 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_16 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_16 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_16 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_16 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_16 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_16 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_16 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_16 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_16 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_16 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_16 = rob_uop__30_ldst_val;
      default:
        casez_tmp_16 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_17 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_17 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_17 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_17 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_17 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_17 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_17 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_17 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_17 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_17 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_17 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_17 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_17 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_17 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_17 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_17 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_17 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_17 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_17 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_17 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_17 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_17 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_17 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_17 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_17 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_17 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_17 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_17 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_17 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_17 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_17 = rob_uop__30_pdst;
      default:
        casez_tmp_17 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1860 = _GEN_8 & casez_tmp_16 & casez_tmp_17 != io_wb_resps_1_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_18 = rob_val__0;
      5'b00001:
        casez_tmp_18 = rob_val__1;
      5'b00010:
        casez_tmp_18 = rob_val__2;
      5'b00011:
        casez_tmp_18 = rob_val__3;
      5'b00100:
        casez_tmp_18 = rob_val__4;
      5'b00101:
        casez_tmp_18 = rob_val__5;
      5'b00110:
        casez_tmp_18 = rob_val__6;
      5'b00111:
        casez_tmp_18 = rob_val__7;
      5'b01000:
        casez_tmp_18 = rob_val__8;
      5'b01001:
        casez_tmp_18 = rob_val__9;
      5'b01010:
        casez_tmp_18 = rob_val__10;
      5'b01011:
        casez_tmp_18 = rob_val__11;
      5'b01100:
        casez_tmp_18 = rob_val__12;
      5'b01101:
        casez_tmp_18 = rob_val__13;
      5'b01110:
        casez_tmp_18 = rob_val__14;
      5'b01111:
        casez_tmp_18 = rob_val__15;
      5'b10000:
        casez_tmp_18 = rob_val__16;
      5'b10001:
        casez_tmp_18 = rob_val__17;
      5'b10010:
        casez_tmp_18 = rob_val__18;
      5'b10011:
        casez_tmp_18 = rob_val__19;
      5'b10100:
        casez_tmp_18 = rob_val__20;
      5'b10101:
        casez_tmp_18 = rob_val__21;
      5'b10110:
        casez_tmp_18 = rob_val__22;
      5'b10111:
        casez_tmp_18 = rob_val__23;
      5'b11000:
        casez_tmp_18 = rob_val__24;
      5'b11001:
        casez_tmp_18 = rob_val__25;
      5'b11010:
        casez_tmp_18 = rob_val__26;
      5'b11011:
        casez_tmp_18 = rob_val__27;
      5'b11100:
        casez_tmp_18 = rob_val__28;
      5'b11101:
        casez_tmp_18 = rob_val__29;
      5'b11110:
        casez_tmp_18 = rob_val__30;
      default:
        casez_tmp_18 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1861 = _GEN_458 & ~casez_tmp_18;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_19 = rob_bsy__0;
      5'b00001:
        casez_tmp_19 = rob_bsy__1;
      5'b00010:
        casez_tmp_19 = rob_bsy__2;
      5'b00011:
        casez_tmp_19 = rob_bsy__3;
      5'b00100:
        casez_tmp_19 = rob_bsy__4;
      5'b00101:
        casez_tmp_19 = rob_bsy__5;
      5'b00110:
        casez_tmp_19 = rob_bsy__6;
      5'b00111:
        casez_tmp_19 = rob_bsy__7;
      5'b01000:
        casez_tmp_19 = rob_bsy__8;
      5'b01001:
        casez_tmp_19 = rob_bsy__9;
      5'b01010:
        casez_tmp_19 = rob_bsy__10;
      5'b01011:
        casez_tmp_19 = rob_bsy__11;
      5'b01100:
        casez_tmp_19 = rob_bsy__12;
      5'b01101:
        casez_tmp_19 = rob_bsy__13;
      5'b01110:
        casez_tmp_19 = rob_bsy__14;
      5'b01111:
        casez_tmp_19 = rob_bsy__15;
      5'b10000:
        casez_tmp_19 = rob_bsy__16;
      5'b10001:
        casez_tmp_19 = rob_bsy__17;
      5'b10010:
        casez_tmp_19 = rob_bsy__18;
      5'b10011:
        casez_tmp_19 = rob_bsy__19;
      5'b10100:
        casez_tmp_19 = rob_bsy__20;
      5'b10101:
        casez_tmp_19 = rob_bsy__21;
      5'b10110:
        casez_tmp_19 = rob_bsy__22;
      5'b10111:
        casez_tmp_19 = rob_bsy__23;
      5'b11000:
        casez_tmp_19 = rob_bsy__24;
      5'b11001:
        casez_tmp_19 = rob_bsy__25;
      5'b11010:
        casez_tmp_19 = rob_bsy__26;
      5'b11011:
        casez_tmp_19 = rob_bsy__27;
      5'b11100:
        casez_tmp_19 = rob_bsy__28;
      5'b11101:
        casez_tmp_19 = rob_bsy__29;
      5'b11110:
        casez_tmp_19 = rob_bsy__30;
      default:
        casez_tmp_19 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1862 = _GEN_458 & ~casez_tmp_19;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_20 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_20 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_20 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_20 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_20 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_20 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_20 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_20 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_20 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_20 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_20 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_20 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_20 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_20 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_20 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_20 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_20 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_20 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_20 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_20 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_20 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_20 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_20 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_20 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_20 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_20 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_20 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_20 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_20 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_20 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_20 = rob_uop__30_ldst_val;
      default:
        casez_tmp_20 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_21 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_21 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_21 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_21 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_21 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_21 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_21 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_21 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_21 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_21 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_21 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_21 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_21 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_21 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_21 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_21 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_21 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_21 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_21 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_21 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_21 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_21 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_21 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_21 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_21 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_21 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_21 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_21 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_21 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_21 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_21 = rob_uop__30_pdst;
      default:
        casez_tmp_21 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1863 = _GEN_458 & casez_tmp_20 & casez_tmp_21 != io_wb_resps_2_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_22 = rob_val__0;
      5'b00001:
        casez_tmp_22 = rob_val__1;
      5'b00010:
        casez_tmp_22 = rob_val__2;
      5'b00011:
        casez_tmp_22 = rob_val__3;
      5'b00100:
        casez_tmp_22 = rob_val__4;
      5'b00101:
        casez_tmp_22 = rob_val__5;
      5'b00110:
        casez_tmp_22 = rob_val__6;
      5'b00111:
        casez_tmp_22 = rob_val__7;
      5'b01000:
        casez_tmp_22 = rob_val__8;
      5'b01001:
        casez_tmp_22 = rob_val__9;
      5'b01010:
        casez_tmp_22 = rob_val__10;
      5'b01011:
        casez_tmp_22 = rob_val__11;
      5'b01100:
        casez_tmp_22 = rob_val__12;
      5'b01101:
        casez_tmp_22 = rob_val__13;
      5'b01110:
        casez_tmp_22 = rob_val__14;
      5'b01111:
        casez_tmp_22 = rob_val__15;
      5'b10000:
        casez_tmp_22 = rob_val__16;
      5'b10001:
        casez_tmp_22 = rob_val__17;
      5'b10010:
        casez_tmp_22 = rob_val__18;
      5'b10011:
        casez_tmp_22 = rob_val__19;
      5'b10100:
        casez_tmp_22 = rob_val__20;
      5'b10101:
        casez_tmp_22 = rob_val__21;
      5'b10110:
        casez_tmp_22 = rob_val__22;
      5'b10111:
        casez_tmp_22 = rob_val__23;
      5'b11000:
        casez_tmp_22 = rob_val__24;
      5'b11001:
        casez_tmp_22 = rob_val__25;
      5'b11010:
        casez_tmp_22 = rob_val__26;
      5'b11011:
        casez_tmp_22 = rob_val__27;
      5'b11100:
        casez_tmp_22 = rob_val__28;
      5'b11101:
        casez_tmp_22 = rob_val__29;
      5'b11110:
        casez_tmp_22 = rob_val__30;
      default:
        casez_tmp_22 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1864 = _GEN_7 & ~casez_tmp_22;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_23 = rob_bsy__0;
      5'b00001:
        casez_tmp_23 = rob_bsy__1;
      5'b00010:
        casez_tmp_23 = rob_bsy__2;
      5'b00011:
        casez_tmp_23 = rob_bsy__3;
      5'b00100:
        casez_tmp_23 = rob_bsy__4;
      5'b00101:
        casez_tmp_23 = rob_bsy__5;
      5'b00110:
        casez_tmp_23 = rob_bsy__6;
      5'b00111:
        casez_tmp_23 = rob_bsy__7;
      5'b01000:
        casez_tmp_23 = rob_bsy__8;
      5'b01001:
        casez_tmp_23 = rob_bsy__9;
      5'b01010:
        casez_tmp_23 = rob_bsy__10;
      5'b01011:
        casez_tmp_23 = rob_bsy__11;
      5'b01100:
        casez_tmp_23 = rob_bsy__12;
      5'b01101:
        casez_tmp_23 = rob_bsy__13;
      5'b01110:
        casez_tmp_23 = rob_bsy__14;
      5'b01111:
        casez_tmp_23 = rob_bsy__15;
      5'b10000:
        casez_tmp_23 = rob_bsy__16;
      5'b10001:
        casez_tmp_23 = rob_bsy__17;
      5'b10010:
        casez_tmp_23 = rob_bsy__18;
      5'b10011:
        casez_tmp_23 = rob_bsy__19;
      5'b10100:
        casez_tmp_23 = rob_bsy__20;
      5'b10101:
        casez_tmp_23 = rob_bsy__21;
      5'b10110:
        casez_tmp_23 = rob_bsy__22;
      5'b10111:
        casez_tmp_23 = rob_bsy__23;
      5'b11000:
        casez_tmp_23 = rob_bsy__24;
      5'b11001:
        casez_tmp_23 = rob_bsy__25;
      5'b11010:
        casez_tmp_23 = rob_bsy__26;
      5'b11011:
        casez_tmp_23 = rob_bsy__27;
      5'b11100:
        casez_tmp_23 = rob_bsy__28;
      5'b11101:
        casez_tmp_23 = rob_bsy__29;
      5'b11110:
        casez_tmp_23 = rob_bsy__30;
      default:
        casez_tmp_23 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1865 = _GEN_7 & ~casez_tmp_23;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_24 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_24 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_24 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_24 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_24 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_24 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_24 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_24 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_24 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_24 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_24 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_24 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_24 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_24 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_24 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_24 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_24 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_24 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_24 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_24 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_24 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_24 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_24 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_24 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_24 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_24 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_24 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_24 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_24 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_24 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_24 = rob_uop__30_ldst_val;
      default:
        casez_tmp_24 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_25 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_25 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_25 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_25 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_25 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_25 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_25 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_25 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_25 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_25 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_25 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_25 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_25 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_25 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_25 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_25 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_25 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_25 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_25 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_25 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_25 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_25 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_25 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_25 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_25 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_25 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_25 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_25 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_25 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_25 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_25 = rob_uop__30_pdst;
      default:
        casez_tmp_25 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1866 = _GEN_7 & casez_tmp_24 & casez_tmp_25 != io_wb_resps_3_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_26 = rob_val__0;
      5'b00001:
        casez_tmp_26 = rob_val__1;
      5'b00010:
        casez_tmp_26 = rob_val__2;
      5'b00011:
        casez_tmp_26 = rob_val__3;
      5'b00100:
        casez_tmp_26 = rob_val__4;
      5'b00101:
        casez_tmp_26 = rob_val__5;
      5'b00110:
        casez_tmp_26 = rob_val__6;
      5'b00111:
        casez_tmp_26 = rob_val__7;
      5'b01000:
        casez_tmp_26 = rob_val__8;
      5'b01001:
        casez_tmp_26 = rob_val__9;
      5'b01010:
        casez_tmp_26 = rob_val__10;
      5'b01011:
        casez_tmp_26 = rob_val__11;
      5'b01100:
        casez_tmp_26 = rob_val__12;
      5'b01101:
        casez_tmp_26 = rob_val__13;
      5'b01110:
        casez_tmp_26 = rob_val__14;
      5'b01111:
        casez_tmp_26 = rob_val__15;
      5'b10000:
        casez_tmp_26 = rob_val__16;
      5'b10001:
        casez_tmp_26 = rob_val__17;
      5'b10010:
        casez_tmp_26 = rob_val__18;
      5'b10011:
        casez_tmp_26 = rob_val__19;
      5'b10100:
        casez_tmp_26 = rob_val__20;
      5'b10101:
        casez_tmp_26 = rob_val__21;
      5'b10110:
        casez_tmp_26 = rob_val__22;
      5'b10111:
        casez_tmp_26 = rob_val__23;
      5'b11000:
        casez_tmp_26 = rob_val__24;
      5'b11001:
        casez_tmp_26 = rob_val__25;
      5'b11010:
        casez_tmp_26 = rob_val__26;
      5'b11011:
        casez_tmp_26 = rob_val__27;
      5'b11100:
        casez_tmp_26 = rob_val__28;
      5'b11101:
        casez_tmp_26 = rob_val__29;
      5'b11110:
        casez_tmp_26 = rob_val__30;
      default:
        casez_tmp_26 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1867 = _GEN_459 & ~casez_tmp_26;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_27 = rob_bsy__0;
      5'b00001:
        casez_tmp_27 = rob_bsy__1;
      5'b00010:
        casez_tmp_27 = rob_bsy__2;
      5'b00011:
        casez_tmp_27 = rob_bsy__3;
      5'b00100:
        casez_tmp_27 = rob_bsy__4;
      5'b00101:
        casez_tmp_27 = rob_bsy__5;
      5'b00110:
        casez_tmp_27 = rob_bsy__6;
      5'b00111:
        casez_tmp_27 = rob_bsy__7;
      5'b01000:
        casez_tmp_27 = rob_bsy__8;
      5'b01001:
        casez_tmp_27 = rob_bsy__9;
      5'b01010:
        casez_tmp_27 = rob_bsy__10;
      5'b01011:
        casez_tmp_27 = rob_bsy__11;
      5'b01100:
        casez_tmp_27 = rob_bsy__12;
      5'b01101:
        casez_tmp_27 = rob_bsy__13;
      5'b01110:
        casez_tmp_27 = rob_bsy__14;
      5'b01111:
        casez_tmp_27 = rob_bsy__15;
      5'b10000:
        casez_tmp_27 = rob_bsy__16;
      5'b10001:
        casez_tmp_27 = rob_bsy__17;
      5'b10010:
        casez_tmp_27 = rob_bsy__18;
      5'b10011:
        casez_tmp_27 = rob_bsy__19;
      5'b10100:
        casez_tmp_27 = rob_bsy__20;
      5'b10101:
        casez_tmp_27 = rob_bsy__21;
      5'b10110:
        casez_tmp_27 = rob_bsy__22;
      5'b10111:
        casez_tmp_27 = rob_bsy__23;
      5'b11000:
        casez_tmp_27 = rob_bsy__24;
      5'b11001:
        casez_tmp_27 = rob_bsy__25;
      5'b11010:
        casez_tmp_27 = rob_bsy__26;
      5'b11011:
        casez_tmp_27 = rob_bsy__27;
      5'b11100:
        casez_tmp_27 = rob_bsy__28;
      5'b11101:
        casez_tmp_27 = rob_bsy__29;
      5'b11110:
        casez_tmp_27 = rob_bsy__30;
      default:
        casez_tmp_27 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1868 = _GEN_459 & ~casez_tmp_27;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_28 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_28 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_28 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_28 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_28 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_28 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_28 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_28 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_28 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_28 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_28 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_28 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_28 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_28 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_28 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_28 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_28 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_28 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_28 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_28 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_28 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_28 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_28 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_28 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_28 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_28 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_28 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_28 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_28 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_28 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_28 = rob_uop__30_ldst_val;
      default:
        casez_tmp_28 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_29 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_29 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_29 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_29 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_29 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_29 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_29 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_29 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_29 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_29 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_29 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_29 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_29 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_29 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_29 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_29 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_29 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_29 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_29 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_29 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_29 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_29 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_29 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_29 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_29 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_29 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_29 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_29 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_29 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_29 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_29 = rob_uop__30_pdst;
      default:
        casez_tmp_29 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1869 = _GEN_459 & casez_tmp_28 & casez_tmp_29 != io_wb_resps_4_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_30 = rob_val__0;
      5'b00001:
        casez_tmp_30 = rob_val__1;
      5'b00010:
        casez_tmp_30 = rob_val__2;
      5'b00011:
        casez_tmp_30 = rob_val__3;
      5'b00100:
        casez_tmp_30 = rob_val__4;
      5'b00101:
        casez_tmp_30 = rob_val__5;
      5'b00110:
        casez_tmp_30 = rob_val__6;
      5'b00111:
        casez_tmp_30 = rob_val__7;
      5'b01000:
        casez_tmp_30 = rob_val__8;
      5'b01001:
        casez_tmp_30 = rob_val__9;
      5'b01010:
        casez_tmp_30 = rob_val__10;
      5'b01011:
        casez_tmp_30 = rob_val__11;
      5'b01100:
        casez_tmp_30 = rob_val__12;
      5'b01101:
        casez_tmp_30 = rob_val__13;
      5'b01110:
        casez_tmp_30 = rob_val__14;
      5'b01111:
        casez_tmp_30 = rob_val__15;
      5'b10000:
        casez_tmp_30 = rob_val__16;
      5'b10001:
        casez_tmp_30 = rob_val__17;
      5'b10010:
        casez_tmp_30 = rob_val__18;
      5'b10011:
        casez_tmp_30 = rob_val__19;
      5'b10100:
        casez_tmp_30 = rob_val__20;
      5'b10101:
        casez_tmp_30 = rob_val__21;
      5'b10110:
        casez_tmp_30 = rob_val__22;
      5'b10111:
        casez_tmp_30 = rob_val__23;
      5'b11000:
        casez_tmp_30 = rob_val__24;
      5'b11001:
        casez_tmp_30 = rob_val__25;
      5'b11010:
        casez_tmp_30 = rob_val__26;
      5'b11011:
        casez_tmp_30 = rob_val__27;
      5'b11100:
        casez_tmp_30 = rob_val__28;
      5'b11101:
        casez_tmp_30 = rob_val__29;
      5'b11110:
        casez_tmp_30 = rob_val__30;
      default:
        casez_tmp_30 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1870 = _GEN_6 & ~casez_tmp_30;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_31 = rob_bsy__0;
      5'b00001:
        casez_tmp_31 = rob_bsy__1;
      5'b00010:
        casez_tmp_31 = rob_bsy__2;
      5'b00011:
        casez_tmp_31 = rob_bsy__3;
      5'b00100:
        casez_tmp_31 = rob_bsy__4;
      5'b00101:
        casez_tmp_31 = rob_bsy__5;
      5'b00110:
        casez_tmp_31 = rob_bsy__6;
      5'b00111:
        casez_tmp_31 = rob_bsy__7;
      5'b01000:
        casez_tmp_31 = rob_bsy__8;
      5'b01001:
        casez_tmp_31 = rob_bsy__9;
      5'b01010:
        casez_tmp_31 = rob_bsy__10;
      5'b01011:
        casez_tmp_31 = rob_bsy__11;
      5'b01100:
        casez_tmp_31 = rob_bsy__12;
      5'b01101:
        casez_tmp_31 = rob_bsy__13;
      5'b01110:
        casez_tmp_31 = rob_bsy__14;
      5'b01111:
        casez_tmp_31 = rob_bsy__15;
      5'b10000:
        casez_tmp_31 = rob_bsy__16;
      5'b10001:
        casez_tmp_31 = rob_bsy__17;
      5'b10010:
        casez_tmp_31 = rob_bsy__18;
      5'b10011:
        casez_tmp_31 = rob_bsy__19;
      5'b10100:
        casez_tmp_31 = rob_bsy__20;
      5'b10101:
        casez_tmp_31 = rob_bsy__21;
      5'b10110:
        casez_tmp_31 = rob_bsy__22;
      5'b10111:
        casez_tmp_31 = rob_bsy__23;
      5'b11000:
        casez_tmp_31 = rob_bsy__24;
      5'b11001:
        casez_tmp_31 = rob_bsy__25;
      5'b11010:
        casez_tmp_31 = rob_bsy__26;
      5'b11011:
        casez_tmp_31 = rob_bsy__27;
      5'b11100:
        casez_tmp_31 = rob_bsy__28;
      5'b11101:
        casez_tmp_31 = rob_bsy__29;
      5'b11110:
        casez_tmp_31 = rob_bsy__30;
      default:
        casez_tmp_31 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1871 = _GEN_6 & ~casez_tmp_31;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_32 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_32 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_32 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_32 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_32 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_32 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_32 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_32 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_32 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_32 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_32 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_32 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_32 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_32 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_32 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_32 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_32 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_32 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_32 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_32 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_32 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_32 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_32 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_32 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_32 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_32 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_32 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_32 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_32 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_32 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_32 = rob_uop__30_ldst_val;
      default:
        casez_tmp_32 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_33 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_33 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_33 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_33 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_33 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_33 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_33 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_33 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_33 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_33 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_33 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_33 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_33 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_33 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_33 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_33 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_33 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_33 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_33 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_33 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_33 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_33 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_33 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_33 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_33 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_33 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_33 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_33 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_33 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_33 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_33 = rob_uop__30_pdst;
      default:
        casez_tmp_33 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1872 = _GEN_6 & casez_tmp_32 & casez_tmp_33 != io_wb_resps_5_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_34 = rob_val__0;
      5'b00001:
        casez_tmp_34 = rob_val__1;
      5'b00010:
        casez_tmp_34 = rob_val__2;
      5'b00011:
        casez_tmp_34 = rob_val__3;
      5'b00100:
        casez_tmp_34 = rob_val__4;
      5'b00101:
        casez_tmp_34 = rob_val__5;
      5'b00110:
        casez_tmp_34 = rob_val__6;
      5'b00111:
        casez_tmp_34 = rob_val__7;
      5'b01000:
        casez_tmp_34 = rob_val__8;
      5'b01001:
        casez_tmp_34 = rob_val__9;
      5'b01010:
        casez_tmp_34 = rob_val__10;
      5'b01011:
        casez_tmp_34 = rob_val__11;
      5'b01100:
        casez_tmp_34 = rob_val__12;
      5'b01101:
        casez_tmp_34 = rob_val__13;
      5'b01110:
        casez_tmp_34 = rob_val__14;
      5'b01111:
        casez_tmp_34 = rob_val__15;
      5'b10000:
        casez_tmp_34 = rob_val__16;
      5'b10001:
        casez_tmp_34 = rob_val__17;
      5'b10010:
        casez_tmp_34 = rob_val__18;
      5'b10011:
        casez_tmp_34 = rob_val__19;
      5'b10100:
        casez_tmp_34 = rob_val__20;
      5'b10101:
        casez_tmp_34 = rob_val__21;
      5'b10110:
        casez_tmp_34 = rob_val__22;
      5'b10111:
        casez_tmp_34 = rob_val__23;
      5'b11000:
        casez_tmp_34 = rob_val__24;
      5'b11001:
        casez_tmp_34 = rob_val__25;
      5'b11010:
        casez_tmp_34 = rob_val__26;
      5'b11011:
        casez_tmp_34 = rob_val__27;
      5'b11100:
        casez_tmp_34 = rob_val__28;
      5'b11101:
        casez_tmp_34 = rob_val__29;
      5'b11110:
        casez_tmp_34 = rob_val__30;
      default:
        casez_tmp_34 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1873 = _GEN_460 & ~casez_tmp_34;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_35 = rob_bsy__0;
      5'b00001:
        casez_tmp_35 = rob_bsy__1;
      5'b00010:
        casez_tmp_35 = rob_bsy__2;
      5'b00011:
        casez_tmp_35 = rob_bsy__3;
      5'b00100:
        casez_tmp_35 = rob_bsy__4;
      5'b00101:
        casez_tmp_35 = rob_bsy__5;
      5'b00110:
        casez_tmp_35 = rob_bsy__6;
      5'b00111:
        casez_tmp_35 = rob_bsy__7;
      5'b01000:
        casez_tmp_35 = rob_bsy__8;
      5'b01001:
        casez_tmp_35 = rob_bsy__9;
      5'b01010:
        casez_tmp_35 = rob_bsy__10;
      5'b01011:
        casez_tmp_35 = rob_bsy__11;
      5'b01100:
        casez_tmp_35 = rob_bsy__12;
      5'b01101:
        casez_tmp_35 = rob_bsy__13;
      5'b01110:
        casez_tmp_35 = rob_bsy__14;
      5'b01111:
        casez_tmp_35 = rob_bsy__15;
      5'b10000:
        casez_tmp_35 = rob_bsy__16;
      5'b10001:
        casez_tmp_35 = rob_bsy__17;
      5'b10010:
        casez_tmp_35 = rob_bsy__18;
      5'b10011:
        casez_tmp_35 = rob_bsy__19;
      5'b10100:
        casez_tmp_35 = rob_bsy__20;
      5'b10101:
        casez_tmp_35 = rob_bsy__21;
      5'b10110:
        casez_tmp_35 = rob_bsy__22;
      5'b10111:
        casez_tmp_35 = rob_bsy__23;
      5'b11000:
        casez_tmp_35 = rob_bsy__24;
      5'b11001:
        casez_tmp_35 = rob_bsy__25;
      5'b11010:
        casez_tmp_35 = rob_bsy__26;
      5'b11011:
        casez_tmp_35 = rob_bsy__27;
      5'b11100:
        casez_tmp_35 = rob_bsy__28;
      5'b11101:
        casez_tmp_35 = rob_bsy__29;
      5'b11110:
        casez_tmp_35 = rob_bsy__30;
      default:
        casez_tmp_35 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1874 = _GEN_460 & ~casez_tmp_35;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_36 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_36 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_36 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_36 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_36 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_36 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_36 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_36 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_36 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_36 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_36 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_36 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_36 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_36 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_36 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_36 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_36 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_36 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_36 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_36 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_36 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_36 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_36 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_36 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_36 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_36 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_36 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_36 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_36 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_36 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_36 = rob_uop__30_ldst_val;
      default:
        casez_tmp_36 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_37 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_37 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_37 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_37 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_37 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_37 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_37 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_37 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_37 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_37 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_37 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_37 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_37 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_37 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_37 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_37 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_37 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_37 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_37 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_37 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_37 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_37 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_37 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_37 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_37 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_37 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_37 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_37 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_37 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_37 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_37 = rob_uop__30_pdst;
      default:
        casez_tmp_37 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1875 = _GEN_460 & casez_tmp_36 & casez_tmp_37 != io_wb_resps_6_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_38 = rob_val__0;
      5'b00001:
        casez_tmp_38 = rob_val__1;
      5'b00010:
        casez_tmp_38 = rob_val__2;
      5'b00011:
        casez_tmp_38 = rob_val__3;
      5'b00100:
        casez_tmp_38 = rob_val__4;
      5'b00101:
        casez_tmp_38 = rob_val__5;
      5'b00110:
        casez_tmp_38 = rob_val__6;
      5'b00111:
        casez_tmp_38 = rob_val__7;
      5'b01000:
        casez_tmp_38 = rob_val__8;
      5'b01001:
        casez_tmp_38 = rob_val__9;
      5'b01010:
        casez_tmp_38 = rob_val__10;
      5'b01011:
        casez_tmp_38 = rob_val__11;
      5'b01100:
        casez_tmp_38 = rob_val__12;
      5'b01101:
        casez_tmp_38 = rob_val__13;
      5'b01110:
        casez_tmp_38 = rob_val__14;
      5'b01111:
        casez_tmp_38 = rob_val__15;
      5'b10000:
        casez_tmp_38 = rob_val__16;
      5'b10001:
        casez_tmp_38 = rob_val__17;
      5'b10010:
        casez_tmp_38 = rob_val__18;
      5'b10011:
        casez_tmp_38 = rob_val__19;
      5'b10100:
        casez_tmp_38 = rob_val__20;
      5'b10101:
        casez_tmp_38 = rob_val__21;
      5'b10110:
        casez_tmp_38 = rob_val__22;
      5'b10111:
        casez_tmp_38 = rob_val__23;
      5'b11000:
        casez_tmp_38 = rob_val__24;
      5'b11001:
        casez_tmp_38 = rob_val__25;
      5'b11010:
        casez_tmp_38 = rob_val__26;
      5'b11011:
        casez_tmp_38 = rob_val__27;
      5'b11100:
        casez_tmp_38 = rob_val__28;
      5'b11101:
        casez_tmp_38 = rob_val__29;
      5'b11110:
        casez_tmp_38 = rob_val__30;
      default:
        casez_tmp_38 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1876 = _GEN_5 & ~casez_tmp_38;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_39 = rob_bsy__0;
      5'b00001:
        casez_tmp_39 = rob_bsy__1;
      5'b00010:
        casez_tmp_39 = rob_bsy__2;
      5'b00011:
        casez_tmp_39 = rob_bsy__3;
      5'b00100:
        casez_tmp_39 = rob_bsy__4;
      5'b00101:
        casez_tmp_39 = rob_bsy__5;
      5'b00110:
        casez_tmp_39 = rob_bsy__6;
      5'b00111:
        casez_tmp_39 = rob_bsy__7;
      5'b01000:
        casez_tmp_39 = rob_bsy__8;
      5'b01001:
        casez_tmp_39 = rob_bsy__9;
      5'b01010:
        casez_tmp_39 = rob_bsy__10;
      5'b01011:
        casez_tmp_39 = rob_bsy__11;
      5'b01100:
        casez_tmp_39 = rob_bsy__12;
      5'b01101:
        casez_tmp_39 = rob_bsy__13;
      5'b01110:
        casez_tmp_39 = rob_bsy__14;
      5'b01111:
        casez_tmp_39 = rob_bsy__15;
      5'b10000:
        casez_tmp_39 = rob_bsy__16;
      5'b10001:
        casez_tmp_39 = rob_bsy__17;
      5'b10010:
        casez_tmp_39 = rob_bsy__18;
      5'b10011:
        casez_tmp_39 = rob_bsy__19;
      5'b10100:
        casez_tmp_39 = rob_bsy__20;
      5'b10101:
        casez_tmp_39 = rob_bsy__21;
      5'b10110:
        casez_tmp_39 = rob_bsy__22;
      5'b10111:
        casez_tmp_39 = rob_bsy__23;
      5'b11000:
        casez_tmp_39 = rob_bsy__24;
      5'b11001:
        casez_tmp_39 = rob_bsy__25;
      5'b11010:
        casez_tmp_39 = rob_bsy__26;
      5'b11011:
        casez_tmp_39 = rob_bsy__27;
      5'b11100:
        casez_tmp_39 = rob_bsy__28;
      5'b11101:
        casez_tmp_39 = rob_bsy__29;
      5'b11110:
        casez_tmp_39 = rob_bsy__30;
      default:
        casez_tmp_39 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1877 = _GEN_5 & ~casez_tmp_39;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_40 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_40 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_40 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_40 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_40 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_40 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_40 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_40 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_40 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_40 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_40 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_40 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_40 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_40 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_40 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_40 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_40 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_40 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_40 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_40 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_40 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_40 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_40 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_40 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_40 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_40 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_40 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_40 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_40 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_40 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_40 = rob_uop__30_ldst_val;
      default:
        casez_tmp_40 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_41 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_41 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_41 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_41 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_41 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_41 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_41 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_41 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_41 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_41 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_41 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_41 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_41 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_41 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_41 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_41 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_41 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_41 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_41 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_41 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_41 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_41 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_41 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_41 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_41 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_41 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_41 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_41 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_41 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_41 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_41 = rob_uop__30_pdst;
      default:
        casez_tmp_41 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1878 = _GEN_5 & casez_tmp_40 & casez_tmp_41 != io_wb_resps_7_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_42 = rob_val__0;
      5'b00001:
        casez_tmp_42 = rob_val__1;
      5'b00010:
        casez_tmp_42 = rob_val__2;
      5'b00011:
        casez_tmp_42 = rob_val__3;
      5'b00100:
        casez_tmp_42 = rob_val__4;
      5'b00101:
        casez_tmp_42 = rob_val__5;
      5'b00110:
        casez_tmp_42 = rob_val__6;
      5'b00111:
        casez_tmp_42 = rob_val__7;
      5'b01000:
        casez_tmp_42 = rob_val__8;
      5'b01001:
        casez_tmp_42 = rob_val__9;
      5'b01010:
        casez_tmp_42 = rob_val__10;
      5'b01011:
        casez_tmp_42 = rob_val__11;
      5'b01100:
        casez_tmp_42 = rob_val__12;
      5'b01101:
        casez_tmp_42 = rob_val__13;
      5'b01110:
        casez_tmp_42 = rob_val__14;
      5'b01111:
        casez_tmp_42 = rob_val__15;
      5'b10000:
        casez_tmp_42 = rob_val__16;
      5'b10001:
        casez_tmp_42 = rob_val__17;
      5'b10010:
        casez_tmp_42 = rob_val__18;
      5'b10011:
        casez_tmp_42 = rob_val__19;
      5'b10100:
        casez_tmp_42 = rob_val__20;
      5'b10101:
        casez_tmp_42 = rob_val__21;
      5'b10110:
        casez_tmp_42 = rob_val__22;
      5'b10111:
        casez_tmp_42 = rob_val__23;
      5'b11000:
        casez_tmp_42 = rob_val__24;
      5'b11001:
        casez_tmp_42 = rob_val__25;
      5'b11010:
        casez_tmp_42 = rob_val__26;
      5'b11011:
        casez_tmp_42 = rob_val__27;
      5'b11100:
        casez_tmp_42 = rob_val__28;
      5'b11101:
        casez_tmp_42 = rob_val__29;
      5'b11110:
        casez_tmp_42 = rob_val__30;
      default:
        casez_tmp_42 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1879 = _GEN_461 & ~casez_tmp_42;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_43 = rob_bsy__0;
      5'b00001:
        casez_tmp_43 = rob_bsy__1;
      5'b00010:
        casez_tmp_43 = rob_bsy__2;
      5'b00011:
        casez_tmp_43 = rob_bsy__3;
      5'b00100:
        casez_tmp_43 = rob_bsy__4;
      5'b00101:
        casez_tmp_43 = rob_bsy__5;
      5'b00110:
        casez_tmp_43 = rob_bsy__6;
      5'b00111:
        casez_tmp_43 = rob_bsy__7;
      5'b01000:
        casez_tmp_43 = rob_bsy__8;
      5'b01001:
        casez_tmp_43 = rob_bsy__9;
      5'b01010:
        casez_tmp_43 = rob_bsy__10;
      5'b01011:
        casez_tmp_43 = rob_bsy__11;
      5'b01100:
        casez_tmp_43 = rob_bsy__12;
      5'b01101:
        casez_tmp_43 = rob_bsy__13;
      5'b01110:
        casez_tmp_43 = rob_bsy__14;
      5'b01111:
        casez_tmp_43 = rob_bsy__15;
      5'b10000:
        casez_tmp_43 = rob_bsy__16;
      5'b10001:
        casez_tmp_43 = rob_bsy__17;
      5'b10010:
        casez_tmp_43 = rob_bsy__18;
      5'b10011:
        casez_tmp_43 = rob_bsy__19;
      5'b10100:
        casez_tmp_43 = rob_bsy__20;
      5'b10101:
        casez_tmp_43 = rob_bsy__21;
      5'b10110:
        casez_tmp_43 = rob_bsy__22;
      5'b10111:
        casez_tmp_43 = rob_bsy__23;
      5'b11000:
        casez_tmp_43 = rob_bsy__24;
      5'b11001:
        casez_tmp_43 = rob_bsy__25;
      5'b11010:
        casez_tmp_43 = rob_bsy__26;
      5'b11011:
        casez_tmp_43 = rob_bsy__27;
      5'b11100:
        casez_tmp_43 = rob_bsy__28;
      5'b11101:
        casez_tmp_43 = rob_bsy__29;
      5'b11110:
        casez_tmp_43 = rob_bsy__30;
      default:
        casez_tmp_43 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1880 = _GEN_461 & ~casez_tmp_43;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_44 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_44 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_44 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_44 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_44 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_44 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_44 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_44 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_44 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_44 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_44 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_44 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_44 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_44 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_44 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_44 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_44 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_44 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_44 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_44 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_44 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_44 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_44 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_44 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_44 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_44 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_44 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_44 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_44 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_44 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_44 = rob_uop__30_ldst_val;
      default:
        casez_tmp_44 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_45 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_45 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_45 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_45 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_45 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_45 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_45 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_45 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_45 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_45 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_45 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_45 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_45 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_45 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_45 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_45 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_45 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_45 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_45 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_45 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_45 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_45 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_45 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_45 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_45 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_45 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_45 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_45 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_45 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_45 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_45 = rob_uop__30_pdst;
      default:
        casez_tmp_45 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1881 = _GEN_461 & casez_tmp_44 & casez_tmp_45 != io_wb_resps_8_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_46 = rob_val__0;
      5'b00001:
        casez_tmp_46 = rob_val__1;
      5'b00010:
        casez_tmp_46 = rob_val__2;
      5'b00011:
        casez_tmp_46 = rob_val__3;
      5'b00100:
        casez_tmp_46 = rob_val__4;
      5'b00101:
        casez_tmp_46 = rob_val__5;
      5'b00110:
        casez_tmp_46 = rob_val__6;
      5'b00111:
        casez_tmp_46 = rob_val__7;
      5'b01000:
        casez_tmp_46 = rob_val__8;
      5'b01001:
        casez_tmp_46 = rob_val__9;
      5'b01010:
        casez_tmp_46 = rob_val__10;
      5'b01011:
        casez_tmp_46 = rob_val__11;
      5'b01100:
        casez_tmp_46 = rob_val__12;
      5'b01101:
        casez_tmp_46 = rob_val__13;
      5'b01110:
        casez_tmp_46 = rob_val__14;
      5'b01111:
        casez_tmp_46 = rob_val__15;
      5'b10000:
        casez_tmp_46 = rob_val__16;
      5'b10001:
        casez_tmp_46 = rob_val__17;
      5'b10010:
        casez_tmp_46 = rob_val__18;
      5'b10011:
        casez_tmp_46 = rob_val__19;
      5'b10100:
        casez_tmp_46 = rob_val__20;
      5'b10101:
        casez_tmp_46 = rob_val__21;
      5'b10110:
        casez_tmp_46 = rob_val__22;
      5'b10111:
        casez_tmp_46 = rob_val__23;
      5'b11000:
        casez_tmp_46 = rob_val__24;
      5'b11001:
        casez_tmp_46 = rob_val__25;
      5'b11010:
        casez_tmp_46 = rob_val__26;
      5'b11011:
        casez_tmp_46 = rob_val__27;
      5'b11100:
        casez_tmp_46 = rob_val__28;
      5'b11101:
        casez_tmp_46 = rob_val__29;
      5'b11110:
        casez_tmp_46 = rob_val__30;
      default:
        casez_tmp_46 = rob_val__31;
    endcase
  end // always @(*)
  wire       _GEN_1882 = _GEN_4 & ~casez_tmp_46;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_47 = rob_bsy__0;
      5'b00001:
        casez_tmp_47 = rob_bsy__1;
      5'b00010:
        casez_tmp_47 = rob_bsy__2;
      5'b00011:
        casez_tmp_47 = rob_bsy__3;
      5'b00100:
        casez_tmp_47 = rob_bsy__4;
      5'b00101:
        casez_tmp_47 = rob_bsy__5;
      5'b00110:
        casez_tmp_47 = rob_bsy__6;
      5'b00111:
        casez_tmp_47 = rob_bsy__7;
      5'b01000:
        casez_tmp_47 = rob_bsy__8;
      5'b01001:
        casez_tmp_47 = rob_bsy__9;
      5'b01010:
        casez_tmp_47 = rob_bsy__10;
      5'b01011:
        casez_tmp_47 = rob_bsy__11;
      5'b01100:
        casez_tmp_47 = rob_bsy__12;
      5'b01101:
        casez_tmp_47 = rob_bsy__13;
      5'b01110:
        casez_tmp_47 = rob_bsy__14;
      5'b01111:
        casez_tmp_47 = rob_bsy__15;
      5'b10000:
        casez_tmp_47 = rob_bsy__16;
      5'b10001:
        casez_tmp_47 = rob_bsy__17;
      5'b10010:
        casez_tmp_47 = rob_bsy__18;
      5'b10011:
        casez_tmp_47 = rob_bsy__19;
      5'b10100:
        casez_tmp_47 = rob_bsy__20;
      5'b10101:
        casez_tmp_47 = rob_bsy__21;
      5'b10110:
        casez_tmp_47 = rob_bsy__22;
      5'b10111:
        casez_tmp_47 = rob_bsy__23;
      5'b11000:
        casez_tmp_47 = rob_bsy__24;
      5'b11001:
        casez_tmp_47 = rob_bsy__25;
      5'b11010:
        casez_tmp_47 = rob_bsy__26;
      5'b11011:
        casez_tmp_47 = rob_bsy__27;
      5'b11100:
        casez_tmp_47 = rob_bsy__28;
      5'b11101:
        casez_tmp_47 = rob_bsy__29;
      5'b11110:
        casez_tmp_47 = rob_bsy__30;
      default:
        casez_tmp_47 = rob_bsy__31;
    endcase
  end // always @(*)
  wire       _GEN_1883 = _GEN_4 & ~casez_tmp_47;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_48 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_48 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_48 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_48 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_48 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_48 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_48 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_48 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_48 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_48 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_48 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_48 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_48 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_48 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_48 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_48 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_48 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_48 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_48 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_48 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_48 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_48 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_48 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_48 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_48 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_48 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_48 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_48 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_48 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_48 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_48 = rob_uop__30_ldst_val;
      default:
        casez_tmp_48 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_49 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_49 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_49 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_49 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_49 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_49 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_49 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_49 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_49 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_49 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_49 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_49 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_49 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_49 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_49 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_49 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_49 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_49 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_49 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_49 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_49 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_49 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_49 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_49 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_49 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_49 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_49 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_49 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_49 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_49 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_49 = rob_uop__30_pdst;
      default:
        casez_tmp_49 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1884 = _GEN_4 & casez_tmp_48 & casez_tmp_49 != io_wb_resps_9_bits_uop_pdst;
  reg        rob_unsafe_1_0;
  reg        rob_unsafe_1_1;
  reg        rob_unsafe_1_2;
  reg        rob_unsafe_1_3;
  reg        rob_unsafe_1_4;
  reg        rob_unsafe_1_5;
  reg        rob_unsafe_1_6;
  reg        rob_unsafe_1_7;
  reg        rob_unsafe_1_8;
  reg        rob_unsafe_1_9;
  reg        rob_unsafe_1_10;
  reg        rob_unsafe_1_11;
  reg        rob_unsafe_1_12;
  reg        rob_unsafe_1_13;
  reg        rob_unsafe_1_14;
  reg        rob_unsafe_1_15;
  reg        rob_unsafe_1_16;
  reg        rob_unsafe_1_17;
  reg        rob_unsafe_1_18;
  reg        rob_unsafe_1_19;
  reg        rob_unsafe_1_20;
  reg        rob_unsafe_1_21;
  reg        rob_unsafe_1_22;
  reg        rob_unsafe_1_23;
  reg        rob_unsafe_1_24;
  reg        rob_unsafe_1_25;
  reg        rob_unsafe_1_26;
  reg        rob_unsafe_1_27;
  reg        rob_unsafe_1_28;
  reg        rob_unsafe_1_29;
  reg        rob_unsafe_1_30;
  reg        rob_unsafe_1_31;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp_50 = rob_val_1_0;
      5'b00001:
        casez_tmp_50 = rob_val_1_1;
      5'b00010:
        casez_tmp_50 = rob_val_1_2;
      5'b00011:
        casez_tmp_50 = rob_val_1_3;
      5'b00100:
        casez_tmp_50 = rob_val_1_4;
      5'b00101:
        casez_tmp_50 = rob_val_1_5;
      5'b00110:
        casez_tmp_50 = rob_val_1_6;
      5'b00111:
        casez_tmp_50 = rob_val_1_7;
      5'b01000:
        casez_tmp_50 = rob_val_1_8;
      5'b01001:
        casez_tmp_50 = rob_val_1_9;
      5'b01010:
        casez_tmp_50 = rob_val_1_10;
      5'b01011:
        casez_tmp_50 = rob_val_1_11;
      5'b01100:
        casez_tmp_50 = rob_val_1_12;
      5'b01101:
        casez_tmp_50 = rob_val_1_13;
      5'b01110:
        casez_tmp_50 = rob_val_1_14;
      5'b01111:
        casez_tmp_50 = rob_val_1_15;
      5'b10000:
        casez_tmp_50 = rob_val_1_16;
      5'b10001:
        casez_tmp_50 = rob_val_1_17;
      5'b10010:
        casez_tmp_50 = rob_val_1_18;
      5'b10011:
        casez_tmp_50 = rob_val_1_19;
      5'b10100:
        casez_tmp_50 = rob_val_1_20;
      5'b10101:
        casez_tmp_50 = rob_val_1_21;
      5'b10110:
        casez_tmp_50 = rob_val_1_22;
      5'b10111:
        casez_tmp_50 = rob_val_1_23;
      5'b11000:
        casez_tmp_50 = rob_val_1_24;
      5'b11001:
        casez_tmp_50 = rob_val_1_25;
      5'b11010:
        casez_tmp_50 = rob_val_1_26;
      5'b11011:
        casez_tmp_50 = rob_val_1_27;
      5'b11100:
        casez_tmp_50 = rob_val_1_28;
      5'b11101:
        casez_tmp_50 = rob_val_1_29;
      5'b11110:
        casez_tmp_50 = rob_val_1_30;
      default:
        casez_tmp_50 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1885 = io_enq_uops_1_rob_idx[6:2] == rob_tail;
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_51 = rob_val_1_0;
      5'b00001:
        casez_tmp_51 = rob_val_1_1;
      5'b00010:
        casez_tmp_51 = rob_val_1_2;
      5'b00011:
        casez_tmp_51 = rob_val_1_3;
      5'b00100:
        casez_tmp_51 = rob_val_1_4;
      5'b00101:
        casez_tmp_51 = rob_val_1_5;
      5'b00110:
        casez_tmp_51 = rob_val_1_6;
      5'b00111:
        casez_tmp_51 = rob_val_1_7;
      5'b01000:
        casez_tmp_51 = rob_val_1_8;
      5'b01001:
        casez_tmp_51 = rob_val_1_9;
      5'b01010:
        casez_tmp_51 = rob_val_1_10;
      5'b01011:
        casez_tmp_51 = rob_val_1_11;
      5'b01100:
        casez_tmp_51 = rob_val_1_12;
      5'b01101:
        casez_tmp_51 = rob_val_1_13;
      5'b01110:
        casez_tmp_51 = rob_val_1_14;
      5'b01111:
        casez_tmp_51 = rob_val_1_15;
      5'b10000:
        casez_tmp_51 = rob_val_1_16;
      5'b10001:
        casez_tmp_51 = rob_val_1_17;
      5'b10010:
        casez_tmp_51 = rob_val_1_18;
      5'b10011:
        casez_tmp_51 = rob_val_1_19;
      5'b10100:
        casez_tmp_51 = rob_val_1_20;
      5'b10101:
        casez_tmp_51 = rob_val_1_21;
      5'b10110:
        casez_tmp_51 = rob_val_1_22;
      5'b10111:
        casez_tmp_51 = rob_val_1_23;
      5'b11000:
        casez_tmp_51 = rob_val_1_24;
      5'b11001:
        casez_tmp_51 = rob_val_1_25;
      5'b11010:
        casez_tmp_51 = rob_val_1_26;
      5'b11011:
        casez_tmp_51 = rob_val_1_27;
      5'b11100:
        casez_tmp_51 = rob_val_1_28;
      5'b11101:
        casez_tmp_51 = rob_val_1_29;
      5'b11110:
        casez_tmp_51 = rob_val_1_30;
      default:
        casez_tmp_51 = rob_val_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_52 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_52 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_52 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_52 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_52 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_52 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_52 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_52 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_52 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_52 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_52 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_52 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_52 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_52 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_52 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_52 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_52 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_52 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_52 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_52 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_52 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_52 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_52 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_52 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_52 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_52 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_52 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_52 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_52 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_52 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_52 = rob_bsy_1_30;
      default:
        casez_tmp_52 = rob_bsy_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_53 = rob_val_1_0;
      5'b00001:
        casez_tmp_53 = rob_val_1_1;
      5'b00010:
        casez_tmp_53 = rob_val_1_2;
      5'b00011:
        casez_tmp_53 = rob_val_1_3;
      5'b00100:
        casez_tmp_53 = rob_val_1_4;
      5'b00101:
        casez_tmp_53 = rob_val_1_5;
      5'b00110:
        casez_tmp_53 = rob_val_1_6;
      5'b00111:
        casez_tmp_53 = rob_val_1_7;
      5'b01000:
        casez_tmp_53 = rob_val_1_8;
      5'b01001:
        casez_tmp_53 = rob_val_1_9;
      5'b01010:
        casez_tmp_53 = rob_val_1_10;
      5'b01011:
        casez_tmp_53 = rob_val_1_11;
      5'b01100:
        casez_tmp_53 = rob_val_1_12;
      5'b01101:
        casez_tmp_53 = rob_val_1_13;
      5'b01110:
        casez_tmp_53 = rob_val_1_14;
      5'b01111:
        casez_tmp_53 = rob_val_1_15;
      5'b10000:
        casez_tmp_53 = rob_val_1_16;
      5'b10001:
        casez_tmp_53 = rob_val_1_17;
      5'b10010:
        casez_tmp_53 = rob_val_1_18;
      5'b10011:
        casez_tmp_53 = rob_val_1_19;
      5'b10100:
        casez_tmp_53 = rob_val_1_20;
      5'b10101:
        casez_tmp_53 = rob_val_1_21;
      5'b10110:
        casez_tmp_53 = rob_val_1_22;
      5'b10111:
        casez_tmp_53 = rob_val_1_23;
      5'b11000:
        casez_tmp_53 = rob_val_1_24;
      5'b11001:
        casez_tmp_53 = rob_val_1_25;
      5'b11010:
        casez_tmp_53 = rob_val_1_26;
      5'b11011:
        casez_tmp_53 = rob_val_1_27;
      5'b11100:
        casez_tmp_53 = rob_val_1_28;
      5'b11101:
        casez_tmp_53 = rob_val_1_29;
      5'b11110:
        casez_tmp_53 = rob_val_1_30;
      default:
        casez_tmp_53 = rob_val_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_54 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_54 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_54 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_54 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_54 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_54 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_54 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_54 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_54 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_54 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_54 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_54 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_54 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_54 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_54 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_54 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_54 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_54 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_54 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_54 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_54 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_54 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_54 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_54 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_54 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_54 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_54 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_54 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_54 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_54 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_54 = rob_bsy_1_30;
      default:
        casez_tmp_54 = rob_bsy_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_55 = rob_val_1_0;
      5'b00001:
        casez_tmp_55 = rob_val_1_1;
      5'b00010:
        casez_tmp_55 = rob_val_1_2;
      5'b00011:
        casez_tmp_55 = rob_val_1_3;
      5'b00100:
        casez_tmp_55 = rob_val_1_4;
      5'b00101:
        casez_tmp_55 = rob_val_1_5;
      5'b00110:
        casez_tmp_55 = rob_val_1_6;
      5'b00111:
        casez_tmp_55 = rob_val_1_7;
      5'b01000:
        casez_tmp_55 = rob_val_1_8;
      5'b01001:
        casez_tmp_55 = rob_val_1_9;
      5'b01010:
        casez_tmp_55 = rob_val_1_10;
      5'b01011:
        casez_tmp_55 = rob_val_1_11;
      5'b01100:
        casez_tmp_55 = rob_val_1_12;
      5'b01101:
        casez_tmp_55 = rob_val_1_13;
      5'b01110:
        casez_tmp_55 = rob_val_1_14;
      5'b01111:
        casez_tmp_55 = rob_val_1_15;
      5'b10000:
        casez_tmp_55 = rob_val_1_16;
      5'b10001:
        casez_tmp_55 = rob_val_1_17;
      5'b10010:
        casez_tmp_55 = rob_val_1_18;
      5'b10011:
        casez_tmp_55 = rob_val_1_19;
      5'b10100:
        casez_tmp_55 = rob_val_1_20;
      5'b10101:
        casez_tmp_55 = rob_val_1_21;
      5'b10110:
        casez_tmp_55 = rob_val_1_22;
      5'b10111:
        casez_tmp_55 = rob_val_1_23;
      5'b11000:
        casez_tmp_55 = rob_val_1_24;
      5'b11001:
        casez_tmp_55 = rob_val_1_25;
      5'b11010:
        casez_tmp_55 = rob_val_1_26;
      5'b11011:
        casez_tmp_55 = rob_val_1_27;
      5'b11100:
        casez_tmp_55 = rob_val_1_28;
      5'b11101:
        casez_tmp_55 = rob_val_1_29;
      5'b11110:
        casez_tmp_55 = rob_val_1_30;
      default:
        casez_tmp_55 = rob_val_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_56 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_56 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_56 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_56 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_56 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_56 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_56 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_56 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_56 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_56 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_56 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_56 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_56 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_56 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_56 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_56 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_56 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_56 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_56 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_56 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_56 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_56 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_56 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_56 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_56 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_56 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_56 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_56 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_56 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_56 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_56 = rob_bsy_1_30;
      default:
        casez_tmp_56 = rob_bsy_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_2)
      5'b00000:
        casez_tmp_57 = rob_unsafe_1_0;
      5'b00001:
        casez_tmp_57 = rob_unsafe_1_1;
      5'b00010:
        casez_tmp_57 = rob_unsafe_1_2;
      5'b00011:
        casez_tmp_57 = rob_unsafe_1_3;
      5'b00100:
        casez_tmp_57 = rob_unsafe_1_4;
      5'b00101:
        casez_tmp_57 = rob_unsafe_1_5;
      5'b00110:
        casez_tmp_57 = rob_unsafe_1_6;
      5'b00111:
        casez_tmp_57 = rob_unsafe_1_7;
      5'b01000:
        casez_tmp_57 = rob_unsafe_1_8;
      5'b01001:
        casez_tmp_57 = rob_unsafe_1_9;
      5'b01010:
        casez_tmp_57 = rob_unsafe_1_10;
      5'b01011:
        casez_tmp_57 = rob_unsafe_1_11;
      5'b01100:
        casez_tmp_57 = rob_unsafe_1_12;
      5'b01101:
        casez_tmp_57 = rob_unsafe_1_13;
      5'b01110:
        casez_tmp_57 = rob_unsafe_1_14;
      5'b01111:
        casez_tmp_57 = rob_unsafe_1_15;
      5'b10000:
        casez_tmp_57 = rob_unsafe_1_16;
      5'b10001:
        casez_tmp_57 = rob_unsafe_1_17;
      5'b10010:
        casez_tmp_57 = rob_unsafe_1_18;
      5'b10011:
        casez_tmp_57 = rob_unsafe_1_19;
      5'b10100:
        casez_tmp_57 = rob_unsafe_1_20;
      5'b10101:
        casez_tmp_57 = rob_unsafe_1_21;
      5'b10110:
        casez_tmp_57 = rob_unsafe_1_22;
      5'b10111:
        casez_tmp_57 = rob_unsafe_1_23;
      5'b11000:
        casez_tmp_57 = rob_unsafe_1_24;
      5'b11001:
        casez_tmp_57 = rob_unsafe_1_25;
      5'b11010:
        casez_tmp_57 = rob_unsafe_1_26;
      5'b11011:
        casez_tmp_57 = rob_unsafe_1_27;
      5'b11100:
        casez_tmp_57 = rob_unsafe_1_28;
      5'b11101:
        casez_tmp_57 = rob_unsafe_1_29;
      5'b11110:
        casez_tmp_57 = rob_unsafe_1_30;
      default:
        casez_tmp_57 = rob_unsafe_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_58 = rob_unsafe_1_0;
      5'b00001:
        casez_tmp_58 = rob_unsafe_1_1;
      5'b00010:
        casez_tmp_58 = rob_unsafe_1_2;
      5'b00011:
        casez_tmp_58 = rob_unsafe_1_3;
      5'b00100:
        casez_tmp_58 = rob_unsafe_1_4;
      5'b00101:
        casez_tmp_58 = rob_unsafe_1_5;
      5'b00110:
        casez_tmp_58 = rob_unsafe_1_6;
      5'b00111:
        casez_tmp_58 = rob_unsafe_1_7;
      5'b01000:
        casez_tmp_58 = rob_unsafe_1_8;
      5'b01001:
        casez_tmp_58 = rob_unsafe_1_9;
      5'b01010:
        casez_tmp_58 = rob_unsafe_1_10;
      5'b01011:
        casez_tmp_58 = rob_unsafe_1_11;
      5'b01100:
        casez_tmp_58 = rob_unsafe_1_12;
      5'b01101:
        casez_tmp_58 = rob_unsafe_1_13;
      5'b01110:
        casez_tmp_58 = rob_unsafe_1_14;
      5'b01111:
        casez_tmp_58 = rob_unsafe_1_15;
      5'b10000:
        casez_tmp_58 = rob_unsafe_1_16;
      5'b10001:
        casez_tmp_58 = rob_unsafe_1_17;
      5'b10010:
        casez_tmp_58 = rob_unsafe_1_18;
      5'b10011:
        casez_tmp_58 = rob_unsafe_1_19;
      5'b10100:
        casez_tmp_58 = rob_unsafe_1_20;
      5'b10101:
        casez_tmp_58 = rob_unsafe_1_21;
      5'b10110:
        casez_tmp_58 = rob_unsafe_1_22;
      5'b10111:
        casez_tmp_58 = rob_unsafe_1_23;
      5'b11000:
        casez_tmp_58 = rob_unsafe_1_24;
      5'b11001:
        casez_tmp_58 = rob_unsafe_1_25;
      5'b11010:
        casez_tmp_58 = rob_unsafe_1_26;
      5'b11011:
        casez_tmp_58 = rob_unsafe_1_27;
      5'b11100:
        casez_tmp_58 = rob_unsafe_1_28;
      5'b11101:
        casez_tmp_58 = rob_unsafe_1_29;
      5'b11110:
        casez_tmp_58 = rob_unsafe_1_30;
      default:
        casez_tmp_58 = rob_unsafe_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_59 = rob_exception_1_0;
      5'b00001:
        casez_tmp_59 = rob_exception_1_1;
      5'b00010:
        casez_tmp_59 = rob_exception_1_2;
      5'b00011:
        casez_tmp_59 = rob_exception_1_3;
      5'b00100:
        casez_tmp_59 = rob_exception_1_4;
      5'b00101:
        casez_tmp_59 = rob_exception_1_5;
      5'b00110:
        casez_tmp_59 = rob_exception_1_6;
      5'b00111:
        casez_tmp_59 = rob_exception_1_7;
      5'b01000:
        casez_tmp_59 = rob_exception_1_8;
      5'b01001:
        casez_tmp_59 = rob_exception_1_9;
      5'b01010:
        casez_tmp_59 = rob_exception_1_10;
      5'b01011:
        casez_tmp_59 = rob_exception_1_11;
      5'b01100:
        casez_tmp_59 = rob_exception_1_12;
      5'b01101:
        casez_tmp_59 = rob_exception_1_13;
      5'b01110:
        casez_tmp_59 = rob_exception_1_14;
      5'b01111:
        casez_tmp_59 = rob_exception_1_15;
      5'b10000:
        casez_tmp_59 = rob_exception_1_16;
      5'b10001:
        casez_tmp_59 = rob_exception_1_17;
      5'b10010:
        casez_tmp_59 = rob_exception_1_18;
      5'b10011:
        casez_tmp_59 = rob_exception_1_19;
      5'b10100:
        casez_tmp_59 = rob_exception_1_20;
      5'b10101:
        casez_tmp_59 = rob_exception_1_21;
      5'b10110:
        casez_tmp_59 = rob_exception_1_22;
      5'b10111:
        casez_tmp_59 = rob_exception_1_23;
      5'b11000:
        casez_tmp_59 = rob_exception_1_24;
      5'b11001:
        casez_tmp_59 = rob_exception_1_25;
      5'b11010:
        casez_tmp_59 = rob_exception_1_26;
      5'b11011:
        casez_tmp_59 = rob_exception_1_27;
      5'b11100:
        casez_tmp_59 = rob_exception_1_28;
      5'b11101:
        casez_tmp_59 = rob_exception_1_29;
      5'b11110:
        casez_tmp_59 = rob_exception_1_30;
      default:
        casez_tmp_59 = rob_exception_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_60 = rob_val_1_0;
      5'b00001:
        casez_tmp_60 = rob_val_1_1;
      5'b00010:
        casez_tmp_60 = rob_val_1_2;
      5'b00011:
        casez_tmp_60 = rob_val_1_3;
      5'b00100:
        casez_tmp_60 = rob_val_1_4;
      5'b00101:
        casez_tmp_60 = rob_val_1_5;
      5'b00110:
        casez_tmp_60 = rob_val_1_6;
      5'b00111:
        casez_tmp_60 = rob_val_1_7;
      5'b01000:
        casez_tmp_60 = rob_val_1_8;
      5'b01001:
        casez_tmp_60 = rob_val_1_9;
      5'b01010:
        casez_tmp_60 = rob_val_1_10;
      5'b01011:
        casez_tmp_60 = rob_val_1_11;
      5'b01100:
        casez_tmp_60 = rob_val_1_12;
      5'b01101:
        casez_tmp_60 = rob_val_1_13;
      5'b01110:
        casez_tmp_60 = rob_val_1_14;
      5'b01111:
        casez_tmp_60 = rob_val_1_15;
      5'b10000:
        casez_tmp_60 = rob_val_1_16;
      5'b10001:
        casez_tmp_60 = rob_val_1_17;
      5'b10010:
        casez_tmp_60 = rob_val_1_18;
      5'b10011:
        casez_tmp_60 = rob_val_1_19;
      5'b10100:
        casez_tmp_60 = rob_val_1_20;
      5'b10101:
        casez_tmp_60 = rob_val_1_21;
      5'b10110:
        casez_tmp_60 = rob_val_1_22;
      5'b10111:
        casez_tmp_60 = rob_val_1_23;
      5'b11000:
        casez_tmp_60 = rob_val_1_24;
      5'b11001:
        casez_tmp_60 = rob_val_1_25;
      5'b11010:
        casez_tmp_60 = rob_val_1_26;
      5'b11011:
        casez_tmp_60 = rob_val_1_27;
      5'b11100:
        casez_tmp_60 = rob_val_1_28;
      5'b11101:
        casez_tmp_60 = rob_val_1_29;
      5'b11110:
        casez_tmp_60 = rob_val_1_30;
      default:
        casez_tmp_60 = rob_val_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_61 = rob_val_1_0;
      5'b00001:
        casez_tmp_61 = rob_val_1_1;
      5'b00010:
        casez_tmp_61 = rob_val_1_2;
      5'b00011:
        casez_tmp_61 = rob_val_1_3;
      5'b00100:
        casez_tmp_61 = rob_val_1_4;
      5'b00101:
        casez_tmp_61 = rob_val_1_5;
      5'b00110:
        casez_tmp_61 = rob_val_1_6;
      5'b00111:
        casez_tmp_61 = rob_val_1_7;
      5'b01000:
        casez_tmp_61 = rob_val_1_8;
      5'b01001:
        casez_tmp_61 = rob_val_1_9;
      5'b01010:
        casez_tmp_61 = rob_val_1_10;
      5'b01011:
        casez_tmp_61 = rob_val_1_11;
      5'b01100:
        casez_tmp_61 = rob_val_1_12;
      5'b01101:
        casez_tmp_61 = rob_val_1_13;
      5'b01110:
        casez_tmp_61 = rob_val_1_14;
      5'b01111:
        casez_tmp_61 = rob_val_1_15;
      5'b10000:
        casez_tmp_61 = rob_val_1_16;
      5'b10001:
        casez_tmp_61 = rob_val_1_17;
      5'b10010:
        casez_tmp_61 = rob_val_1_18;
      5'b10011:
        casez_tmp_61 = rob_val_1_19;
      5'b10100:
        casez_tmp_61 = rob_val_1_20;
      5'b10101:
        casez_tmp_61 = rob_val_1_21;
      5'b10110:
        casez_tmp_61 = rob_val_1_22;
      5'b10111:
        casez_tmp_61 = rob_val_1_23;
      5'b11000:
        casez_tmp_61 = rob_val_1_24;
      5'b11001:
        casez_tmp_61 = rob_val_1_25;
      5'b11010:
        casez_tmp_61 = rob_val_1_26;
      5'b11011:
        casez_tmp_61 = rob_val_1_27;
      5'b11100:
        casez_tmp_61 = rob_val_1_28;
      5'b11101:
        casez_tmp_61 = rob_val_1_29;
      5'b11110:
        casez_tmp_61 = rob_val_1_30;
      default:
        casez_tmp_61 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1886 = _GEN_916 & ~casez_tmp_61;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_62 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_62 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_62 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_62 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_62 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_62 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_62 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_62 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_62 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_62 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_62 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_62 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_62 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_62 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_62 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_62 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_62 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_62 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_62 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_62 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_62 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_62 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_62 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_62 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_62 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_62 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_62 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_62 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_62 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_62 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_62 = rob_bsy_1_30;
      default:
        casez_tmp_62 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1887 = _GEN_916 & ~casez_tmp_62;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_63 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_63 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_63 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_63 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_63 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_63 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_63 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_63 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_63 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_63 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_63 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_63 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_63 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_63 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_63 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_63 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_63 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_63 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_63 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_63 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_63 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_63 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_63 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_63 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_63 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_63 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_63 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_63 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_63 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_63 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_63 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_63 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_64 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_64 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_64 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_64 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_64 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_64 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_64 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_64 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_64 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_64 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_64 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_64 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_64 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_64 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_64 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_64 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_64 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_64 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_64 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_64 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_64 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_64 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_64 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_64 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_64 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_64 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_64 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_64 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_64 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_64 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_64 = rob_uop_1_30_pdst;
      default:
        casez_tmp_64 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1888 = _GEN_916 & casez_tmp_63 & casez_tmp_64 != io_wb_resps_0_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_65 = rob_val_1_0;
      5'b00001:
        casez_tmp_65 = rob_val_1_1;
      5'b00010:
        casez_tmp_65 = rob_val_1_2;
      5'b00011:
        casez_tmp_65 = rob_val_1_3;
      5'b00100:
        casez_tmp_65 = rob_val_1_4;
      5'b00101:
        casez_tmp_65 = rob_val_1_5;
      5'b00110:
        casez_tmp_65 = rob_val_1_6;
      5'b00111:
        casez_tmp_65 = rob_val_1_7;
      5'b01000:
        casez_tmp_65 = rob_val_1_8;
      5'b01001:
        casez_tmp_65 = rob_val_1_9;
      5'b01010:
        casez_tmp_65 = rob_val_1_10;
      5'b01011:
        casez_tmp_65 = rob_val_1_11;
      5'b01100:
        casez_tmp_65 = rob_val_1_12;
      5'b01101:
        casez_tmp_65 = rob_val_1_13;
      5'b01110:
        casez_tmp_65 = rob_val_1_14;
      5'b01111:
        casez_tmp_65 = rob_val_1_15;
      5'b10000:
        casez_tmp_65 = rob_val_1_16;
      5'b10001:
        casez_tmp_65 = rob_val_1_17;
      5'b10010:
        casez_tmp_65 = rob_val_1_18;
      5'b10011:
        casez_tmp_65 = rob_val_1_19;
      5'b10100:
        casez_tmp_65 = rob_val_1_20;
      5'b10101:
        casez_tmp_65 = rob_val_1_21;
      5'b10110:
        casez_tmp_65 = rob_val_1_22;
      5'b10111:
        casez_tmp_65 = rob_val_1_23;
      5'b11000:
        casez_tmp_65 = rob_val_1_24;
      5'b11001:
        casez_tmp_65 = rob_val_1_25;
      5'b11010:
        casez_tmp_65 = rob_val_1_26;
      5'b11011:
        casez_tmp_65 = rob_val_1_27;
      5'b11100:
        casez_tmp_65 = rob_val_1_28;
      5'b11101:
        casez_tmp_65 = rob_val_1_29;
      5'b11110:
        casez_tmp_65 = rob_val_1_30;
      default:
        casez_tmp_65 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1889 = _GEN_467 & ~casez_tmp_65;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_66 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_66 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_66 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_66 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_66 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_66 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_66 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_66 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_66 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_66 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_66 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_66 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_66 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_66 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_66 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_66 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_66 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_66 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_66 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_66 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_66 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_66 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_66 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_66 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_66 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_66 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_66 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_66 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_66 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_66 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_66 = rob_bsy_1_30;
      default:
        casez_tmp_66 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1890 = _GEN_467 & ~casez_tmp_66;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_67 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_67 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_67 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_67 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_67 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_67 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_67 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_67 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_67 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_67 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_67 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_67 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_67 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_67 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_67 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_67 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_67 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_67 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_67 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_67 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_67 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_67 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_67 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_67 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_67 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_67 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_67 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_67 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_67 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_67 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_67 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_67 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_68 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_68 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_68 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_68 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_68 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_68 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_68 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_68 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_68 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_68 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_68 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_68 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_68 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_68 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_68 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_68 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_68 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_68 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_68 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_68 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_68 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_68 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_68 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_68 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_68 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_68 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_68 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_68 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_68 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_68 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_68 = rob_uop_1_30_pdst;
      default:
        casez_tmp_68 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1891 = _GEN_467 & casez_tmp_67 & casez_tmp_68 != io_wb_resps_1_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_69 = rob_val_1_0;
      5'b00001:
        casez_tmp_69 = rob_val_1_1;
      5'b00010:
        casez_tmp_69 = rob_val_1_2;
      5'b00011:
        casez_tmp_69 = rob_val_1_3;
      5'b00100:
        casez_tmp_69 = rob_val_1_4;
      5'b00101:
        casez_tmp_69 = rob_val_1_5;
      5'b00110:
        casez_tmp_69 = rob_val_1_6;
      5'b00111:
        casez_tmp_69 = rob_val_1_7;
      5'b01000:
        casez_tmp_69 = rob_val_1_8;
      5'b01001:
        casez_tmp_69 = rob_val_1_9;
      5'b01010:
        casez_tmp_69 = rob_val_1_10;
      5'b01011:
        casez_tmp_69 = rob_val_1_11;
      5'b01100:
        casez_tmp_69 = rob_val_1_12;
      5'b01101:
        casez_tmp_69 = rob_val_1_13;
      5'b01110:
        casez_tmp_69 = rob_val_1_14;
      5'b01111:
        casez_tmp_69 = rob_val_1_15;
      5'b10000:
        casez_tmp_69 = rob_val_1_16;
      5'b10001:
        casez_tmp_69 = rob_val_1_17;
      5'b10010:
        casez_tmp_69 = rob_val_1_18;
      5'b10011:
        casez_tmp_69 = rob_val_1_19;
      5'b10100:
        casez_tmp_69 = rob_val_1_20;
      5'b10101:
        casez_tmp_69 = rob_val_1_21;
      5'b10110:
        casez_tmp_69 = rob_val_1_22;
      5'b10111:
        casez_tmp_69 = rob_val_1_23;
      5'b11000:
        casez_tmp_69 = rob_val_1_24;
      5'b11001:
        casez_tmp_69 = rob_val_1_25;
      5'b11010:
        casez_tmp_69 = rob_val_1_26;
      5'b11011:
        casez_tmp_69 = rob_val_1_27;
      5'b11100:
        casez_tmp_69 = rob_val_1_28;
      5'b11101:
        casez_tmp_69 = rob_val_1_29;
      5'b11110:
        casez_tmp_69 = rob_val_1_30;
      default:
        casez_tmp_69 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1892 = _GEN_917 & ~casez_tmp_69;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_70 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_70 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_70 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_70 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_70 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_70 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_70 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_70 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_70 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_70 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_70 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_70 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_70 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_70 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_70 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_70 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_70 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_70 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_70 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_70 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_70 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_70 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_70 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_70 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_70 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_70 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_70 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_70 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_70 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_70 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_70 = rob_bsy_1_30;
      default:
        casez_tmp_70 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1893 = _GEN_917 & ~casez_tmp_70;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_71 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_71 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_71 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_71 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_71 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_71 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_71 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_71 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_71 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_71 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_71 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_71 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_71 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_71 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_71 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_71 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_71 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_71 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_71 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_71 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_71 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_71 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_71 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_71 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_71 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_71 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_71 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_71 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_71 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_71 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_71 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_71 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_72 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_72 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_72 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_72 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_72 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_72 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_72 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_72 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_72 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_72 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_72 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_72 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_72 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_72 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_72 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_72 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_72 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_72 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_72 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_72 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_72 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_72 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_72 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_72 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_72 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_72 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_72 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_72 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_72 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_72 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_72 = rob_uop_1_30_pdst;
      default:
        casez_tmp_72 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1894 = _GEN_917 & casez_tmp_71 & casez_tmp_72 != io_wb_resps_2_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_73 = rob_val_1_0;
      5'b00001:
        casez_tmp_73 = rob_val_1_1;
      5'b00010:
        casez_tmp_73 = rob_val_1_2;
      5'b00011:
        casez_tmp_73 = rob_val_1_3;
      5'b00100:
        casez_tmp_73 = rob_val_1_4;
      5'b00101:
        casez_tmp_73 = rob_val_1_5;
      5'b00110:
        casez_tmp_73 = rob_val_1_6;
      5'b00111:
        casez_tmp_73 = rob_val_1_7;
      5'b01000:
        casez_tmp_73 = rob_val_1_8;
      5'b01001:
        casez_tmp_73 = rob_val_1_9;
      5'b01010:
        casez_tmp_73 = rob_val_1_10;
      5'b01011:
        casez_tmp_73 = rob_val_1_11;
      5'b01100:
        casez_tmp_73 = rob_val_1_12;
      5'b01101:
        casez_tmp_73 = rob_val_1_13;
      5'b01110:
        casez_tmp_73 = rob_val_1_14;
      5'b01111:
        casez_tmp_73 = rob_val_1_15;
      5'b10000:
        casez_tmp_73 = rob_val_1_16;
      5'b10001:
        casez_tmp_73 = rob_val_1_17;
      5'b10010:
        casez_tmp_73 = rob_val_1_18;
      5'b10011:
        casez_tmp_73 = rob_val_1_19;
      5'b10100:
        casez_tmp_73 = rob_val_1_20;
      5'b10101:
        casez_tmp_73 = rob_val_1_21;
      5'b10110:
        casez_tmp_73 = rob_val_1_22;
      5'b10111:
        casez_tmp_73 = rob_val_1_23;
      5'b11000:
        casez_tmp_73 = rob_val_1_24;
      5'b11001:
        casez_tmp_73 = rob_val_1_25;
      5'b11010:
        casez_tmp_73 = rob_val_1_26;
      5'b11011:
        casez_tmp_73 = rob_val_1_27;
      5'b11100:
        casez_tmp_73 = rob_val_1_28;
      5'b11101:
        casez_tmp_73 = rob_val_1_29;
      5'b11110:
        casez_tmp_73 = rob_val_1_30;
      default:
        casez_tmp_73 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1895 = _GEN_466 & ~casez_tmp_73;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_74 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_74 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_74 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_74 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_74 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_74 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_74 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_74 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_74 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_74 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_74 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_74 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_74 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_74 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_74 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_74 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_74 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_74 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_74 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_74 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_74 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_74 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_74 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_74 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_74 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_74 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_74 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_74 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_74 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_74 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_74 = rob_bsy_1_30;
      default:
        casez_tmp_74 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1896 = _GEN_466 & ~casez_tmp_74;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_75 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_75 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_75 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_75 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_75 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_75 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_75 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_75 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_75 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_75 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_75 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_75 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_75 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_75 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_75 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_75 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_75 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_75 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_75 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_75 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_75 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_75 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_75 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_75 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_75 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_75 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_75 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_75 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_75 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_75 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_75 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_75 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_76 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_76 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_76 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_76 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_76 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_76 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_76 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_76 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_76 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_76 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_76 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_76 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_76 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_76 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_76 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_76 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_76 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_76 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_76 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_76 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_76 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_76 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_76 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_76 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_76 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_76 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_76 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_76 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_76 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_76 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_76 = rob_uop_1_30_pdst;
      default:
        casez_tmp_76 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1897 = _GEN_466 & casez_tmp_75 & casez_tmp_76 != io_wb_resps_3_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_77 = rob_val_1_0;
      5'b00001:
        casez_tmp_77 = rob_val_1_1;
      5'b00010:
        casez_tmp_77 = rob_val_1_2;
      5'b00011:
        casez_tmp_77 = rob_val_1_3;
      5'b00100:
        casez_tmp_77 = rob_val_1_4;
      5'b00101:
        casez_tmp_77 = rob_val_1_5;
      5'b00110:
        casez_tmp_77 = rob_val_1_6;
      5'b00111:
        casez_tmp_77 = rob_val_1_7;
      5'b01000:
        casez_tmp_77 = rob_val_1_8;
      5'b01001:
        casez_tmp_77 = rob_val_1_9;
      5'b01010:
        casez_tmp_77 = rob_val_1_10;
      5'b01011:
        casez_tmp_77 = rob_val_1_11;
      5'b01100:
        casez_tmp_77 = rob_val_1_12;
      5'b01101:
        casez_tmp_77 = rob_val_1_13;
      5'b01110:
        casez_tmp_77 = rob_val_1_14;
      5'b01111:
        casez_tmp_77 = rob_val_1_15;
      5'b10000:
        casez_tmp_77 = rob_val_1_16;
      5'b10001:
        casez_tmp_77 = rob_val_1_17;
      5'b10010:
        casez_tmp_77 = rob_val_1_18;
      5'b10011:
        casez_tmp_77 = rob_val_1_19;
      5'b10100:
        casez_tmp_77 = rob_val_1_20;
      5'b10101:
        casez_tmp_77 = rob_val_1_21;
      5'b10110:
        casez_tmp_77 = rob_val_1_22;
      5'b10111:
        casez_tmp_77 = rob_val_1_23;
      5'b11000:
        casez_tmp_77 = rob_val_1_24;
      5'b11001:
        casez_tmp_77 = rob_val_1_25;
      5'b11010:
        casez_tmp_77 = rob_val_1_26;
      5'b11011:
        casez_tmp_77 = rob_val_1_27;
      5'b11100:
        casez_tmp_77 = rob_val_1_28;
      5'b11101:
        casez_tmp_77 = rob_val_1_29;
      5'b11110:
        casez_tmp_77 = rob_val_1_30;
      default:
        casez_tmp_77 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1898 = _GEN_918 & ~casez_tmp_77;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_78 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_78 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_78 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_78 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_78 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_78 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_78 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_78 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_78 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_78 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_78 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_78 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_78 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_78 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_78 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_78 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_78 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_78 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_78 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_78 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_78 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_78 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_78 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_78 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_78 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_78 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_78 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_78 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_78 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_78 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_78 = rob_bsy_1_30;
      default:
        casez_tmp_78 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1899 = _GEN_918 & ~casez_tmp_78;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_79 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_79 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_79 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_79 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_79 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_79 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_79 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_79 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_79 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_79 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_79 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_79 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_79 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_79 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_79 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_79 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_79 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_79 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_79 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_79 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_79 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_79 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_79 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_79 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_79 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_79 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_79 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_79 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_79 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_79 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_79 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_79 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_80 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_80 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_80 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_80 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_80 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_80 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_80 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_80 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_80 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_80 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_80 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_80 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_80 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_80 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_80 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_80 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_80 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_80 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_80 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_80 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_80 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_80 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_80 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_80 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_80 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_80 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_80 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_80 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_80 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_80 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_80 = rob_uop_1_30_pdst;
      default:
        casez_tmp_80 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1900 = _GEN_918 & casez_tmp_79 & casez_tmp_80 != io_wb_resps_4_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_81 = rob_val_1_0;
      5'b00001:
        casez_tmp_81 = rob_val_1_1;
      5'b00010:
        casez_tmp_81 = rob_val_1_2;
      5'b00011:
        casez_tmp_81 = rob_val_1_3;
      5'b00100:
        casez_tmp_81 = rob_val_1_4;
      5'b00101:
        casez_tmp_81 = rob_val_1_5;
      5'b00110:
        casez_tmp_81 = rob_val_1_6;
      5'b00111:
        casez_tmp_81 = rob_val_1_7;
      5'b01000:
        casez_tmp_81 = rob_val_1_8;
      5'b01001:
        casez_tmp_81 = rob_val_1_9;
      5'b01010:
        casez_tmp_81 = rob_val_1_10;
      5'b01011:
        casez_tmp_81 = rob_val_1_11;
      5'b01100:
        casez_tmp_81 = rob_val_1_12;
      5'b01101:
        casez_tmp_81 = rob_val_1_13;
      5'b01110:
        casez_tmp_81 = rob_val_1_14;
      5'b01111:
        casez_tmp_81 = rob_val_1_15;
      5'b10000:
        casez_tmp_81 = rob_val_1_16;
      5'b10001:
        casez_tmp_81 = rob_val_1_17;
      5'b10010:
        casez_tmp_81 = rob_val_1_18;
      5'b10011:
        casez_tmp_81 = rob_val_1_19;
      5'b10100:
        casez_tmp_81 = rob_val_1_20;
      5'b10101:
        casez_tmp_81 = rob_val_1_21;
      5'b10110:
        casez_tmp_81 = rob_val_1_22;
      5'b10111:
        casez_tmp_81 = rob_val_1_23;
      5'b11000:
        casez_tmp_81 = rob_val_1_24;
      5'b11001:
        casez_tmp_81 = rob_val_1_25;
      5'b11010:
        casez_tmp_81 = rob_val_1_26;
      5'b11011:
        casez_tmp_81 = rob_val_1_27;
      5'b11100:
        casez_tmp_81 = rob_val_1_28;
      5'b11101:
        casez_tmp_81 = rob_val_1_29;
      5'b11110:
        casez_tmp_81 = rob_val_1_30;
      default:
        casez_tmp_81 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1901 = _GEN_465 & ~casez_tmp_81;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_82 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_82 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_82 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_82 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_82 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_82 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_82 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_82 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_82 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_82 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_82 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_82 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_82 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_82 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_82 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_82 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_82 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_82 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_82 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_82 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_82 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_82 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_82 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_82 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_82 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_82 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_82 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_82 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_82 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_82 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_82 = rob_bsy_1_30;
      default:
        casez_tmp_82 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1902 = _GEN_465 & ~casez_tmp_82;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_83 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_83 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_83 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_83 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_83 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_83 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_83 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_83 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_83 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_83 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_83 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_83 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_83 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_83 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_83 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_83 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_83 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_83 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_83 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_83 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_83 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_83 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_83 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_83 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_83 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_83 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_83 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_83 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_83 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_83 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_83 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_83 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_84 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_84 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_84 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_84 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_84 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_84 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_84 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_84 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_84 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_84 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_84 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_84 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_84 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_84 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_84 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_84 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_84 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_84 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_84 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_84 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_84 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_84 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_84 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_84 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_84 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_84 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_84 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_84 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_84 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_84 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_84 = rob_uop_1_30_pdst;
      default:
        casez_tmp_84 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1903 = _GEN_465 & casez_tmp_83 & casez_tmp_84 != io_wb_resps_5_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_85 = rob_val_1_0;
      5'b00001:
        casez_tmp_85 = rob_val_1_1;
      5'b00010:
        casez_tmp_85 = rob_val_1_2;
      5'b00011:
        casez_tmp_85 = rob_val_1_3;
      5'b00100:
        casez_tmp_85 = rob_val_1_4;
      5'b00101:
        casez_tmp_85 = rob_val_1_5;
      5'b00110:
        casez_tmp_85 = rob_val_1_6;
      5'b00111:
        casez_tmp_85 = rob_val_1_7;
      5'b01000:
        casez_tmp_85 = rob_val_1_8;
      5'b01001:
        casez_tmp_85 = rob_val_1_9;
      5'b01010:
        casez_tmp_85 = rob_val_1_10;
      5'b01011:
        casez_tmp_85 = rob_val_1_11;
      5'b01100:
        casez_tmp_85 = rob_val_1_12;
      5'b01101:
        casez_tmp_85 = rob_val_1_13;
      5'b01110:
        casez_tmp_85 = rob_val_1_14;
      5'b01111:
        casez_tmp_85 = rob_val_1_15;
      5'b10000:
        casez_tmp_85 = rob_val_1_16;
      5'b10001:
        casez_tmp_85 = rob_val_1_17;
      5'b10010:
        casez_tmp_85 = rob_val_1_18;
      5'b10011:
        casez_tmp_85 = rob_val_1_19;
      5'b10100:
        casez_tmp_85 = rob_val_1_20;
      5'b10101:
        casez_tmp_85 = rob_val_1_21;
      5'b10110:
        casez_tmp_85 = rob_val_1_22;
      5'b10111:
        casez_tmp_85 = rob_val_1_23;
      5'b11000:
        casez_tmp_85 = rob_val_1_24;
      5'b11001:
        casez_tmp_85 = rob_val_1_25;
      5'b11010:
        casez_tmp_85 = rob_val_1_26;
      5'b11011:
        casez_tmp_85 = rob_val_1_27;
      5'b11100:
        casez_tmp_85 = rob_val_1_28;
      5'b11101:
        casez_tmp_85 = rob_val_1_29;
      5'b11110:
        casez_tmp_85 = rob_val_1_30;
      default:
        casez_tmp_85 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1904 = _GEN_919 & ~casez_tmp_85;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_86 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_86 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_86 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_86 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_86 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_86 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_86 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_86 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_86 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_86 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_86 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_86 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_86 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_86 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_86 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_86 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_86 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_86 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_86 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_86 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_86 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_86 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_86 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_86 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_86 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_86 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_86 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_86 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_86 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_86 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_86 = rob_bsy_1_30;
      default:
        casez_tmp_86 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1905 = _GEN_919 & ~casez_tmp_86;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_87 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_87 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_87 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_87 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_87 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_87 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_87 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_87 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_87 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_87 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_87 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_87 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_87 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_87 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_87 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_87 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_87 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_87 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_87 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_87 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_87 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_87 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_87 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_87 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_87 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_87 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_87 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_87 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_87 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_87 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_87 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_87 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_88 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_88 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_88 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_88 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_88 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_88 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_88 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_88 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_88 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_88 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_88 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_88 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_88 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_88 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_88 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_88 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_88 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_88 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_88 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_88 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_88 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_88 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_88 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_88 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_88 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_88 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_88 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_88 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_88 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_88 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_88 = rob_uop_1_30_pdst;
      default:
        casez_tmp_88 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1906 = _GEN_919 & casez_tmp_87 & casez_tmp_88 != io_wb_resps_6_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_89 = rob_val_1_0;
      5'b00001:
        casez_tmp_89 = rob_val_1_1;
      5'b00010:
        casez_tmp_89 = rob_val_1_2;
      5'b00011:
        casez_tmp_89 = rob_val_1_3;
      5'b00100:
        casez_tmp_89 = rob_val_1_4;
      5'b00101:
        casez_tmp_89 = rob_val_1_5;
      5'b00110:
        casez_tmp_89 = rob_val_1_6;
      5'b00111:
        casez_tmp_89 = rob_val_1_7;
      5'b01000:
        casez_tmp_89 = rob_val_1_8;
      5'b01001:
        casez_tmp_89 = rob_val_1_9;
      5'b01010:
        casez_tmp_89 = rob_val_1_10;
      5'b01011:
        casez_tmp_89 = rob_val_1_11;
      5'b01100:
        casez_tmp_89 = rob_val_1_12;
      5'b01101:
        casez_tmp_89 = rob_val_1_13;
      5'b01110:
        casez_tmp_89 = rob_val_1_14;
      5'b01111:
        casez_tmp_89 = rob_val_1_15;
      5'b10000:
        casez_tmp_89 = rob_val_1_16;
      5'b10001:
        casez_tmp_89 = rob_val_1_17;
      5'b10010:
        casez_tmp_89 = rob_val_1_18;
      5'b10011:
        casez_tmp_89 = rob_val_1_19;
      5'b10100:
        casez_tmp_89 = rob_val_1_20;
      5'b10101:
        casez_tmp_89 = rob_val_1_21;
      5'b10110:
        casez_tmp_89 = rob_val_1_22;
      5'b10111:
        casez_tmp_89 = rob_val_1_23;
      5'b11000:
        casez_tmp_89 = rob_val_1_24;
      5'b11001:
        casez_tmp_89 = rob_val_1_25;
      5'b11010:
        casez_tmp_89 = rob_val_1_26;
      5'b11011:
        casez_tmp_89 = rob_val_1_27;
      5'b11100:
        casez_tmp_89 = rob_val_1_28;
      5'b11101:
        casez_tmp_89 = rob_val_1_29;
      5'b11110:
        casez_tmp_89 = rob_val_1_30;
      default:
        casez_tmp_89 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1907 = _GEN_464 & ~casez_tmp_89;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_90 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_90 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_90 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_90 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_90 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_90 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_90 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_90 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_90 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_90 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_90 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_90 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_90 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_90 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_90 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_90 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_90 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_90 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_90 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_90 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_90 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_90 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_90 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_90 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_90 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_90 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_90 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_90 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_90 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_90 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_90 = rob_bsy_1_30;
      default:
        casez_tmp_90 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1908 = _GEN_464 & ~casez_tmp_90;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_91 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_91 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_91 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_91 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_91 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_91 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_91 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_91 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_91 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_91 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_91 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_91 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_91 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_91 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_91 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_91 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_91 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_91 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_91 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_91 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_91 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_91 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_91 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_91 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_91 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_91 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_91 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_91 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_91 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_91 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_91 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_91 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_92 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_92 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_92 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_92 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_92 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_92 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_92 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_92 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_92 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_92 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_92 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_92 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_92 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_92 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_92 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_92 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_92 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_92 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_92 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_92 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_92 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_92 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_92 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_92 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_92 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_92 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_92 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_92 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_92 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_92 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_92 = rob_uop_1_30_pdst;
      default:
        casez_tmp_92 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1909 = _GEN_464 & casez_tmp_91 & casez_tmp_92 != io_wb_resps_7_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_93 = rob_val_1_0;
      5'b00001:
        casez_tmp_93 = rob_val_1_1;
      5'b00010:
        casez_tmp_93 = rob_val_1_2;
      5'b00011:
        casez_tmp_93 = rob_val_1_3;
      5'b00100:
        casez_tmp_93 = rob_val_1_4;
      5'b00101:
        casez_tmp_93 = rob_val_1_5;
      5'b00110:
        casez_tmp_93 = rob_val_1_6;
      5'b00111:
        casez_tmp_93 = rob_val_1_7;
      5'b01000:
        casez_tmp_93 = rob_val_1_8;
      5'b01001:
        casez_tmp_93 = rob_val_1_9;
      5'b01010:
        casez_tmp_93 = rob_val_1_10;
      5'b01011:
        casez_tmp_93 = rob_val_1_11;
      5'b01100:
        casez_tmp_93 = rob_val_1_12;
      5'b01101:
        casez_tmp_93 = rob_val_1_13;
      5'b01110:
        casez_tmp_93 = rob_val_1_14;
      5'b01111:
        casez_tmp_93 = rob_val_1_15;
      5'b10000:
        casez_tmp_93 = rob_val_1_16;
      5'b10001:
        casez_tmp_93 = rob_val_1_17;
      5'b10010:
        casez_tmp_93 = rob_val_1_18;
      5'b10011:
        casez_tmp_93 = rob_val_1_19;
      5'b10100:
        casez_tmp_93 = rob_val_1_20;
      5'b10101:
        casez_tmp_93 = rob_val_1_21;
      5'b10110:
        casez_tmp_93 = rob_val_1_22;
      5'b10111:
        casez_tmp_93 = rob_val_1_23;
      5'b11000:
        casez_tmp_93 = rob_val_1_24;
      5'b11001:
        casez_tmp_93 = rob_val_1_25;
      5'b11010:
        casez_tmp_93 = rob_val_1_26;
      5'b11011:
        casez_tmp_93 = rob_val_1_27;
      5'b11100:
        casez_tmp_93 = rob_val_1_28;
      5'b11101:
        casez_tmp_93 = rob_val_1_29;
      5'b11110:
        casez_tmp_93 = rob_val_1_30;
      default:
        casez_tmp_93 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1910 = _GEN_920 & ~casez_tmp_93;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_94 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_94 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_94 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_94 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_94 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_94 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_94 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_94 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_94 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_94 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_94 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_94 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_94 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_94 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_94 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_94 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_94 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_94 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_94 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_94 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_94 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_94 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_94 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_94 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_94 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_94 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_94 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_94 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_94 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_94 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_94 = rob_bsy_1_30;
      default:
        casez_tmp_94 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1911 = _GEN_920 & ~casez_tmp_94;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_95 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_95 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_95 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_95 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_95 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_95 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_95 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_95 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_95 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_95 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_95 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_95 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_95 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_95 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_95 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_95 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_95 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_95 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_95 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_95 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_95 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_95 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_95 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_95 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_95 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_95 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_95 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_95 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_95 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_95 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_95 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_95 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_96 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_96 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_96 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_96 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_96 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_96 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_96 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_96 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_96 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_96 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_96 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_96 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_96 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_96 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_96 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_96 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_96 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_96 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_96 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_96 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_96 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_96 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_96 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_96 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_96 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_96 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_96 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_96 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_96 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_96 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_96 = rob_uop_1_30_pdst;
      default:
        casez_tmp_96 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1912 = _GEN_920 & casez_tmp_95 & casez_tmp_96 != io_wb_resps_8_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_97 = rob_val_1_0;
      5'b00001:
        casez_tmp_97 = rob_val_1_1;
      5'b00010:
        casez_tmp_97 = rob_val_1_2;
      5'b00011:
        casez_tmp_97 = rob_val_1_3;
      5'b00100:
        casez_tmp_97 = rob_val_1_4;
      5'b00101:
        casez_tmp_97 = rob_val_1_5;
      5'b00110:
        casez_tmp_97 = rob_val_1_6;
      5'b00111:
        casez_tmp_97 = rob_val_1_7;
      5'b01000:
        casez_tmp_97 = rob_val_1_8;
      5'b01001:
        casez_tmp_97 = rob_val_1_9;
      5'b01010:
        casez_tmp_97 = rob_val_1_10;
      5'b01011:
        casez_tmp_97 = rob_val_1_11;
      5'b01100:
        casez_tmp_97 = rob_val_1_12;
      5'b01101:
        casez_tmp_97 = rob_val_1_13;
      5'b01110:
        casez_tmp_97 = rob_val_1_14;
      5'b01111:
        casez_tmp_97 = rob_val_1_15;
      5'b10000:
        casez_tmp_97 = rob_val_1_16;
      5'b10001:
        casez_tmp_97 = rob_val_1_17;
      5'b10010:
        casez_tmp_97 = rob_val_1_18;
      5'b10011:
        casez_tmp_97 = rob_val_1_19;
      5'b10100:
        casez_tmp_97 = rob_val_1_20;
      5'b10101:
        casez_tmp_97 = rob_val_1_21;
      5'b10110:
        casez_tmp_97 = rob_val_1_22;
      5'b10111:
        casez_tmp_97 = rob_val_1_23;
      5'b11000:
        casez_tmp_97 = rob_val_1_24;
      5'b11001:
        casez_tmp_97 = rob_val_1_25;
      5'b11010:
        casez_tmp_97 = rob_val_1_26;
      5'b11011:
        casez_tmp_97 = rob_val_1_27;
      5'b11100:
        casez_tmp_97 = rob_val_1_28;
      5'b11101:
        casez_tmp_97 = rob_val_1_29;
      5'b11110:
        casez_tmp_97 = rob_val_1_30;
      default:
        casez_tmp_97 = rob_val_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1913 = _GEN_463 & ~casez_tmp_97;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_98 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_98 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_98 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_98 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_98 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_98 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_98 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_98 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_98 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_98 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_98 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_98 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_98 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_98 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_98 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_98 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_98 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_98 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_98 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_98 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_98 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_98 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_98 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_98 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_98 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_98 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_98 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_98 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_98 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_98 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_98 = rob_bsy_1_30;
      default:
        casez_tmp_98 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire       _GEN_1914 = _GEN_463 & ~casez_tmp_98;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_99 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_99 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_99 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_99 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_99 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_99 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_99 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_99 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_99 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_99 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_99 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_99 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_99 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_99 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_99 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_99 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_99 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_99 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_99 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_99 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_99 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_99 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_99 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_99 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_99 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_99 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_99 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_99 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_99 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_99 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_99 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_99 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_100 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_100 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_100 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_100 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_100 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_100 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_100 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_100 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_100 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_100 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_100 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_100 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_100 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_100 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_100 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_100 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_100 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_100 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_100 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_100 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_100 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_100 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_100 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_100 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_100 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_100 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_100 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_100 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_100 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_100 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_100 = rob_uop_1_30_pdst;
      default:
        casez_tmp_100 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1915 = _GEN_463 & casez_tmp_99 & casez_tmp_100 != io_wb_resps_9_bits_uop_pdst;
  reg        rob_unsafe_2_0;
  reg        rob_unsafe_2_1;
  reg        rob_unsafe_2_2;
  reg        rob_unsafe_2_3;
  reg        rob_unsafe_2_4;
  reg        rob_unsafe_2_5;
  reg        rob_unsafe_2_6;
  reg        rob_unsafe_2_7;
  reg        rob_unsafe_2_8;
  reg        rob_unsafe_2_9;
  reg        rob_unsafe_2_10;
  reg        rob_unsafe_2_11;
  reg        rob_unsafe_2_12;
  reg        rob_unsafe_2_13;
  reg        rob_unsafe_2_14;
  reg        rob_unsafe_2_15;
  reg        rob_unsafe_2_16;
  reg        rob_unsafe_2_17;
  reg        rob_unsafe_2_18;
  reg        rob_unsafe_2_19;
  reg        rob_unsafe_2_20;
  reg        rob_unsafe_2_21;
  reg        rob_unsafe_2_22;
  reg        rob_unsafe_2_23;
  reg        rob_unsafe_2_24;
  reg        rob_unsafe_2_25;
  reg        rob_unsafe_2_26;
  reg        rob_unsafe_2_27;
  reg        rob_unsafe_2_28;
  reg        rob_unsafe_2_29;
  reg        rob_unsafe_2_30;
  reg        rob_unsafe_2_31;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp_101 = rob_val_2_0;
      5'b00001:
        casez_tmp_101 = rob_val_2_1;
      5'b00010:
        casez_tmp_101 = rob_val_2_2;
      5'b00011:
        casez_tmp_101 = rob_val_2_3;
      5'b00100:
        casez_tmp_101 = rob_val_2_4;
      5'b00101:
        casez_tmp_101 = rob_val_2_5;
      5'b00110:
        casez_tmp_101 = rob_val_2_6;
      5'b00111:
        casez_tmp_101 = rob_val_2_7;
      5'b01000:
        casez_tmp_101 = rob_val_2_8;
      5'b01001:
        casez_tmp_101 = rob_val_2_9;
      5'b01010:
        casez_tmp_101 = rob_val_2_10;
      5'b01011:
        casez_tmp_101 = rob_val_2_11;
      5'b01100:
        casez_tmp_101 = rob_val_2_12;
      5'b01101:
        casez_tmp_101 = rob_val_2_13;
      5'b01110:
        casez_tmp_101 = rob_val_2_14;
      5'b01111:
        casez_tmp_101 = rob_val_2_15;
      5'b10000:
        casez_tmp_101 = rob_val_2_16;
      5'b10001:
        casez_tmp_101 = rob_val_2_17;
      5'b10010:
        casez_tmp_101 = rob_val_2_18;
      5'b10011:
        casez_tmp_101 = rob_val_2_19;
      5'b10100:
        casez_tmp_101 = rob_val_2_20;
      5'b10101:
        casez_tmp_101 = rob_val_2_21;
      5'b10110:
        casez_tmp_101 = rob_val_2_22;
      5'b10111:
        casez_tmp_101 = rob_val_2_23;
      5'b11000:
        casez_tmp_101 = rob_val_2_24;
      5'b11001:
        casez_tmp_101 = rob_val_2_25;
      5'b11010:
        casez_tmp_101 = rob_val_2_26;
      5'b11011:
        casez_tmp_101 = rob_val_2_27;
      5'b11100:
        casez_tmp_101 = rob_val_2_28;
      5'b11101:
        casez_tmp_101 = rob_val_2_29;
      5'b11110:
        casez_tmp_101 = rob_val_2_30;
      default:
        casez_tmp_101 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1916 = io_enq_uops_2_rob_idx[6:2] == rob_tail;
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_102 = rob_val_2_0;
      5'b00001:
        casez_tmp_102 = rob_val_2_1;
      5'b00010:
        casez_tmp_102 = rob_val_2_2;
      5'b00011:
        casez_tmp_102 = rob_val_2_3;
      5'b00100:
        casez_tmp_102 = rob_val_2_4;
      5'b00101:
        casez_tmp_102 = rob_val_2_5;
      5'b00110:
        casez_tmp_102 = rob_val_2_6;
      5'b00111:
        casez_tmp_102 = rob_val_2_7;
      5'b01000:
        casez_tmp_102 = rob_val_2_8;
      5'b01001:
        casez_tmp_102 = rob_val_2_9;
      5'b01010:
        casez_tmp_102 = rob_val_2_10;
      5'b01011:
        casez_tmp_102 = rob_val_2_11;
      5'b01100:
        casez_tmp_102 = rob_val_2_12;
      5'b01101:
        casez_tmp_102 = rob_val_2_13;
      5'b01110:
        casez_tmp_102 = rob_val_2_14;
      5'b01111:
        casez_tmp_102 = rob_val_2_15;
      5'b10000:
        casez_tmp_102 = rob_val_2_16;
      5'b10001:
        casez_tmp_102 = rob_val_2_17;
      5'b10010:
        casez_tmp_102 = rob_val_2_18;
      5'b10011:
        casez_tmp_102 = rob_val_2_19;
      5'b10100:
        casez_tmp_102 = rob_val_2_20;
      5'b10101:
        casez_tmp_102 = rob_val_2_21;
      5'b10110:
        casez_tmp_102 = rob_val_2_22;
      5'b10111:
        casez_tmp_102 = rob_val_2_23;
      5'b11000:
        casez_tmp_102 = rob_val_2_24;
      5'b11001:
        casez_tmp_102 = rob_val_2_25;
      5'b11010:
        casez_tmp_102 = rob_val_2_26;
      5'b11011:
        casez_tmp_102 = rob_val_2_27;
      5'b11100:
        casez_tmp_102 = rob_val_2_28;
      5'b11101:
        casez_tmp_102 = rob_val_2_29;
      5'b11110:
        casez_tmp_102 = rob_val_2_30;
      default:
        casez_tmp_102 = rob_val_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_103 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_103 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_103 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_103 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_103 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_103 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_103 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_103 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_103 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_103 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_103 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_103 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_103 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_103 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_103 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_103 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_103 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_103 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_103 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_103 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_103 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_103 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_103 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_103 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_103 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_103 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_103 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_103 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_103 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_103 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_103 = rob_bsy_2_30;
      default:
        casez_tmp_103 = rob_bsy_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_104 = rob_val_2_0;
      5'b00001:
        casez_tmp_104 = rob_val_2_1;
      5'b00010:
        casez_tmp_104 = rob_val_2_2;
      5'b00011:
        casez_tmp_104 = rob_val_2_3;
      5'b00100:
        casez_tmp_104 = rob_val_2_4;
      5'b00101:
        casez_tmp_104 = rob_val_2_5;
      5'b00110:
        casez_tmp_104 = rob_val_2_6;
      5'b00111:
        casez_tmp_104 = rob_val_2_7;
      5'b01000:
        casez_tmp_104 = rob_val_2_8;
      5'b01001:
        casez_tmp_104 = rob_val_2_9;
      5'b01010:
        casez_tmp_104 = rob_val_2_10;
      5'b01011:
        casez_tmp_104 = rob_val_2_11;
      5'b01100:
        casez_tmp_104 = rob_val_2_12;
      5'b01101:
        casez_tmp_104 = rob_val_2_13;
      5'b01110:
        casez_tmp_104 = rob_val_2_14;
      5'b01111:
        casez_tmp_104 = rob_val_2_15;
      5'b10000:
        casez_tmp_104 = rob_val_2_16;
      5'b10001:
        casez_tmp_104 = rob_val_2_17;
      5'b10010:
        casez_tmp_104 = rob_val_2_18;
      5'b10011:
        casez_tmp_104 = rob_val_2_19;
      5'b10100:
        casez_tmp_104 = rob_val_2_20;
      5'b10101:
        casez_tmp_104 = rob_val_2_21;
      5'b10110:
        casez_tmp_104 = rob_val_2_22;
      5'b10111:
        casez_tmp_104 = rob_val_2_23;
      5'b11000:
        casez_tmp_104 = rob_val_2_24;
      5'b11001:
        casez_tmp_104 = rob_val_2_25;
      5'b11010:
        casez_tmp_104 = rob_val_2_26;
      5'b11011:
        casez_tmp_104 = rob_val_2_27;
      5'b11100:
        casez_tmp_104 = rob_val_2_28;
      5'b11101:
        casez_tmp_104 = rob_val_2_29;
      5'b11110:
        casez_tmp_104 = rob_val_2_30;
      default:
        casez_tmp_104 = rob_val_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_105 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_105 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_105 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_105 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_105 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_105 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_105 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_105 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_105 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_105 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_105 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_105 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_105 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_105 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_105 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_105 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_105 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_105 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_105 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_105 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_105 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_105 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_105 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_105 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_105 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_105 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_105 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_105 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_105 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_105 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_105 = rob_bsy_2_30;
      default:
        casez_tmp_105 = rob_bsy_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_106 = rob_val_2_0;
      5'b00001:
        casez_tmp_106 = rob_val_2_1;
      5'b00010:
        casez_tmp_106 = rob_val_2_2;
      5'b00011:
        casez_tmp_106 = rob_val_2_3;
      5'b00100:
        casez_tmp_106 = rob_val_2_4;
      5'b00101:
        casez_tmp_106 = rob_val_2_5;
      5'b00110:
        casez_tmp_106 = rob_val_2_6;
      5'b00111:
        casez_tmp_106 = rob_val_2_7;
      5'b01000:
        casez_tmp_106 = rob_val_2_8;
      5'b01001:
        casez_tmp_106 = rob_val_2_9;
      5'b01010:
        casez_tmp_106 = rob_val_2_10;
      5'b01011:
        casez_tmp_106 = rob_val_2_11;
      5'b01100:
        casez_tmp_106 = rob_val_2_12;
      5'b01101:
        casez_tmp_106 = rob_val_2_13;
      5'b01110:
        casez_tmp_106 = rob_val_2_14;
      5'b01111:
        casez_tmp_106 = rob_val_2_15;
      5'b10000:
        casez_tmp_106 = rob_val_2_16;
      5'b10001:
        casez_tmp_106 = rob_val_2_17;
      5'b10010:
        casez_tmp_106 = rob_val_2_18;
      5'b10011:
        casez_tmp_106 = rob_val_2_19;
      5'b10100:
        casez_tmp_106 = rob_val_2_20;
      5'b10101:
        casez_tmp_106 = rob_val_2_21;
      5'b10110:
        casez_tmp_106 = rob_val_2_22;
      5'b10111:
        casez_tmp_106 = rob_val_2_23;
      5'b11000:
        casez_tmp_106 = rob_val_2_24;
      5'b11001:
        casez_tmp_106 = rob_val_2_25;
      5'b11010:
        casez_tmp_106 = rob_val_2_26;
      5'b11011:
        casez_tmp_106 = rob_val_2_27;
      5'b11100:
        casez_tmp_106 = rob_val_2_28;
      5'b11101:
        casez_tmp_106 = rob_val_2_29;
      5'b11110:
        casez_tmp_106 = rob_val_2_30;
      default:
        casez_tmp_106 = rob_val_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_107 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_107 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_107 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_107 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_107 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_107 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_107 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_107 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_107 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_107 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_107 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_107 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_107 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_107 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_107 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_107 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_107 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_107 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_107 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_107 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_107 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_107 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_107 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_107 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_107 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_107 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_107 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_107 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_107 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_107 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_107 = rob_bsy_2_30;
      default:
        casez_tmp_107 = rob_bsy_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_2)
      5'b00000:
        casez_tmp_108 = rob_unsafe_2_0;
      5'b00001:
        casez_tmp_108 = rob_unsafe_2_1;
      5'b00010:
        casez_tmp_108 = rob_unsafe_2_2;
      5'b00011:
        casez_tmp_108 = rob_unsafe_2_3;
      5'b00100:
        casez_tmp_108 = rob_unsafe_2_4;
      5'b00101:
        casez_tmp_108 = rob_unsafe_2_5;
      5'b00110:
        casez_tmp_108 = rob_unsafe_2_6;
      5'b00111:
        casez_tmp_108 = rob_unsafe_2_7;
      5'b01000:
        casez_tmp_108 = rob_unsafe_2_8;
      5'b01001:
        casez_tmp_108 = rob_unsafe_2_9;
      5'b01010:
        casez_tmp_108 = rob_unsafe_2_10;
      5'b01011:
        casez_tmp_108 = rob_unsafe_2_11;
      5'b01100:
        casez_tmp_108 = rob_unsafe_2_12;
      5'b01101:
        casez_tmp_108 = rob_unsafe_2_13;
      5'b01110:
        casez_tmp_108 = rob_unsafe_2_14;
      5'b01111:
        casez_tmp_108 = rob_unsafe_2_15;
      5'b10000:
        casez_tmp_108 = rob_unsafe_2_16;
      5'b10001:
        casez_tmp_108 = rob_unsafe_2_17;
      5'b10010:
        casez_tmp_108 = rob_unsafe_2_18;
      5'b10011:
        casez_tmp_108 = rob_unsafe_2_19;
      5'b10100:
        casez_tmp_108 = rob_unsafe_2_20;
      5'b10101:
        casez_tmp_108 = rob_unsafe_2_21;
      5'b10110:
        casez_tmp_108 = rob_unsafe_2_22;
      5'b10111:
        casez_tmp_108 = rob_unsafe_2_23;
      5'b11000:
        casez_tmp_108 = rob_unsafe_2_24;
      5'b11001:
        casez_tmp_108 = rob_unsafe_2_25;
      5'b11010:
        casez_tmp_108 = rob_unsafe_2_26;
      5'b11011:
        casez_tmp_108 = rob_unsafe_2_27;
      5'b11100:
        casez_tmp_108 = rob_unsafe_2_28;
      5'b11101:
        casez_tmp_108 = rob_unsafe_2_29;
      5'b11110:
        casez_tmp_108 = rob_unsafe_2_30;
      default:
        casez_tmp_108 = rob_unsafe_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_109 = rob_unsafe_2_0;
      5'b00001:
        casez_tmp_109 = rob_unsafe_2_1;
      5'b00010:
        casez_tmp_109 = rob_unsafe_2_2;
      5'b00011:
        casez_tmp_109 = rob_unsafe_2_3;
      5'b00100:
        casez_tmp_109 = rob_unsafe_2_4;
      5'b00101:
        casez_tmp_109 = rob_unsafe_2_5;
      5'b00110:
        casez_tmp_109 = rob_unsafe_2_6;
      5'b00111:
        casez_tmp_109 = rob_unsafe_2_7;
      5'b01000:
        casez_tmp_109 = rob_unsafe_2_8;
      5'b01001:
        casez_tmp_109 = rob_unsafe_2_9;
      5'b01010:
        casez_tmp_109 = rob_unsafe_2_10;
      5'b01011:
        casez_tmp_109 = rob_unsafe_2_11;
      5'b01100:
        casez_tmp_109 = rob_unsafe_2_12;
      5'b01101:
        casez_tmp_109 = rob_unsafe_2_13;
      5'b01110:
        casez_tmp_109 = rob_unsafe_2_14;
      5'b01111:
        casez_tmp_109 = rob_unsafe_2_15;
      5'b10000:
        casez_tmp_109 = rob_unsafe_2_16;
      5'b10001:
        casez_tmp_109 = rob_unsafe_2_17;
      5'b10010:
        casez_tmp_109 = rob_unsafe_2_18;
      5'b10011:
        casez_tmp_109 = rob_unsafe_2_19;
      5'b10100:
        casez_tmp_109 = rob_unsafe_2_20;
      5'b10101:
        casez_tmp_109 = rob_unsafe_2_21;
      5'b10110:
        casez_tmp_109 = rob_unsafe_2_22;
      5'b10111:
        casez_tmp_109 = rob_unsafe_2_23;
      5'b11000:
        casez_tmp_109 = rob_unsafe_2_24;
      5'b11001:
        casez_tmp_109 = rob_unsafe_2_25;
      5'b11010:
        casez_tmp_109 = rob_unsafe_2_26;
      5'b11011:
        casez_tmp_109 = rob_unsafe_2_27;
      5'b11100:
        casez_tmp_109 = rob_unsafe_2_28;
      5'b11101:
        casez_tmp_109 = rob_unsafe_2_29;
      5'b11110:
        casez_tmp_109 = rob_unsafe_2_30;
      default:
        casez_tmp_109 = rob_unsafe_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_110 = rob_exception_2_0;
      5'b00001:
        casez_tmp_110 = rob_exception_2_1;
      5'b00010:
        casez_tmp_110 = rob_exception_2_2;
      5'b00011:
        casez_tmp_110 = rob_exception_2_3;
      5'b00100:
        casez_tmp_110 = rob_exception_2_4;
      5'b00101:
        casez_tmp_110 = rob_exception_2_5;
      5'b00110:
        casez_tmp_110 = rob_exception_2_6;
      5'b00111:
        casez_tmp_110 = rob_exception_2_7;
      5'b01000:
        casez_tmp_110 = rob_exception_2_8;
      5'b01001:
        casez_tmp_110 = rob_exception_2_9;
      5'b01010:
        casez_tmp_110 = rob_exception_2_10;
      5'b01011:
        casez_tmp_110 = rob_exception_2_11;
      5'b01100:
        casez_tmp_110 = rob_exception_2_12;
      5'b01101:
        casez_tmp_110 = rob_exception_2_13;
      5'b01110:
        casez_tmp_110 = rob_exception_2_14;
      5'b01111:
        casez_tmp_110 = rob_exception_2_15;
      5'b10000:
        casez_tmp_110 = rob_exception_2_16;
      5'b10001:
        casez_tmp_110 = rob_exception_2_17;
      5'b10010:
        casez_tmp_110 = rob_exception_2_18;
      5'b10011:
        casez_tmp_110 = rob_exception_2_19;
      5'b10100:
        casez_tmp_110 = rob_exception_2_20;
      5'b10101:
        casez_tmp_110 = rob_exception_2_21;
      5'b10110:
        casez_tmp_110 = rob_exception_2_22;
      5'b10111:
        casez_tmp_110 = rob_exception_2_23;
      5'b11000:
        casez_tmp_110 = rob_exception_2_24;
      5'b11001:
        casez_tmp_110 = rob_exception_2_25;
      5'b11010:
        casez_tmp_110 = rob_exception_2_26;
      5'b11011:
        casez_tmp_110 = rob_exception_2_27;
      5'b11100:
        casez_tmp_110 = rob_exception_2_28;
      5'b11101:
        casez_tmp_110 = rob_exception_2_29;
      5'b11110:
        casez_tmp_110 = rob_exception_2_30;
      default:
        casez_tmp_110 = rob_exception_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_111 = rob_val_2_0;
      5'b00001:
        casez_tmp_111 = rob_val_2_1;
      5'b00010:
        casez_tmp_111 = rob_val_2_2;
      5'b00011:
        casez_tmp_111 = rob_val_2_3;
      5'b00100:
        casez_tmp_111 = rob_val_2_4;
      5'b00101:
        casez_tmp_111 = rob_val_2_5;
      5'b00110:
        casez_tmp_111 = rob_val_2_6;
      5'b00111:
        casez_tmp_111 = rob_val_2_7;
      5'b01000:
        casez_tmp_111 = rob_val_2_8;
      5'b01001:
        casez_tmp_111 = rob_val_2_9;
      5'b01010:
        casez_tmp_111 = rob_val_2_10;
      5'b01011:
        casez_tmp_111 = rob_val_2_11;
      5'b01100:
        casez_tmp_111 = rob_val_2_12;
      5'b01101:
        casez_tmp_111 = rob_val_2_13;
      5'b01110:
        casez_tmp_111 = rob_val_2_14;
      5'b01111:
        casez_tmp_111 = rob_val_2_15;
      5'b10000:
        casez_tmp_111 = rob_val_2_16;
      5'b10001:
        casez_tmp_111 = rob_val_2_17;
      5'b10010:
        casez_tmp_111 = rob_val_2_18;
      5'b10011:
        casez_tmp_111 = rob_val_2_19;
      5'b10100:
        casez_tmp_111 = rob_val_2_20;
      5'b10101:
        casez_tmp_111 = rob_val_2_21;
      5'b10110:
        casez_tmp_111 = rob_val_2_22;
      5'b10111:
        casez_tmp_111 = rob_val_2_23;
      5'b11000:
        casez_tmp_111 = rob_val_2_24;
      5'b11001:
        casez_tmp_111 = rob_val_2_25;
      5'b11010:
        casez_tmp_111 = rob_val_2_26;
      5'b11011:
        casez_tmp_111 = rob_val_2_27;
      5'b11100:
        casez_tmp_111 = rob_val_2_28;
      5'b11101:
        casez_tmp_111 = rob_val_2_29;
      5'b11110:
        casez_tmp_111 = rob_val_2_30;
      default:
        casez_tmp_111 = rob_val_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_112 = rob_val_2_0;
      5'b00001:
        casez_tmp_112 = rob_val_2_1;
      5'b00010:
        casez_tmp_112 = rob_val_2_2;
      5'b00011:
        casez_tmp_112 = rob_val_2_3;
      5'b00100:
        casez_tmp_112 = rob_val_2_4;
      5'b00101:
        casez_tmp_112 = rob_val_2_5;
      5'b00110:
        casez_tmp_112 = rob_val_2_6;
      5'b00111:
        casez_tmp_112 = rob_val_2_7;
      5'b01000:
        casez_tmp_112 = rob_val_2_8;
      5'b01001:
        casez_tmp_112 = rob_val_2_9;
      5'b01010:
        casez_tmp_112 = rob_val_2_10;
      5'b01011:
        casez_tmp_112 = rob_val_2_11;
      5'b01100:
        casez_tmp_112 = rob_val_2_12;
      5'b01101:
        casez_tmp_112 = rob_val_2_13;
      5'b01110:
        casez_tmp_112 = rob_val_2_14;
      5'b01111:
        casez_tmp_112 = rob_val_2_15;
      5'b10000:
        casez_tmp_112 = rob_val_2_16;
      5'b10001:
        casez_tmp_112 = rob_val_2_17;
      5'b10010:
        casez_tmp_112 = rob_val_2_18;
      5'b10011:
        casez_tmp_112 = rob_val_2_19;
      5'b10100:
        casez_tmp_112 = rob_val_2_20;
      5'b10101:
        casez_tmp_112 = rob_val_2_21;
      5'b10110:
        casez_tmp_112 = rob_val_2_22;
      5'b10111:
        casez_tmp_112 = rob_val_2_23;
      5'b11000:
        casez_tmp_112 = rob_val_2_24;
      5'b11001:
        casez_tmp_112 = rob_val_2_25;
      5'b11010:
        casez_tmp_112 = rob_val_2_26;
      5'b11011:
        casez_tmp_112 = rob_val_2_27;
      5'b11100:
        casez_tmp_112 = rob_val_2_28;
      5'b11101:
        casez_tmp_112 = rob_val_2_29;
      5'b11110:
        casez_tmp_112 = rob_val_2_30;
      default:
        casez_tmp_112 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1917 = _GEN_1375 & ~casez_tmp_112;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_113 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_113 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_113 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_113 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_113 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_113 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_113 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_113 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_113 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_113 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_113 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_113 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_113 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_113 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_113 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_113 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_113 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_113 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_113 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_113 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_113 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_113 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_113 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_113 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_113 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_113 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_113 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_113 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_113 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_113 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_113 = rob_bsy_2_30;
      default:
        casez_tmp_113 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1918 = _GEN_1375 & ~casez_tmp_113;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_114 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_114 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_114 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_114 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_114 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_114 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_114 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_114 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_114 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_114 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_114 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_114 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_114 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_114 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_114 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_114 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_114 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_114 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_114 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_114 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_114 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_114 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_114 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_114 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_114 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_114 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_114 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_114 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_114 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_114 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_114 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_114 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_115 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_115 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_115 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_115 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_115 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_115 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_115 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_115 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_115 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_115 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_115 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_115 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_115 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_115 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_115 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_115 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_115 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_115 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_115 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_115 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_115 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_115 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_115 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_115 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_115 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_115 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_115 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_115 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_115 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_115 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_115 = rob_uop_2_30_pdst;
      default:
        casez_tmp_115 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1919 = _GEN_1375 & casez_tmp_114 & casez_tmp_115 != io_wb_resps_0_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_116 = rob_val_2_0;
      5'b00001:
        casez_tmp_116 = rob_val_2_1;
      5'b00010:
        casez_tmp_116 = rob_val_2_2;
      5'b00011:
        casez_tmp_116 = rob_val_2_3;
      5'b00100:
        casez_tmp_116 = rob_val_2_4;
      5'b00101:
        casez_tmp_116 = rob_val_2_5;
      5'b00110:
        casez_tmp_116 = rob_val_2_6;
      5'b00111:
        casez_tmp_116 = rob_val_2_7;
      5'b01000:
        casez_tmp_116 = rob_val_2_8;
      5'b01001:
        casez_tmp_116 = rob_val_2_9;
      5'b01010:
        casez_tmp_116 = rob_val_2_10;
      5'b01011:
        casez_tmp_116 = rob_val_2_11;
      5'b01100:
        casez_tmp_116 = rob_val_2_12;
      5'b01101:
        casez_tmp_116 = rob_val_2_13;
      5'b01110:
        casez_tmp_116 = rob_val_2_14;
      5'b01111:
        casez_tmp_116 = rob_val_2_15;
      5'b10000:
        casez_tmp_116 = rob_val_2_16;
      5'b10001:
        casez_tmp_116 = rob_val_2_17;
      5'b10010:
        casez_tmp_116 = rob_val_2_18;
      5'b10011:
        casez_tmp_116 = rob_val_2_19;
      5'b10100:
        casez_tmp_116 = rob_val_2_20;
      5'b10101:
        casez_tmp_116 = rob_val_2_21;
      5'b10110:
        casez_tmp_116 = rob_val_2_22;
      5'b10111:
        casez_tmp_116 = rob_val_2_23;
      5'b11000:
        casez_tmp_116 = rob_val_2_24;
      5'b11001:
        casez_tmp_116 = rob_val_2_25;
      5'b11010:
        casez_tmp_116 = rob_val_2_26;
      5'b11011:
        casez_tmp_116 = rob_val_2_27;
      5'b11100:
        casez_tmp_116 = rob_val_2_28;
      5'b11101:
        casez_tmp_116 = rob_val_2_29;
      5'b11110:
        casez_tmp_116 = rob_val_2_30;
      default:
        casez_tmp_116 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1920 = _GEN_926 & ~casez_tmp_116;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_117 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_117 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_117 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_117 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_117 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_117 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_117 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_117 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_117 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_117 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_117 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_117 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_117 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_117 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_117 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_117 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_117 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_117 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_117 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_117 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_117 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_117 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_117 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_117 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_117 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_117 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_117 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_117 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_117 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_117 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_117 = rob_bsy_2_30;
      default:
        casez_tmp_117 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1921 = _GEN_926 & ~casez_tmp_117;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_118 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_118 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_118 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_118 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_118 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_118 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_118 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_118 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_118 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_118 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_118 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_118 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_118 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_118 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_118 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_118 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_118 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_118 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_118 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_118 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_118 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_118 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_118 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_118 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_118 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_118 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_118 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_118 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_118 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_118 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_118 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_118 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_119 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_119 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_119 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_119 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_119 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_119 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_119 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_119 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_119 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_119 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_119 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_119 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_119 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_119 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_119 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_119 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_119 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_119 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_119 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_119 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_119 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_119 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_119 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_119 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_119 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_119 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_119 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_119 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_119 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_119 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_119 = rob_uop_2_30_pdst;
      default:
        casez_tmp_119 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1922 = _GEN_926 & casez_tmp_118 & casez_tmp_119 != io_wb_resps_1_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_120 = rob_val_2_0;
      5'b00001:
        casez_tmp_120 = rob_val_2_1;
      5'b00010:
        casez_tmp_120 = rob_val_2_2;
      5'b00011:
        casez_tmp_120 = rob_val_2_3;
      5'b00100:
        casez_tmp_120 = rob_val_2_4;
      5'b00101:
        casez_tmp_120 = rob_val_2_5;
      5'b00110:
        casez_tmp_120 = rob_val_2_6;
      5'b00111:
        casez_tmp_120 = rob_val_2_7;
      5'b01000:
        casez_tmp_120 = rob_val_2_8;
      5'b01001:
        casez_tmp_120 = rob_val_2_9;
      5'b01010:
        casez_tmp_120 = rob_val_2_10;
      5'b01011:
        casez_tmp_120 = rob_val_2_11;
      5'b01100:
        casez_tmp_120 = rob_val_2_12;
      5'b01101:
        casez_tmp_120 = rob_val_2_13;
      5'b01110:
        casez_tmp_120 = rob_val_2_14;
      5'b01111:
        casez_tmp_120 = rob_val_2_15;
      5'b10000:
        casez_tmp_120 = rob_val_2_16;
      5'b10001:
        casez_tmp_120 = rob_val_2_17;
      5'b10010:
        casez_tmp_120 = rob_val_2_18;
      5'b10011:
        casez_tmp_120 = rob_val_2_19;
      5'b10100:
        casez_tmp_120 = rob_val_2_20;
      5'b10101:
        casez_tmp_120 = rob_val_2_21;
      5'b10110:
        casez_tmp_120 = rob_val_2_22;
      5'b10111:
        casez_tmp_120 = rob_val_2_23;
      5'b11000:
        casez_tmp_120 = rob_val_2_24;
      5'b11001:
        casez_tmp_120 = rob_val_2_25;
      5'b11010:
        casez_tmp_120 = rob_val_2_26;
      5'b11011:
        casez_tmp_120 = rob_val_2_27;
      5'b11100:
        casez_tmp_120 = rob_val_2_28;
      5'b11101:
        casez_tmp_120 = rob_val_2_29;
      5'b11110:
        casez_tmp_120 = rob_val_2_30;
      default:
        casez_tmp_120 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1923 = _GEN_1376 & ~casez_tmp_120;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_121 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_121 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_121 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_121 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_121 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_121 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_121 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_121 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_121 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_121 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_121 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_121 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_121 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_121 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_121 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_121 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_121 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_121 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_121 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_121 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_121 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_121 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_121 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_121 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_121 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_121 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_121 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_121 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_121 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_121 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_121 = rob_bsy_2_30;
      default:
        casez_tmp_121 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1924 = _GEN_1376 & ~casez_tmp_121;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_122 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_122 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_122 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_122 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_122 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_122 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_122 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_122 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_122 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_122 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_122 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_122 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_122 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_122 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_122 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_122 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_122 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_122 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_122 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_122 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_122 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_122 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_122 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_122 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_122 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_122 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_122 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_122 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_122 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_122 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_122 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_122 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_123 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_123 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_123 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_123 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_123 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_123 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_123 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_123 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_123 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_123 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_123 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_123 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_123 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_123 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_123 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_123 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_123 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_123 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_123 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_123 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_123 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_123 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_123 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_123 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_123 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_123 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_123 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_123 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_123 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_123 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_123 = rob_uop_2_30_pdst;
      default:
        casez_tmp_123 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1925 = _GEN_1376 & casez_tmp_122 & casez_tmp_123 != io_wb_resps_2_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_124 = rob_val_2_0;
      5'b00001:
        casez_tmp_124 = rob_val_2_1;
      5'b00010:
        casez_tmp_124 = rob_val_2_2;
      5'b00011:
        casez_tmp_124 = rob_val_2_3;
      5'b00100:
        casez_tmp_124 = rob_val_2_4;
      5'b00101:
        casez_tmp_124 = rob_val_2_5;
      5'b00110:
        casez_tmp_124 = rob_val_2_6;
      5'b00111:
        casez_tmp_124 = rob_val_2_7;
      5'b01000:
        casez_tmp_124 = rob_val_2_8;
      5'b01001:
        casez_tmp_124 = rob_val_2_9;
      5'b01010:
        casez_tmp_124 = rob_val_2_10;
      5'b01011:
        casez_tmp_124 = rob_val_2_11;
      5'b01100:
        casez_tmp_124 = rob_val_2_12;
      5'b01101:
        casez_tmp_124 = rob_val_2_13;
      5'b01110:
        casez_tmp_124 = rob_val_2_14;
      5'b01111:
        casez_tmp_124 = rob_val_2_15;
      5'b10000:
        casez_tmp_124 = rob_val_2_16;
      5'b10001:
        casez_tmp_124 = rob_val_2_17;
      5'b10010:
        casez_tmp_124 = rob_val_2_18;
      5'b10011:
        casez_tmp_124 = rob_val_2_19;
      5'b10100:
        casez_tmp_124 = rob_val_2_20;
      5'b10101:
        casez_tmp_124 = rob_val_2_21;
      5'b10110:
        casez_tmp_124 = rob_val_2_22;
      5'b10111:
        casez_tmp_124 = rob_val_2_23;
      5'b11000:
        casez_tmp_124 = rob_val_2_24;
      5'b11001:
        casez_tmp_124 = rob_val_2_25;
      5'b11010:
        casez_tmp_124 = rob_val_2_26;
      5'b11011:
        casez_tmp_124 = rob_val_2_27;
      5'b11100:
        casez_tmp_124 = rob_val_2_28;
      5'b11101:
        casez_tmp_124 = rob_val_2_29;
      5'b11110:
        casez_tmp_124 = rob_val_2_30;
      default:
        casez_tmp_124 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1926 = _GEN_925 & ~casez_tmp_124;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_125 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_125 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_125 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_125 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_125 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_125 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_125 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_125 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_125 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_125 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_125 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_125 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_125 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_125 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_125 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_125 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_125 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_125 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_125 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_125 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_125 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_125 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_125 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_125 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_125 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_125 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_125 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_125 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_125 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_125 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_125 = rob_bsy_2_30;
      default:
        casez_tmp_125 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1927 = _GEN_925 & ~casez_tmp_125;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_126 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_126 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_126 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_126 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_126 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_126 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_126 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_126 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_126 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_126 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_126 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_126 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_126 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_126 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_126 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_126 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_126 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_126 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_126 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_126 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_126 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_126 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_126 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_126 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_126 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_126 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_126 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_126 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_126 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_126 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_126 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_126 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_127 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_127 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_127 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_127 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_127 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_127 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_127 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_127 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_127 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_127 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_127 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_127 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_127 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_127 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_127 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_127 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_127 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_127 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_127 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_127 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_127 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_127 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_127 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_127 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_127 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_127 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_127 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_127 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_127 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_127 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_127 = rob_uop_2_30_pdst;
      default:
        casez_tmp_127 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1928 = _GEN_925 & casez_tmp_126 & casez_tmp_127 != io_wb_resps_3_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_128 = rob_val_2_0;
      5'b00001:
        casez_tmp_128 = rob_val_2_1;
      5'b00010:
        casez_tmp_128 = rob_val_2_2;
      5'b00011:
        casez_tmp_128 = rob_val_2_3;
      5'b00100:
        casez_tmp_128 = rob_val_2_4;
      5'b00101:
        casez_tmp_128 = rob_val_2_5;
      5'b00110:
        casez_tmp_128 = rob_val_2_6;
      5'b00111:
        casez_tmp_128 = rob_val_2_7;
      5'b01000:
        casez_tmp_128 = rob_val_2_8;
      5'b01001:
        casez_tmp_128 = rob_val_2_9;
      5'b01010:
        casez_tmp_128 = rob_val_2_10;
      5'b01011:
        casez_tmp_128 = rob_val_2_11;
      5'b01100:
        casez_tmp_128 = rob_val_2_12;
      5'b01101:
        casez_tmp_128 = rob_val_2_13;
      5'b01110:
        casez_tmp_128 = rob_val_2_14;
      5'b01111:
        casez_tmp_128 = rob_val_2_15;
      5'b10000:
        casez_tmp_128 = rob_val_2_16;
      5'b10001:
        casez_tmp_128 = rob_val_2_17;
      5'b10010:
        casez_tmp_128 = rob_val_2_18;
      5'b10011:
        casez_tmp_128 = rob_val_2_19;
      5'b10100:
        casez_tmp_128 = rob_val_2_20;
      5'b10101:
        casez_tmp_128 = rob_val_2_21;
      5'b10110:
        casez_tmp_128 = rob_val_2_22;
      5'b10111:
        casez_tmp_128 = rob_val_2_23;
      5'b11000:
        casez_tmp_128 = rob_val_2_24;
      5'b11001:
        casez_tmp_128 = rob_val_2_25;
      5'b11010:
        casez_tmp_128 = rob_val_2_26;
      5'b11011:
        casez_tmp_128 = rob_val_2_27;
      5'b11100:
        casez_tmp_128 = rob_val_2_28;
      5'b11101:
        casez_tmp_128 = rob_val_2_29;
      5'b11110:
        casez_tmp_128 = rob_val_2_30;
      default:
        casez_tmp_128 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1929 = _GEN_1377 & ~casez_tmp_128;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_129 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_129 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_129 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_129 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_129 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_129 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_129 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_129 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_129 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_129 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_129 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_129 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_129 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_129 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_129 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_129 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_129 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_129 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_129 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_129 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_129 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_129 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_129 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_129 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_129 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_129 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_129 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_129 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_129 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_129 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_129 = rob_bsy_2_30;
      default:
        casez_tmp_129 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1930 = _GEN_1377 & ~casez_tmp_129;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_130 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_130 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_130 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_130 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_130 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_130 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_130 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_130 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_130 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_130 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_130 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_130 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_130 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_130 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_130 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_130 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_130 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_130 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_130 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_130 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_130 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_130 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_130 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_130 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_130 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_130 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_130 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_130 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_130 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_130 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_130 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_130 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_131 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_131 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_131 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_131 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_131 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_131 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_131 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_131 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_131 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_131 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_131 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_131 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_131 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_131 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_131 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_131 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_131 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_131 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_131 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_131 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_131 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_131 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_131 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_131 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_131 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_131 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_131 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_131 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_131 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_131 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_131 = rob_uop_2_30_pdst;
      default:
        casez_tmp_131 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1931 = _GEN_1377 & casez_tmp_130 & casez_tmp_131 != io_wb_resps_4_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_132 = rob_val_2_0;
      5'b00001:
        casez_tmp_132 = rob_val_2_1;
      5'b00010:
        casez_tmp_132 = rob_val_2_2;
      5'b00011:
        casez_tmp_132 = rob_val_2_3;
      5'b00100:
        casez_tmp_132 = rob_val_2_4;
      5'b00101:
        casez_tmp_132 = rob_val_2_5;
      5'b00110:
        casez_tmp_132 = rob_val_2_6;
      5'b00111:
        casez_tmp_132 = rob_val_2_7;
      5'b01000:
        casez_tmp_132 = rob_val_2_8;
      5'b01001:
        casez_tmp_132 = rob_val_2_9;
      5'b01010:
        casez_tmp_132 = rob_val_2_10;
      5'b01011:
        casez_tmp_132 = rob_val_2_11;
      5'b01100:
        casez_tmp_132 = rob_val_2_12;
      5'b01101:
        casez_tmp_132 = rob_val_2_13;
      5'b01110:
        casez_tmp_132 = rob_val_2_14;
      5'b01111:
        casez_tmp_132 = rob_val_2_15;
      5'b10000:
        casez_tmp_132 = rob_val_2_16;
      5'b10001:
        casez_tmp_132 = rob_val_2_17;
      5'b10010:
        casez_tmp_132 = rob_val_2_18;
      5'b10011:
        casez_tmp_132 = rob_val_2_19;
      5'b10100:
        casez_tmp_132 = rob_val_2_20;
      5'b10101:
        casez_tmp_132 = rob_val_2_21;
      5'b10110:
        casez_tmp_132 = rob_val_2_22;
      5'b10111:
        casez_tmp_132 = rob_val_2_23;
      5'b11000:
        casez_tmp_132 = rob_val_2_24;
      5'b11001:
        casez_tmp_132 = rob_val_2_25;
      5'b11010:
        casez_tmp_132 = rob_val_2_26;
      5'b11011:
        casez_tmp_132 = rob_val_2_27;
      5'b11100:
        casez_tmp_132 = rob_val_2_28;
      5'b11101:
        casez_tmp_132 = rob_val_2_29;
      5'b11110:
        casez_tmp_132 = rob_val_2_30;
      default:
        casez_tmp_132 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1932 = _GEN_924 & ~casez_tmp_132;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_133 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_133 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_133 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_133 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_133 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_133 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_133 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_133 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_133 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_133 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_133 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_133 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_133 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_133 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_133 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_133 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_133 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_133 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_133 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_133 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_133 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_133 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_133 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_133 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_133 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_133 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_133 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_133 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_133 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_133 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_133 = rob_bsy_2_30;
      default:
        casez_tmp_133 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1933 = _GEN_924 & ~casez_tmp_133;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_134 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_134 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_134 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_134 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_134 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_134 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_134 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_134 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_134 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_134 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_134 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_134 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_134 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_134 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_134 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_134 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_134 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_134 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_134 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_134 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_134 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_134 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_134 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_134 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_134 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_134 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_134 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_134 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_134 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_134 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_134 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_134 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_135 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_135 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_135 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_135 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_135 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_135 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_135 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_135 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_135 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_135 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_135 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_135 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_135 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_135 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_135 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_135 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_135 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_135 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_135 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_135 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_135 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_135 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_135 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_135 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_135 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_135 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_135 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_135 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_135 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_135 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_135 = rob_uop_2_30_pdst;
      default:
        casez_tmp_135 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1934 = _GEN_924 & casez_tmp_134 & casez_tmp_135 != io_wb_resps_5_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_136 = rob_val_2_0;
      5'b00001:
        casez_tmp_136 = rob_val_2_1;
      5'b00010:
        casez_tmp_136 = rob_val_2_2;
      5'b00011:
        casez_tmp_136 = rob_val_2_3;
      5'b00100:
        casez_tmp_136 = rob_val_2_4;
      5'b00101:
        casez_tmp_136 = rob_val_2_5;
      5'b00110:
        casez_tmp_136 = rob_val_2_6;
      5'b00111:
        casez_tmp_136 = rob_val_2_7;
      5'b01000:
        casez_tmp_136 = rob_val_2_8;
      5'b01001:
        casez_tmp_136 = rob_val_2_9;
      5'b01010:
        casez_tmp_136 = rob_val_2_10;
      5'b01011:
        casez_tmp_136 = rob_val_2_11;
      5'b01100:
        casez_tmp_136 = rob_val_2_12;
      5'b01101:
        casez_tmp_136 = rob_val_2_13;
      5'b01110:
        casez_tmp_136 = rob_val_2_14;
      5'b01111:
        casez_tmp_136 = rob_val_2_15;
      5'b10000:
        casez_tmp_136 = rob_val_2_16;
      5'b10001:
        casez_tmp_136 = rob_val_2_17;
      5'b10010:
        casez_tmp_136 = rob_val_2_18;
      5'b10011:
        casez_tmp_136 = rob_val_2_19;
      5'b10100:
        casez_tmp_136 = rob_val_2_20;
      5'b10101:
        casez_tmp_136 = rob_val_2_21;
      5'b10110:
        casez_tmp_136 = rob_val_2_22;
      5'b10111:
        casez_tmp_136 = rob_val_2_23;
      5'b11000:
        casez_tmp_136 = rob_val_2_24;
      5'b11001:
        casez_tmp_136 = rob_val_2_25;
      5'b11010:
        casez_tmp_136 = rob_val_2_26;
      5'b11011:
        casez_tmp_136 = rob_val_2_27;
      5'b11100:
        casez_tmp_136 = rob_val_2_28;
      5'b11101:
        casez_tmp_136 = rob_val_2_29;
      5'b11110:
        casez_tmp_136 = rob_val_2_30;
      default:
        casez_tmp_136 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1935 = _GEN_1378 & ~casez_tmp_136;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_137 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_137 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_137 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_137 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_137 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_137 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_137 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_137 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_137 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_137 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_137 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_137 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_137 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_137 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_137 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_137 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_137 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_137 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_137 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_137 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_137 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_137 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_137 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_137 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_137 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_137 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_137 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_137 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_137 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_137 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_137 = rob_bsy_2_30;
      default:
        casez_tmp_137 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1936 = _GEN_1378 & ~casez_tmp_137;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_138 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_138 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_138 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_138 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_138 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_138 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_138 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_138 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_138 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_138 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_138 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_138 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_138 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_138 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_138 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_138 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_138 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_138 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_138 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_138 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_138 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_138 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_138 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_138 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_138 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_138 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_138 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_138 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_138 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_138 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_138 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_138 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_139 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_139 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_139 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_139 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_139 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_139 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_139 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_139 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_139 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_139 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_139 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_139 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_139 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_139 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_139 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_139 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_139 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_139 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_139 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_139 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_139 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_139 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_139 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_139 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_139 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_139 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_139 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_139 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_139 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_139 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_139 = rob_uop_2_30_pdst;
      default:
        casez_tmp_139 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1937 = _GEN_1378 & casez_tmp_138 & casez_tmp_139 != io_wb_resps_6_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_140 = rob_val_2_0;
      5'b00001:
        casez_tmp_140 = rob_val_2_1;
      5'b00010:
        casez_tmp_140 = rob_val_2_2;
      5'b00011:
        casez_tmp_140 = rob_val_2_3;
      5'b00100:
        casez_tmp_140 = rob_val_2_4;
      5'b00101:
        casez_tmp_140 = rob_val_2_5;
      5'b00110:
        casez_tmp_140 = rob_val_2_6;
      5'b00111:
        casez_tmp_140 = rob_val_2_7;
      5'b01000:
        casez_tmp_140 = rob_val_2_8;
      5'b01001:
        casez_tmp_140 = rob_val_2_9;
      5'b01010:
        casez_tmp_140 = rob_val_2_10;
      5'b01011:
        casez_tmp_140 = rob_val_2_11;
      5'b01100:
        casez_tmp_140 = rob_val_2_12;
      5'b01101:
        casez_tmp_140 = rob_val_2_13;
      5'b01110:
        casez_tmp_140 = rob_val_2_14;
      5'b01111:
        casez_tmp_140 = rob_val_2_15;
      5'b10000:
        casez_tmp_140 = rob_val_2_16;
      5'b10001:
        casez_tmp_140 = rob_val_2_17;
      5'b10010:
        casez_tmp_140 = rob_val_2_18;
      5'b10011:
        casez_tmp_140 = rob_val_2_19;
      5'b10100:
        casez_tmp_140 = rob_val_2_20;
      5'b10101:
        casez_tmp_140 = rob_val_2_21;
      5'b10110:
        casez_tmp_140 = rob_val_2_22;
      5'b10111:
        casez_tmp_140 = rob_val_2_23;
      5'b11000:
        casez_tmp_140 = rob_val_2_24;
      5'b11001:
        casez_tmp_140 = rob_val_2_25;
      5'b11010:
        casez_tmp_140 = rob_val_2_26;
      5'b11011:
        casez_tmp_140 = rob_val_2_27;
      5'b11100:
        casez_tmp_140 = rob_val_2_28;
      5'b11101:
        casez_tmp_140 = rob_val_2_29;
      5'b11110:
        casez_tmp_140 = rob_val_2_30;
      default:
        casez_tmp_140 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1938 = _GEN_923 & ~casez_tmp_140;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_141 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_141 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_141 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_141 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_141 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_141 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_141 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_141 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_141 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_141 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_141 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_141 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_141 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_141 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_141 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_141 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_141 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_141 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_141 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_141 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_141 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_141 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_141 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_141 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_141 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_141 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_141 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_141 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_141 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_141 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_141 = rob_bsy_2_30;
      default:
        casez_tmp_141 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1939 = _GEN_923 & ~casez_tmp_141;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_142 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_142 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_142 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_142 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_142 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_142 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_142 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_142 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_142 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_142 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_142 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_142 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_142 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_142 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_142 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_142 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_142 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_142 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_142 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_142 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_142 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_142 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_142 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_142 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_142 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_142 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_142 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_142 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_142 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_142 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_142 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_142 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_143 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_143 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_143 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_143 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_143 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_143 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_143 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_143 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_143 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_143 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_143 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_143 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_143 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_143 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_143 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_143 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_143 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_143 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_143 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_143 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_143 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_143 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_143 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_143 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_143 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_143 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_143 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_143 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_143 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_143 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_143 = rob_uop_2_30_pdst;
      default:
        casez_tmp_143 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1940 = _GEN_923 & casez_tmp_142 & casez_tmp_143 != io_wb_resps_7_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_144 = rob_val_2_0;
      5'b00001:
        casez_tmp_144 = rob_val_2_1;
      5'b00010:
        casez_tmp_144 = rob_val_2_2;
      5'b00011:
        casez_tmp_144 = rob_val_2_3;
      5'b00100:
        casez_tmp_144 = rob_val_2_4;
      5'b00101:
        casez_tmp_144 = rob_val_2_5;
      5'b00110:
        casez_tmp_144 = rob_val_2_6;
      5'b00111:
        casez_tmp_144 = rob_val_2_7;
      5'b01000:
        casez_tmp_144 = rob_val_2_8;
      5'b01001:
        casez_tmp_144 = rob_val_2_9;
      5'b01010:
        casez_tmp_144 = rob_val_2_10;
      5'b01011:
        casez_tmp_144 = rob_val_2_11;
      5'b01100:
        casez_tmp_144 = rob_val_2_12;
      5'b01101:
        casez_tmp_144 = rob_val_2_13;
      5'b01110:
        casez_tmp_144 = rob_val_2_14;
      5'b01111:
        casez_tmp_144 = rob_val_2_15;
      5'b10000:
        casez_tmp_144 = rob_val_2_16;
      5'b10001:
        casez_tmp_144 = rob_val_2_17;
      5'b10010:
        casez_tmp_144 = rob_val_2_18;
      5'b10011:
        casez_tmp_144 = rob_val_2_19;
      5'b10100:
        casez_tmp_144 = rob_val_2_20;
      5'b10101:
        casez_tmp_144 = rob_val_2_21;
      5'b10110:
        casez_tmp_144 = rob_val_2_22;
      5'b10111:
        casez_tmp_144 = rob_val_2_23;
      5'b11000:
        casez_tmp_144 = rob_val_2_24;
      5'b11001:
        casez_tmp_144 = rob_val_2_25;
      5'b11010:
        casez_tmp_144 = rob_val_2_26;
      5'b11011:
        casez_tmp_144 = rob_val_2_27;
      5'b11100:
        casez_tmp_144 = rob_val_2_28;
      5'b11101:
        casez_tmp_144 = rob_val_2_29;
      5'b11110:
        casez_tmp_144 = rob_val_2_30;
      default:
        casez_tmp_144 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1941 = _GEN_1379 & ~casez_tmp_144;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_145 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_145 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_145 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_145 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_145 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_145 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_145 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_145 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_145 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_145 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_145 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_145 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_145 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_145 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_145 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_145 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_145 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_145 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_145 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_145 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_145 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_145 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_145 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_145 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_145 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_145 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_145 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_145 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_145 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_145 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_145 = rob_bsy_2_30;
      default:
        casez_tmp_145 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1942 = _GEN_1379 & ~casez_tmp_145;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_146 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_146 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_146 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_146 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_146 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_146 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_146 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_146 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_146 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_146 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_146 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_146 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_146 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_146 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_146 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_146 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_146 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_146 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_146 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_146 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_146 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_146 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_146 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_146 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_146 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_146 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_146 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_146 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_146 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_146 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_146 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_146 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_147 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_147 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_147 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_147 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_147 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_147 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_147 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_147 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_147 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_147 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_147 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_147 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_147 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_147 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_147 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_147 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_147 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_147 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_147 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_147 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_147 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_147 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_147 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_147 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_147 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_147 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_147 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_147 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_147 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_147 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_147 = rob_uop_2_30_pdst;
      default:
        casez_tmp_147 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1943 = _GEN_1379 & casez_tmp_146 & casez_tmp_147 != io_wb_resps_8_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_148 = rob_val_2_0;
      5'b00001:
        casez_tmp_148 = rob_val_2_1;
      5'b00010:
        casez_tmp_148 = rob_val_2_2;
      5'b00011:
        casez_tmp_148 = rob_val_2_3;
      5'b00100:
        casez_tmp_148 = rob_val_2_4;
      5'b00101:
        casez_tmp_148 = rob_val_2_5;
      5'b00110:
        casez_tmp_148 = rob_val_2_6;
      5'b00111:
        casez_tmp_148 = rob_val_2_7;
      5'b01000:
        casez_tmp_148 = rob_val_2_8;
      5'b01001:
        casez_tmp_148 = rob_val_2_9;
      5'b01010:
        casez_tmp_148 = rob_val_2_10;
      5'b01011:
        casez_tmp_148 = rob_val_2_11;
      5'b01100:
        casez_tmp_148 = rob_val_2_12;
      5'b01101:
        casez_tmp_148 = rob_val_2_13;
      5'b01110:
        casez_tmp_148 = rob_val_2_14;
      5'b01111:
        casez_tmp_148 = rob_val_2_15;
      5'b10000:
        casez_tmp_148 = rob_val_2_16;
      5'b10001:
        casez_tmp_148 = rob_val_2_17;
      5'b10010:
        casez_tmp_148 = rob_val_2_18;
      5'b10011:
        casez_tmp_148 = rob_val_2_19;
      5'b10100:
        casez_tmp_148 = rob_val_2_20;
      5'b10101:
        casez_tmp_148 = rob_val_2_21;
      5'b10110:
        casez_tmp_148 = rob_val_2_22;
      5'b10111:
        casez_tmp_148 = rob_val_2_23;
      5'b11000:
        casez_tmp_148 = rob_val_2_24;
      5'b11001:
        casez_tmp_148 = rob_val_2_25;
      5'b11010:
        casez_tmp_148 = rob_val_2_26;
      5'b11011:
        casez_tmp_148 = rob_val_2_27;
      5'b11100:
        casez_tmp_148 = rob_val_2_28;
      5'b11101:
        casez_tmp_148 = rob_val_2_29;
      5'b11110:
        casez_tmp_148 = rob_val_2_30;
      default:
        casez_tmp_148 = rob_val_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1944 = _GEN_922 & ~casez_tmp_148;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_149 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_149 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_149 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_149 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_149 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_149 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_149 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_149 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_149 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_149 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_149 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_149 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_149 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_149 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_149 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_149 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_149 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_149 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_149 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_149 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_149 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_149 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_149 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_149 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_149 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_149 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_149 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_149 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_149 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_149 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_149 = rob_bsy_2_30;
      default:
        casez_tmp_149 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire       _GEN_1945 = _GEN_922 & ~casez_tmp_149;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_150 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_150 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_150 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_150 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_150 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_150 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_150 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_150 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_150 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_150 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_150 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_150 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_150 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_150 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_150 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_150 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_150 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_150 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_150 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_150 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_150 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_150 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_150 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_150 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_150 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_150 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_150 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_150 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_150 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_150 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_150 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_150 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_151 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_151 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_151 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_151 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_151 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_151 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_151 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_151 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_151 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_151 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_151 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_151 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_151 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_151 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_151 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_151 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_151 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_151 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_151 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_151 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_151 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_151 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_151 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_151 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_151 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_151 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_151 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_151 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_151 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_151 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_151 = rob_uop_2_30_pdst;
      default:
        casez_tmp_151 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1946 = _GEN_922 & casez_tmp_150 & casez_tmp_151 != io_wb_resps_9_bits_uop_pdst;
  reg        rob_unsafe_3_0;
  reg        rob_unsafe_3_1;
  reg        rob_unsafe_3_2;
  reg        rob_unsafe_3_3;
  reg        rob_unsafe_3_4;
  reg        rob_unsafe_3_5;
  reg        rob_unsafe_3_6;
  reg        rob_unsafe_3_7;
  reg        rob_unsafe_3_8;
  reg        rob_unsafe_3_9;
  reg        rob_unsafe_3_10;
  reg        rob_unsafe_3_11;
  reg        rob_unsafe_3_12;
  reg        rob_unsafe_3_13;
  reg        rob_unsafe_3_14;
  reg        rob_unsafe_3_15;
  reg        rob_unsafe_3_16;
  reg        rob_unsafe_3_17;
  reg        rob_unsafe_3_18;
  reg        rob_unsafe_3_19;
  reg        rob_unsafe_3_20;
  reg        rob_unsafe_3_21;
  reg        rob_unsafe_3_22;
  reg        rob_unsafe_3_23;
  reg        rob_unsafe_3_24;
  reg        rob_unsafe_3_25;
  reg        rob_unsafe_3_26;
  reg        rob_unsafe_3_27;
  reg        rob_unsafe_3_28;
  reg        rob_unsafe_3_29;
  reg        rob_unsafe_3_30;
  reg        rob_unsafe_3_31;
  always @(*) begin
    casez (rob_tail)
      5'b00000:
        casez_tmp_152 = rob_val_3_0;
      5'b00001:
        casez_tmp_152 = rob_val_3_1;
      5'b00010:
        casez_tmp_152 = rob_val_3_2;
      5'b00011:
        casez_tmp_152 = rob_val_3_3;
      5'b00100:
        casez_tmp_152 = rob_val_3_4;
      5'b00101:
        casez_tmp_152 = rob_val_3_5;
      5'b00110:
        casez_tmp_152 = rob_val_3_6;
      5'b00111:
        casez_tmp_152 = rob_val_3_7;
      5'b01000:
        casez_tmp_152 = rob_val_3_8;
      5'b01001:
        casez_tmp_152 = rob_val_3_9;
      5'b01010:
        casez_tmp_152 = rob_val_3_10;
      5'b01011:
        casez_tmp_152 = rob_val_3_11;
      5'b01100:
        casez_tmp_152 = rob_val_3_12;
      5'b01101:
        casez_tmp_152 = rob_val_3_13;
      5'b01110:
        casez_tmp_152 = rob_val_3_14;
      5'b01111:
        casez_tmp_152 = rob_val_3_15;
      5'b10000:
        casez_tmp_152 = rob_val_3_16;
      5'b10001:
        casez_tmp_152 = rob_val_3_17;
      5'b10010:
        casez_tmp_152 = rob_val_3_18;
      5'b10011:
        casez_tmp_152 = rob_val_3_19;
      5'b10100:
        casez_tmp_152 = rob_val_3_20;
      5'b10101:
        casez_tmp_152 = rob_val_3_21;
      5'b10110:
        casez_tmp_152 = rob_val_3_22;
      5'b10111:
        casez_tmp_152 = rob_val_3_23;
      5'b11000:
        casez_tmp_152 = rob_val_3_24;
      5'b11001:
        casez_tmp_152 = rob_val_3_25;
      5'b11010:
        casez_tmp_152 = rob_val_3_26;
      5'b11011:
        casez_tmp_152 = rob_val_3_27;
      5'b11100:
        casez_tmp_152 = rob_val_3_28;
      5'b11101:
        casez_tmp_152 = rob_val_3_29;
      5'b11110:
        casez_tmp_152 = rob_val_3_30;
      default:
        casez_tmp_152 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1947 = io_enq_uops_3_rob_idx[6:2] == rob_tail;
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_153 = rob_val_3_0;
      5'b00001:
        casez_tmp_153 = rob_val_3_1;
      5'b00010:
        casez_tmp_153 = rob_val_3_2;
      5'b00011:
        casez_tmp_153 = rob_val_3_3;
      5'b00100:
        casez_tmp_153 = rob_val_3_4;
      5'b00101:
        casez_tmp_153 = rob_val_3_5;
      5'b00110:
        casez_tmp_153 = rob_val_3_6;
      5'b00111:
        casez_tmp_153 = rob_val_3_7;
      5'b01000:
        casez_tmp_153 = rob_val_3_8;
      5'b01001:
        casez_tmp_153 = rob_val_3_9;
      5'b01010:
        casez_tmp_153 = rob_val_3_10;
      5'b01011:
        casez_tmp_153 = rob_val_3_11;
      5'b01100:
        casez_tmp_153 = rob_val_3_12;
      5'b01101:
        casez_tmp_153 = rob_val_3_13;
      5'b01110:
        casez_tmp_153 = rob_val_3_14;
      5'b01111:
        casez_tmp_153 = rob_val_3_15;
      5'b10000:
        casez_tmp_153 = rob_val_3_16;
      5'b10001:
        casez_tmp_153 = rob_val_3_17;
      5'b10010:
        casez_tmp_153 = rob_val_3_18;
      5'b10011:
        casez_tmp_153 = rob_val_3_19;
      5'b10100:
        casez_tmp_153 = rob_val_3_20;
      5'b10101:
        casez_tmp_153 = rob_val_3_21;
      5'b10110:
        casez_tmp_153 = rob_val_3_22;
      5'b10111:
        casez_tmp_153 = rob_val_3_23;
      5'b11000:
        casez_tmp_153 = rob_val_3_24;
      5'b11001:
        casez_tmp_153 = rob_val_3_25;
      5'b11010:
        casez_tmp_153 = rob_val_3_26;
      5'b11011:
        casez_tmp_153 = rob_val_3_27;
      5'b11100:
        casez_tmp_153 = rob_val_3_28;
      5'b11101:
        casez_tmp_153 = rob_val_3_29;
      5'b11110:
        casez_tmp_153 = rob_val_3_30;
      default:
        casez_tmp_153 = rob_val_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_154 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_154 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_154 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_154 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_154 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_154 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_154 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_154 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_154 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_154 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_154 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_154 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_154 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_154 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_154 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_154 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_154 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_154 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_154 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_154 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_154 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_154 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_154 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_154 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_154 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_154 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_154 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_154 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_154 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_154 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_154 = rob_bsy_3_30;
      default:
        casez_tmp_154 = rob_bsy_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_155 = rob_val_3_0;
      5'b00001:
        casez_tmp_155 = rob_val_3_1;
      5'b00010:
        casez_tmp_155 = rob_val_3_2;
      5'b00011:
        casez_tmp_155 = rob_val_3_3;
      5'b00100:
        casez_tmp_155 = rob_val_3_4;
      5'b00101:
        casez_tmp_155 = rob_val_3_5;
      5'b00110:
        casez_tmp_155 = rob_val_3_6;
      5'b00111:
        casez_tmp_155 = rob_val_3_7;
      5'b01000:
        casez_tmp_155 = rob_val_3_8;
      5'b01001:
        casez_tmp_155 = rob_val_3_9;
      5'b01010:
        casez_tmp_155 = rob_val_3_10;
      5'b01011:
        casez_tmp_155 = rob_val_3_11;
      5'b01100:
        casez_tmp_155 = rob_val_3_12;
      5'b01101:
        casez_tmp_155 = rob_val_3_13;
      5'b01110:
        casez_tmp_155 = rob_val_3_14;
      5'b01111:
        casez_tmp_155 = rob_val_3_15;
      5'b10000:
        casez_tmp_155 = rob_val_3_16;
      5'b10001:
        casez_tmp_155 = rob_val_3_17;
      5'b10010:
        casez_tmp_155 = rob_val_3_18;
      5'b10011:
        casez_tmp_155 = rob_val_3_19;
      5'b10100:
        casez_tmp_155 = rob_val_3_20;
      5'b10101:
        casez_tmp_155 = rob_val_3_21;
      5'b10110:
        casez_tmp_155 = rob_val_3_22;
      5'b10111:
        casez_tmp_155 = rob_val_3_23;
      5'b11000:
        casez_tmp_155 = rob_val_3_24;
      5'b11001:
        casez_tmp_155 = rob_val_3_25;
      5'b11010:
        casez_tmp_155 = rob_val_3_26;
      5'b11011:
        casez_tmp_155 = rob_val_3_27;
      5'b11100:
        casez_tmp_155 = rob_val_3_28;
      5'b11101:
        casez_tmp_155 = rob_val_3_29;
      5'b11110:
        casez_tmp_155 = rob_val_3_30;
      default:
        casez_tmp_155 = rob_val_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_156 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_156 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_156 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_156 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_156 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_156 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_156 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_156 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_156 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_156 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_156 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_156 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_156 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_156 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_156 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_156 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_156 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_156 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_156 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_156 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_156 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_156 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_156 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_156 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_156 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_156 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_156 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_156 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_156 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_156 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_156 = rob_bsy_3_30;
      default:
        casez_tmp_156 = rob_bsy_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_157 = rob_val_3_0;
      5'b00001:
        casez_tmp_157 = rob_val_3_1;
      5'b00010:
        casez_tmp_157 = rob_val_3_2;
      5'b00011:
        casez_tmp_157 = rob_val_3_3;
      5'b00100:
        casez_tmp_157 = rob_val_3_4;
      5'b00101:
        casez_tmp_157 = rob_val_3_5;
      5'b00110:
        casez_tmp_157 = rob_val_3_6;
      5'b00111:
        casez_tmp_157 = rob_val_3_7;
      5'b01000:
        casez_tmp_157 = rob_val_3_8;
      5'b01001:
        casez_tmp_157 = rob_val_3_9;
      5'b01010:
        casez_tmp_157 = rob_val_3_10;
      5'b01011:
        casez_tmp_157 = rob_val_3_11;
      5'b01100:
        casez_tmp_157 = rob_val_3_12;
      5'b01101:
        casez_tmp_157 = rob_val_3_13;
      5'b01110:
        casez_tmp_157 = rob_val_3_14;
      5'b01111:
        casez_tmp_157 = rob_val_3_15;
      5'b10000:
        casez_tmp_157 = rob_val_3_16;
      5'b10001:
        casez_tmp_157 = rob_val_3_17;
      5'b10010:
        casez_tmp_157 = rob_val_3_18;
      5'b10011:
        casez_tmp_157 = rob_val_3_19;
      5'b10100:
        casez_tmp_157 = rob_val_3_20;
      5'b10101:
        casez_tmp_157 = rob_val_3_21;
      5'b10110:
        casez_tmp_157 = rob_val_3_22;
      5'b10111:
        casez_tmp_157 = rob_val_3_23;
      5'b11000:
        casez_tmp_157 = rob_val_3_24;
      5'b11001:
        casez_tmp_157 = rob_val_3_25;
      5'b11010:
        casez_tmp_157 = rob_val_3_26;
      5'b11011:
        casez_tmp_157 = rob_val_3_27;
      5'b11100:
        casez_tmp_157 = rob_val_3_28;
      5'b11101:
        casez_tmp_157 = rob_val_3_29;
      5'b11110:
        casez_tmp_157 = rob_val_3_30;
      default:
        casez_tmp_157 = rob_val_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_158 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_158 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_158 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_158 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_158 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_158 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_158 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_158 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_158 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_158 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_158 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_158 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_158 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_158 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_158 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_158 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_158 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_158 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_158 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_158 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_158 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_158 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_158 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_158 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_158 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_158 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_158 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_158 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_158 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_158 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_158 = rob_bsy_3_30;
      default:
        casez_tmp_158 = rob_bsy_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_GEN_2)
      5'b00000:
        casez_tmp_159 = rob_unsafe_3_0;
      5'b00001:
        casez_tmp_159 = rob_unsafe_3_1;
      5'b00010:
        casez_tmp_159 = rob_unsafe_3_2;
      5'b00011:
        casez_tmp_159 = rob_unsafe_3_3;
      5'b00100:
        casez_tmp_159 = rob_unsafe_3_4;
      5'b00101:
        casez_tmp_159 = rob_unsafe_3_5;
      5'b00110:
        casez_tmp_159 = rob_unsafe_3_6;
      5'b00111:
        casez_tmp_159 = rob_unsafe_3_7;
      5'b01000:
        casez_tmp_159 = rob_unsafe_3_8;
      5'b01001:
        casez_tmp_159 = rob_unsafe_3_9;
      5'b01010:
        casez_tmp_159 = rob_unsafe_3_10;
      5'b01011:
        casez_tmp_159 = rob_unsafe_3_11;
      5'b01100:
        casez_tmp_159 = rob_unsafe_3_12;
      5'b01101:
        casez_tmp_159 = rob_unsafe_3_13;
      5'b01110:
        casez_tmp_159 = rob_unsafe_3_14;
      5'b01111:
        casez_tmp_159 = rob_unsafe_3_15;
      5'b10000:
        casez_tmp_159 = rob_unsafe_3_16;
      5'b10001:
        casez_tmp_159 = rob_unsafe_3_17;
      5'b10010:
        casez_tmp_159 = rob_unsafe_3_18;
      5'b10011:
        casez_tmp_159 = rob_unsafe_3_19;
      5'b10100:
        casez_tmp_159 = rob_unsafe_3_20;
      5'b10101:
        casez_tmp_159 = rob_unsafe_3_21;
      5'b10110:
        casez_tmp_159 = rob_unsafe_3_22;
      5'b10111:
        casez_tmp_159 = rob_unsafe_3_23;
      5'b11000:
        casez_tmp_159 = rob_unsafe_3_24;
      5'b11001:
        casez_tmp_159 = rob_unsafe_3_25;
      5'b11010:
        casez_tmp_159 = rob_unsafe_3_26;
      5'b11011:
        casez_tmp_159 = rob_unsafe_3_27;
      5'b11100:
        casez_tmp_159 = rob_unsafe_3_28;
      5'b11101:
        casez_tmp_159 = rob_unsafe_3_29;
      5'b11110:
        casez_tmp_159 = rob_unsafe_3_30;
      default:
        casez_tmp_159 = rob_unsafe_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_160 = rob_unsafe_3_0;
      5'b00001:
        casez_tmp_160 = rob_unsafe_3_1;
      5'b00010:
        casez_tmp_160 = rob_unsafe_3_2;
      5'b00011:
        casez_tmp_160 = rob_unsafe_3_3;
      5'b00100:
        casez_tmp_160 = rob_unsafe_3_4;
      5'b00101:
        casez_tmp_160 = rob_unsafe_3_5;
      5'b00110:
        casez_tmp_160 = rob_unsafe_3_6;
      5'b00111:
        casez_tmp_160 = rob_unsafe_3_7;
      5'b01000:
        casez_tmp_160 = rob_unsafe_3_8;
      5'b01001:
        casez_tmp_160 = rob_unsafe_3_9;
      5'b01010:
        casez_tmp_160 = rob_unsafe_3_10;
      5'b01011:
        casez_tmp_160 = rob_unsafe_3_11;
      5'b01100:
        casez_tmp_160 = rob_unsafe_3_12;
      5'b01101:
        casez_tmp_160 = rob_unsafe_3_13;
      5'b01110:
        casez_tmp_160 = rob_unsafe_3_14;
      5'b01111:
        casez_tmp_160 = rob_unsafe_3_15;
      5'b10000:
        casez_tmp_160 = rob_unsafe_3_16;
      5'b10001:
        casez_tmp_160 = rob_unsafe_3_17;
      5'b10010:
        casez_tmp_160 = rob_unsafe_3_18;
      5'b10011:
        casez_tmp_160 = rob_unsafe_3_19;
      5'b10100:
        casez_tmp_160 = rob_unsafe_3_20;
      5'b10101:
        casez_tmp_160 = rob_unsafe_3_21;
      5'b10110:
        casez_tmp_160 = rob_unsafe_3_22;
      5'b10111:
        casez_tmp_160 = rob_unsafe_3_23;
      5'b11000:
        casez_tmp_160 = rob_unsafe_3_24;
      5'b11001:
        casez_tmp_160 = rob_unsafe_3_25;
      5'b11010:
        casez_tmp_160 = rob_unsafe_3_26;
      5'b11011:
        casez_tmp_160 = rob_unsafe_3_27;
      5'b11100:
        casez_tmp_160 = rob_unsafe_3_28;
      5'b11101:
        casez_tmp_160 = rob_unsafe_3_29;
      5'b11110:
        casez_tmp_160 = rob_unsafe_3_30;
      default:
        casez_tmp_160 = rob_unsafe_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_161 = rob_exception_3_0;
      5'b00001:
        casez_tmp_161 = rob_exception_3_1;
      5'b00010:
        casez_tmp_161 = rob_exception_3_2;
      5'b00011:
        casez_tmp_161 = rob_exception_3_3;
      5'b00100:
        casez_tmp_161 = rob_exception_3_4;
      5'b00101:
        casez_tmp_161 = rob_exception_3_5;
      5'b00110:
        casez_tmp_161 = rob_exception_3_6;
      5'b00111:
        casez_tmp_161 = rob_exception_3_7;
      5'b01000:
        casez_tmp_161 = rob_exception_3_8;
      5'b01001:
        casez_tmp_161 = rob_exception_3_9;
      5'b01010:
        casez_tmp_161 = rob_exception_3_10;
      5'b01011:
        casez_tmp_161 = rob_exception_3_11;
      5'b01100:
        casez_tmp_161 = rob_exception_3_12;
      5'b01101:
        casez_tmp_161 = rob_exception_3_13;
      5'b01110:
        casez_tmp_161 = rob_exception_3_14;
      5'b01111:
        casez_tmp_161 = rob_exception_3_15;
      5'b10000:
        casez_tmp_161 = rob_exception_3_16;
      5'b10001:
        casez_tmp_161 = rob_exception_3_17;
      5'b10010:
        casez_tmp_161 = rob_exception_3_18;
      5'b10011:
        casez_tmp_161 = rob_exception_3_19;
      5'b10100:
        casez_tmp_161 = rob_exception_3_20;
      5'b10101:
        casez_tmp_161 = rob_exception_3_21;
      5'b10110:
        casez_tmp_161 = rob_exception_3_22;
      5'b10111:
        casez_tmp_161 = rob_exception_3_23;
      5'b11000:
        casez_tmp_161 = rob_exception_3_24;
      5'b11001:
        casez_tmp_161 = rob_exception_3_25;
      5'b11010:
        casez_tmp_161 = rob_exception_3_26;
      5'b11011:
        casez_tmp_161 = rob_exception_3_27;
      5'b11100:
        casez_tmp_161 = rob_exception_3_28;
      5'b11101:
        casez_tmp_161 = rob_exception_3_29;
      5'b11110:
        casez_tmp_161 = rob_exception_3_30;
      default:
        casez_tmp_161 = rob_exception_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_pnr)
      5'b00000:
        casez_tmp_162 = rob_val_3_0;
      5'b00001:
        casez_tmp_162 = rob_val_3_1;
      5'b00010:
        casez_tmp_162 = rob_val_3_2;
      5'b00011:
        casez_tmp_162 = rob_val_3_3;
      5'b00100:
        casez_tmp_162 = rob_val_3_4;
      5'b00101:
        casez_tmp_162 = rob_val_3_5;
      5'b00110:
        casez_tmp_162 = rob_val_3_6;
      5'b00111:
        casez_tmp_162 = rob_val_3_7;
      5'b01000:
        casez_tmp_162 = rob_val_3_8;
      5'b01001:
        casez_tmp_162 = rob_val_3_9;
      5'b01010:
        casez_tmp_162 = rob_val_3_10;
      5'b01011:
        casez_tmp_162 = rob_val_3_11;
      5'b01100:
        casez_tmp_162 = rob_val_3_12;
      5'b01101:
        casez_tmp_162 = rob_val_3_13;
      5'b01110:
        casez_tmp_162 = rob_val_3_14;
      5'b01111:
        casez_tmp_162 = rob_val_3_15;
      5'b10000:
        casez_tmp_162 = rob_val_3_16;
      5'b10001:
        casez_tmp_162 = rob_val_3_17;
      5'b10010:
        casez_tmp_162 = rob_val_3_18;
      5'b10011:
        casez_tmp_162 = rob_val_3_19;
      5'b10100:
        casez_tmp_162 = rob_val_3_20;
      5'b10101:
        casez_tmp_162 = rob_val_3_21;
      5'b10110:
        casez_tmp_162 = rob_val_3_22;
      5'b10111:
        casez_tmp_162 = rob_val_3_23;
      5'b11000:
        casez_tmp_162 = rob_val_3_24;
      5'b11001:
        casez_tmp_162 = rob_val_3_25;
      5'b11010:
        casez_tmp_162 = rob_val_3_26;
      5'b11011:
        casez_tmp_162 = rob_val_3_27;
      5'b11100:
        casez_tmp_162 = rob_val_3_28;
      5'b11101:
        casez_tmp_162 = rob_val_3_29;
      5'b11110:
        casez_tmp_162 = rob_val_3_30;
      default:
        casez_tmp_162 = rob_val_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_163 = rob_val_3_0;
      5'b00001:
        casez_tmp_163 = rob_val_3_1;
      5'b00010:
        casez_tmp_163 = rob_val_3_2;
      5'b00011:
        casez_tmp_163 = rob_val_3_3;
      5'b00100:
        casez_tmp_163 = rob_val_3_4;
      5'b00101:
        casez_tmp_163 = rob_val_3_5;
      5'b00110:
        casez_tmp_163 = rob_val_3_6;
      5'b00111:
        casez_tmp_163 = rob_val_3_7;
      5'b01000:
        casez_tmp_163 = rob_val_3_8;
      5'b01001:
        casez_tmp_163 = rob_val_3_9;
      5'b01010:
        casez_tmp_163 = rob_val_3_10;
      5'b01011:
        casez_tmp_163 = rob_val_3_11;
      5'b01100:
        casez_tmp_163 = rob_val_3_12;
      5'b01101:
        casez_tmp_163 = rob_val_3_13;
      5'b01110:
        casez_tmp_163 = rob_val_3_14;
      5'b01111:
        casez_tmp_163 = rob_val_3_15;
      5'b10000:
        casez_tmp_163 = rob_val_3_16;
      5'b10001:
        casez_tmp_163 = rob_val_3_17;
      5'b10010:
        casez_tmp_163 = rob_val_3_18;
      5'b10011:
        casez_tmp_163 = rob_val_3_19;
      5'b10100:
        casez_tmp_163 = rob_val_3_20;
      5'b10101:
        casez_tmp_163 = rob_val_3_21;
      5'b10110:
        casez_tmp_163 = rob_val_3_22;
      5'b10111:
        casez_tmp_163 = rob_val_3_23;
      5'b11000:
        casez_tmp_163 = rob_val_3_24;
      5'b11001:
        casez_tmp_163 = rob_val_3_25;
      5'b11010:
        casez_tmp_163 = rob_val_3_26;
      5'b11011:
        casez_tmp_163 = rob_val_3_27;
      5'b11100:
        casez_tmp_163 = rob_val_3_28;
      5'b11101:
        casez_tmp_163 = rob_val_3_29;
      5'b11110:
        casez_tmp_163 = rob_val_3_30;
      default:
        casez_tmp_163 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1948 = _GEN_1834 & ~casez_tmp_163;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_164 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_164 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_164 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_164 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_164 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_164 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_164 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_164 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_164 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_164 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_164 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_164 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_164 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_164 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_164 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_164 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_164 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_164 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_164 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_164 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_164 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_164 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_164 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_164 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_164 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_164 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_164 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_164 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_164 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_164 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_164 = rob_bsy_3_30;
      default:
        casez_tmp_164 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1949 = _GEN_1834 & ~casez_tmp_164;
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_165 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_165 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_165 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_165 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_165 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_165 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_165 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_165 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_165 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_165 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_165 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_165 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_165 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_165 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_165 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_165 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_165 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_165 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_165 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_165 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_165 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_165 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_165 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_165 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_165 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_165 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_165 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_165 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_165 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_165 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_165 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_165 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_61)
      5'b00000:
        casez_tmp_166 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_166 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_166 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_166 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_166 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_166 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_166 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_166 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_166 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_166 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_166 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_166 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_166 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_166 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_166 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_166 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_166 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_166 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_166 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_166 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_166 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_166 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_166 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_166 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_166 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_166 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_166 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_166 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_166 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_166 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_166 = rob_uop_3_30_pdst;
      default:
        casez_tmp_166 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1950 = _GEN_1834 & casez_tmp_165 & casez_tmp_166 != io_wb_resps_0_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_167 = rob_val_3_0;
      5'b00001:
        casez_tmp_167 = rob_val_3_1;
      5'b00010:
        casez_tmp_167 = rob_val_3_2;
      5'b00011:
        casez_tmp_167 = rob_val_3_3;
      5'b00100:
        casez_tmp_167 = rob_val_3_4;
      5'b00101:
        casez_tmp_167 = rob_val_3_5;
      5'b00110:
        casez_tmp_167 = rob_val_3_6;
      5'b00111:
        casez_tmp_167 = rob_val_3_7;
      5'b01000:
        casez_tmp_167 = rob_val_3_8;
      5'b01001:
        casez_tmp_167 = rob_val_3_9;
      5'b01010:
        casez_tmp_167 = rob_val_3_10;
      5'b01011:
        casez_tmp_167 = rob_val_3_11;
      5'b01100:
        casez_tmp_167 = rob_val_3_12;
      5'b01101:
        casez_tmp_167 = rob_val_3_13;
      5'b01110:
        casez_tmp_167 = rob_val_3_14;
      5'b01111:
        casez_tmp_167 = rob_val_3_15;
      5'b10000:
        casez_tmp_167 = rob_val_3_16;
      5'b10001:
        casez_tmp_167 = rob_val_3_17;
      5'b10010:
        casez_tmp_167 = rob_val_3_18;
      5'b10011:
        casez_tmp_167 = rob_val_3_19;
      5'b10100:
        casez_tmp_167 = rob_val_3_20;
      5'b10101:
        casez_tmp_167 = rob_val_3_21;
      5'b10110:
        casez_tmp_167 = rob_val_3_22;
      5'b10111:
        casez_tmp_167 = rob_val_3_23;
      5'b11000:
        casez_tmp_167 = rob_val_3_24;
      5'b11001:
        casez_tmp_167 = rob_val_3_25;
      5'b11010:
        casez_tmp_167 = rob_val_3_26;
      5'b11011:
        casez_tmp_167 = rob_val_3_27;
      5'b11100:
        casez_tmp_167 = rob_val_3_28;
      5'b11101:
        casez_tmp_167 = rob_val_3_29;
      5'b11110:
        casez_tmp_167 = rob_val_3_30;
      default:
        casez_tmp_167 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1951 = _GEN_1385 & ~casez_tmp_167;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_168 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_168 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_168 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_168 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_168 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_168 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_168 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_168 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_168 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_168 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_168 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_168 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_168 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_168 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_168 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_168 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_168 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_168 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_168 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_168 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_168 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_168 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_168 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_168 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_168 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_168 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_168 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_168 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_168 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_168 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_168 = rob_bsy_3_30;
      default:
        casez_tmp_168 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1952 = _GEN_1385 & ~casez_tmp_168;
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_169 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_169 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_169 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_169 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_169 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_169 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_169 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_169 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_169 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_169 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_169 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_169 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_169 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_169 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_169 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_169 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_169 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_169 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_169 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_169 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_169 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_169 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_169 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_169 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_169 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_169 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_169 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_169 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_169 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_169 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_169 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_169 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_63)
      5'b00000:
        casez_tmp_170 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_170 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_170 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_170 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_170 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_170 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_170 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_170 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_170 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_170 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_170 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_170 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_170 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_170 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_170 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_170 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_170 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_170 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_170 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_170 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_170 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_170 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_170 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_170 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_170 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_170 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_170 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_170 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_170 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_170 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_170 = rob_uop_3_30_pdst;
      default:
        casez_tmp_170 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1953 = _GEN_1385 & casez_tmp_169 & casez_tmp_170 != io_wb_resps_1_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_171 = rob_val_3_0;
      5'b00001:
        casez_tmp_171 = rob_val_3_1;
      5'b00010:
        casez_tmp_171 = rob_val_3_2;
      5'b00011:
        casez_tmp_171 = rob_val_3_3;
      5'b00100:
        casez_tmp_171 = rob_val_3_4;
      5'b00101:
        casez_tmp_171 = rob_val_3_5;
      5'b00110:
        casez_tmp_171 = rob_val_3_6;
      5'b00111:
        casez_tmp_171 = rob_val_3_7;
      5'b01000:
        casez_tmp_171 = rob_val_3_8;
      5'b01001:
        casez_tmp_171 = rob_val_3_9;
      5'b01010:
        casez_tmp_171 = rob_val_3_10;
      5'b01011:
        casez_tmp_171 = rob_val_3_11;
      5'b01100:
        casez_tmp_171 = rob_val_3_12;
      5'b01101:
        casez_tmp_171 = rob_val_3_13;
      5'b01110:
        casez_tmp_171 = rob_val_3_14;
      5'b01111:
        casez_tmp_171 = rob_val_3_15;
      5'b10000:
        casez_tmp_171 = rob_val_3_16;
      5'b10001:
        casez_tmp_171 = rob_val_3_17;
      5'b10010:
        casez_tmp_171 = rob_val_3_18;
      5'b10011:
        casez_tmp_171 = rob_val_3_19;
      5'b10100:
        casez_tmp_171 = rob_val_3_20;
      5'b10101:
        casez_tmp_171 = rob_val_3_21;
      5'b10110:
        casez_tmp_171 = rob_val_3_22;
      5'b10111:
        casez_tmp_171 = rob_val_3_23;
      5'b11000:
        casez_tmp_171 = rob_val_3_24;
      5'b11001:
        casez_tmp_171 = rob_val_3_25;
      5'b11010:
        casez_tmp_171 = rob_val_3_26;
      5'b11011:
        casez_tmp_171 = rob_val_3_27;
      5'b11100:
        casez_tmp_171 = rob_val_3_28;
      5'b11101:
        casez_tmp_171 = rob_val_3_29;
      5'b11110:
        casez_tmp_171 = rob_val_3_30;
      default:
        casez_tmp_171 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1954 = _GEN_1835 & ~casez_tmp_171;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_172 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_172 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_172 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_172 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_172 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_172 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_172 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_172 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_172 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_172 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_172 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_172 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_172 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_172 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_172 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_172 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_172 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_172 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_172 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_172 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_172 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_172 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_172 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_172 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_172 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_172 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_172 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_172 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_172 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_172 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_172 = rob_bsy_3_30;
      default:
        casez_tmp_172 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1955 = _GEN_1835 & ~casez_tmp_172;
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_173 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_173 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_173 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_173 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_173 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_173 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_173 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_173 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_173 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_173 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_173 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_173 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_173 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_173 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_173 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_173 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_173 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_173 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_173 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_173 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_173 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_173 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_173 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_173 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_173 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_173 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_173 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_173 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_173 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_173 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_173 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_173 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_65)
      5'b00000:
        casez_tmp_174 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_174 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_174 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_174 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_174 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_174 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_174 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_174 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_174 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_174 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_174 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_174 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_174 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_174 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_174 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_174 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_174 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_174 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_174 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_174 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_174 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_174 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_174 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_174 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_174 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_174 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_174 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_174 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_174 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_174 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_174 = rob_uop_3_30_pdst;
      default:
        casez_tmp_174 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1956 = _GEN_1835 & casez_tmp_173 & casez_tmp_174 != io_wb_resps_2_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_175 = rob_val_3_0;
      5'b00001:
        casez_tmp_175 = rob_val_3_1;
      5'b00010:
        casez_tmp_175 = rob_val_3_2;
      5'b00011:
        casez_tmp_175 = rob_val_3_3;
      5'b00100:
        casez_tmp_175 = rob_val_3_4;
      5'b00101:
        casez_tmp_175 = rob_val_3_5;
      5'b00110:
        casez_tmp_175 = rob_val_3_6;
      5'b00111:
        casez_tmp_175 = rob_val_3_7;
      5'b01000:
        casez_tmp_175 = rob_val_3_8;
      5'b01001:
        casez_tmp_175 = rob_val_3_9;
      5'b01010:
        casez_tmp_175 = rob_val_3_10;
      5'b01011:
        casez_tmp_175 = rob_val_3_11;
      5'b01100:
        casez_tmp_175 = rob_val_3_12;
      5'b01101:
        casez_tmp_175 = rob_val_3_13;
      5'b01110:
        casez_tmp_175 = rob_val_3_14;
      5'b01111:
        casez_tmp_175 = rob_val_3_15;
      5'b10000:
        casez_tmp_175 = rob_val_3_16;
      5'b10001:
        casez_tmp_175 = rob_val_3_17;
      5'b10010:
        casez_tmp_175 = rob_val_3_18;
      5'b10011:
        casez_tmp_175 = rob_val_3_19;
      5'b10100:
        casez_tmp_175 = rob_val_3_20;
      5'b10101:
        casez_tmp_175 = rob_val_3_21;
      5'b10110:
        casez_tmp_175 = rob_val_3_22;
      5'b10111:
        casez_tmp_175 = rob_val_3_23;
      5'b11000:
        casez_tmp_175 = rob_val_3_24;
      5'b11001:
        casez_tmp_175 = rob_val_3_25;
      5'b11010:
        casez_tmp_175 = rob_val_3_26;
      5'b11011:
        casez_tmp_175 = rob_val_3_27;
      5'b11100:
        casez_tmp_175 = rob_val_3_28;
      5'b11101:
        casez_tmp_175 = rob_val_3_29;
      5'b11110:
        casez_tmp_175 = rob_val_3_30;
      default:
        casez_tmp_175 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1957 = _GEN_1384 & ~casez_tmp_175;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_176 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_176 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_176 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_176 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_176 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_176 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_176 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_176 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_176 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_176 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_176 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_176 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_176 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_176 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_176 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_176 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_176 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_176 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_176 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_176 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_176 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_176 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_176 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_176 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_176 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_176 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_176 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_176 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_176 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_176 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_176 = rob_bsy_3_30;
      default:
        casez_tmp_176 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1958 = _GEN_1384 & ~casez_tmp_176;
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_177 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_177 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_177 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_177 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_177 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_177 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_177 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_177 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_177 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_177 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_177 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_177 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_177 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_177 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_177 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_177 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_177 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_177 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_177 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_177 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_177 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_177 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_177 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_177 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_177 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_177 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_177 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_177 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_177 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_177 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_177 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_177 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_67)
      5'b00000:
        casez_tmp_178 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_178 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_178 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_178 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_178 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_178 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_178 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_178 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_178 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_178 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_178 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_178 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_178 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_178 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_178 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_178 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_178 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_178 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_178 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_178 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_178 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_178 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_178 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_178 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_178 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_178 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_178 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_178 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_178 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_178 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_178 = rob_uop_3_30_pdst;
      default:
        casez_tmp_178 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1959 = _GEN_1384 & casez_tmp_177 & casez_tmp_178 != io_wb_resps_3_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_179 = rob_val_3_0;
      5'b00001:
        casez_tmp_179 = rob_val_3_1;
      5'b00010:
        casez_tmp_179 = rob_val_3_2;
      5'b00011:
        casez_tmp_179 = rob_val_3_3;
      5'b00100:
        casez_tmp_179 = rob_val_3_4;
      5'b00101:
        casez_tmp_179 = rob_val_3_5;
      5'b00110:
        casez_tmp_179 = rob_val_3_6;
      5'b00111:
        casez_tmp_179 = rob_val_3_7;
      5'b01000:
        casez_tmp_179 = rob_val_3_8;
      5'b01001:
        casez_tmp_179 = rob_val_3_9;
      5'b01010:
        casez_tmp_179 = rob_val_3_10;
      5'b01011:
        casez_tmp_179 = rob_val_3_11;
      5'b01100:
        casez_tmp_179 = rob_val_3_12;
      5'b01101:
        casez_tmp_179 = rob_val_3_13;
      5'b01110:
        casez_tmp_179 = rob_val_3_14;
      5'b01111:
        casez_tmp_179 = rob_val_3_15;
      5'b10000:
        casez_tmp_179 = rob_val_3_16;
      5'b10001:
        casez_tmp_179 = rob_val_3_17;
      5'b10010:
        casez_tmp_179 = rob_val_3_18;
      5'b10011:
        casez_tmp_179 = rob_val_3_19;
      5'b10100:
        casez_tmp_179 = rob_val_3_20;
      5'b10101:
        casez_tmp_179 = rob_val_3_21;
      5'b10110:
        casez_tmp_179 = rob_val_3_22;
      5'b10111:
        casez_tmp_179 = rob_val_3_23;
      5'b11000:
        casez_tmp_179 = rob_val_3_24;
      5'b11001:
        casez_tmp_179 = rob_val_3_25;
      5'b11010:
        casez_tmp_179 = rob_val_3_26;
      5'b11011:
        casez_tmp_179 = rob_val_3_27;
      5'b11100:
        casez_tmp_179 = rob_val_3_28;
      5'b11101:
        casez_tmp_179 = rob_val_3_29;
      5'b11110:
        casez_tmp_179 = rob_val_3_30;
      default:
        casez_tmp_179 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1960 = _GEN_1836 & ~casez_tmp_179;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_180 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_180 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_180 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_180 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_180 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_180 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_180 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_180 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_180 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_180 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_180 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_180 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_180 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_180 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_180 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_180 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_180 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_180 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_180 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_180 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_180 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_180 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_180 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_180 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_180 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_180 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_180 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_180 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_180 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_180 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_180 = rob_bsy_3_30;
      default:
        casez_tmp_180 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1961 = _GEN_1836 & ~casez_tmp_180;
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_181 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_181 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_181 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_181 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_181 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_181 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_181 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_181 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_181 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_181 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_181 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_181 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_181 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_181 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_181 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_181 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_181 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_181 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_181 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_181 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_181 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_181 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_181 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_181 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_181 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_181 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_181 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_181 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_181 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_181 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_181 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_181 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_69)
      5'b00000:
        casez_tmp_182 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_182 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_182 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_182 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_182 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_182 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_182 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_182 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_182 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_182 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_182 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_182 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_182 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_182 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_182 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_182 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_182 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_182 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_182 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_182 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_182 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_182 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_182 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_182 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_182 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_182 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_182 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_182 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_182 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_182 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_182 = rob_uop_3_30_pdst;
      default:
        casez_tmp_182 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1962 = _GEN_1836 & casez_tmp_181 & casez_tmp_182 != io_wb_resps_4_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_183 = rob_val_3_0;
      5'b00001:
        casez_tmp_183 = rob_val_3_1;
      5'b00010:
        casez_tmp_183 = rob_val_3_2;
      5'b00011:
        casez_tmp_183 = rob_val_3_3;
      5'b00100:
        casez_tmp_183 = rob_val_3_4;
      5'b00101:
        casez_tmp_183 = rob_val_3_5;
      5'b00110:
        casez_tmp_183 = rob_val_3_6;
      5'b00111:
        casez_tmp_183 = rob_val_3_7;
      5'b01000:
        casez_tmp_183 = rob_val_3_8;
      5'b01001:
        casez_tmp_183 = rob_val_3_9;
      5'b01010:
        casez_tmp_183 = rob_val_3_10;
      5'b01011:
        casez_tmp_183 = rob_val_3_11;
      5'b01100:
        casez_tmp_183 = rob_val_3_12;
      5'b01101:
        casez_tmp_183 = rob_val_3_13;
      5'b01110:
        casez_tmp_183 = rob_val_3_14;
      5'b01111:
        casez_tmp_183 = rob_val_3_15;
      5'b10000:
        casez_tmp_183 = rob_val_3_16;
      5'b10001:
        casez_tmp_183 = rob_val_3_17;
      5'b10010:
        casez_tmp_183 = rob_val_3_18;
      5'b10011:
        casez_tmp_183 = rob_val_3_19;
      5'b10100:
        casez_tmp_183 = rob_val_3_20;
      5'b10101:
        casez_tmp_183 = rob_val_3_21;
      5'b10110:
        casez_tmp_183 = rob_val_3_22;
      5'b10111:
        casez_tmp_183 = rob_val_3_23;
      5'b11000:
        casez_tmp_183 = rob_val_3_24;
      5'b11001:
        casez_tmp_183 = rob_val_3_25;
      5'b11010:
        casez_tmp_183 = rob_val_3_26;
      5'b11011:
        casez_tmp_183 = rob_val_3_27;
      5'b11100:
        casez_tmp_183 = rob_val_3_28;
      5'b11101:
        casez_tmp_183 = rob_val_3_29;
      5'b11110:
        casez_tmp_183 = rob_val_3_30;
      default:
        casez_tmp_183 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1963 = _GEN_1383 & ~casez_tmp_183;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_184 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_184 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_184 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_184 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_184 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_184 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_184 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_184 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_184 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_184 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_184 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_184 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_184 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_184 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_184 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_184 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_184 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_184 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_184 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_184 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_184 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_184 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_184 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_184 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_184 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_184 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_184 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_184 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_184 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_184 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_184 = rob_bsy_3_30;
      default:
        casez_tmp_184 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1964 = _GEN_1383 & ~casez_tmp_184;
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_185 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_185 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_185 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_185 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_185 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_185 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_185 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_185 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_185 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_185 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_185 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_185 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_185 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_185 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_185 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_185 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_185 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_185 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_185 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_185 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_185 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_185 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_185 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_185 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_185 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_185 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_185 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_185 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_185 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_185 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_185 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_185 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_71)
      5'b00000:
        casez_tmp_186 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_186 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_186 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_186 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_186 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_186 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_186 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_186 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_186 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_186 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_186 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_186 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_186 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_186 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_186 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_186 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_186 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_186 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_186 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_186 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_186 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_186 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_186 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_186 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_186 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_186 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_186 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_186 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_186 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_186 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_186 = rob_uop_3_30_pdst;
      default:
        casez_tmp_186 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1965 = _GEN_1383 & casez_tmp_185 & casez_tmp_186 != io_wb_resps_5_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_187 = rob_val_3_0;
      5'b00001:
        casez_tmp_187 = rob_val_3_1;
      5'b00010:
        casez_tmp_187 = rob_val_3_2;
      5'b00011:
        casez_tmp_187 = rob_val_3_3;
      5'b00100:
        casez_tmp_187 = rob_val_3_4;
      5'b00101:
        casez_tmp_187 = rob_val_3_5;
      5'b00110:
        casez_tmp_187 = rob_val_3_6;
      5'b00111:
        casez_tmp_187 = rob_val_3_7;
      5'b01000:
        casez_tmp_187 = rob_val_3_8;
      5'b01001:
        casez_tmp_187 = rob_val_3_9;
      5'b01010:
        casez_tmp_187 = rob_val_3_10;
      5'b01011:
        casez_tmp_187 = rob_val_3_11;
      5'b01100:
        casez_tmp_187 = rob_val_3_12;
      5'b01101:
        casez_tmp_187 = rob_val_3_13;
      5'b01110:
        casez_tmp_187 = rob_val_3_14;
      5'b01111:
        casez_tmp_187 = rob_val_3_15;
      5'b10000:
        casez_tmp_187 = rob_val_3_16;
      5'b10001:
        casez_tmp_187 = rob_val_3_17;
      5'b10010:
        casez_tmp_187 = rob_val_3_18;
      5'b10011:
        casez_tmp_187 = rob_val_3_19;
      5'b10100:
        casez_tmp_187 = rob_val_3_20;
      5'b10101:
        casez_tmp_187 = rob_val_3_21;
      5'b10110:
        casez_tmp_187 = rob_val_3_22;
      5'b10111:
        casez_tmp_187 = rob_val_3_23;
      5'b11000:
        casez_tmp_187 = rob_val_3_24;
      5'b11001:
        casez_tmp_187 = rob_val_3_25;
      5'b11010:
        casez_tmp_187 = rob_val_3_26;
      5'b11011:
        casez_tmp_187 = rob_val_3_27;
      5'b11100:
        casez_tmp_187 = rob_val_3_28;
      5'b11101:
        casez_tmp_187 = rob_val_3_29;
      5'b11110:
        casez_tmp_187 = rob_val_3_30;
      default:
        casez_tmp_187 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1966 = _GEN_1837 & ~casez_tmp_187;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_188 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_188 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_188 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_188 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_188 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_188 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_188 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_188 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_188 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_188 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_188 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_188 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_188 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_188 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_188 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_188 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_188 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_188 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_188 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_188 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_188 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_188 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_188 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_188 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_188 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_188 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_188 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_188 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_188 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_188 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_188 = rob_bsy_3_30;
      default:
        casez_tmp_188 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1967 = _GEN_1837 & ~casez_tmp_188;
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_189 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_189 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_189 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_189 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_189 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_189 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_189 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_189 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_189 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_189 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_189 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_189 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_189 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_189 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_189 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_189 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_189 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_189 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_189 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_189 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_189 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_189 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_189 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_189 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_189 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_189 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_189 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_189 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_189 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_189 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_189 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_189 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_73)
      5'b00000:
        casez_tmp_190 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_190 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_190 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_190 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_190 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_190 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_190 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_190 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_190 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_190 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_190 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_190 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_190 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_190 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_190 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_190 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_190 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_190 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_190 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_190 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_190 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_190 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_190 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_190 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_190 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_190 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_190 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_190 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_190 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_190 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_190 = rob_uop_3_30_pdst;
      default:
        casez_tmp_190 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1968 = _GEN_1837 & casez_tmp_189 & casez_tmp_190 != io_wb_resps_6_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_191 = rob_val_3_0;
      5'b00001:
        casez_tmp_191 = rob_val_3_1;
      5'b00010:
        casez_tmp_191 = rob_val_3_2;
      5'b00011:
        casez_tmp_191 = rob_val_3_3;
      5'b00100:
        casez_tmp_191 = rob_val_3_4;
      5'b00101:
        casez_tmp_191 = rob_val_3_5;
      5'b00110:
        casez_tmp_191 = rob_val_3_6;
      5'b00111:
        casez_tmp_191 = rob_val_3_7;
      5'b01000:
        casez_tmp_191 = rob_val_3_8;
      5'b01001:
        casez_tmp_191 = rob_val_3_9;
      5'b01010:
        casez_tmp_191 = rob_val_3_10;
      5'b01011:
        casez_tmp_191 = rob_val_3_11;
      5'b01100:
        casez_tmp_191 = rob_val_3_12;
      5'b01101:
        casez_tmp_191 = rob_val_3_13;
      5'b01110:
        casez_tmp_191 = rob_val_3_14;
      5'b01111:
        casez_tmp_191 = rob_val_3_15;
      5'b10000:
        casez_tmp_191 = rob_val_3_16;
      5'b10001:
        casez_tmp_191 = rob_val_3_17;
      5'b10010:
        casez_tmp_191 = rob_val_3_18;
      5'b10011:
        casez_tmp_191 = rob_val_3_19;
      5'b10100:
        casez_tmp_191 = rob_val_3_20;
      5'b10101:
        casez_tmp_191 = rob_val_3_21;
      5'b10110:
        casez_tmp_191 = rob_val_3_22;
      5'b10111:
        casez_tmp_191 = rob_val_3_23;
      5'b11000:
        casez_tmp_191 = rob_val_3_24;
      5'b11001:
        casez_tmp_191 = rob_val_3_25;
      5'b11010:
        casez_tmp_191 = rob_val_3_26;
      5'b11011:
        casez_tmp_191 = rob_val_3_27;
      5'b11100:
        casez_tmp_191 = rob_val_3_28;
      5'b11101:
        casez_tmp_191 = rob_val_3_29;
      5'b11110:
        casez_tmp_191 = rob_val_3_30;
      default:
        casez_tmp_191 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1969 = _GEN_1382 & ~casez_tmp_191;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_192 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_192 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_192 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_192 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_192 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_192 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_192 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_192 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_192 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_192 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_192 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_192 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_192 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_192 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_192 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_192 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_192 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_192 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_192 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_192 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_192 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_192 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_192 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_192 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_192 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_192 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_192 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_192 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_192 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_192 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_192 = rob_bsy_3_30;
      default:
        casez_tmp_192 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1970 = _GEN_1382 & ~casez_tmp_192;
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_193 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_193 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_193 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_193 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_193 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_193 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_193 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_193 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_193 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_193 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_193 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_193 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_193 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_193 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_193 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_193 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_193 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_193 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_193 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_193 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_193 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_193 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_193 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_193 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_193 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_193 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_193 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_193 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_193 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_193 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_193 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_193 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_75)
      5'b00000:
        casez_tmp_194 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_194 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_194 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_194 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_194 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_194 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_194 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_194 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_194 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_194 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_194 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_194 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_194 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_194 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_194 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_194 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_194 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_194 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_194 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_194 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_194 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_194 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_194 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_194 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_194 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_194 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_194 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_194 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_194 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_194 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_194 = rob_uop_3_30_pdst;
      default:
        casez_tmp_194 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1971 = _GEN_1382 & casez_tmp_193 & casez_tmp_194 != io_wb_resps_7_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_195 = rob_val_3_0;
      5'b00001:
        casez_tmp_195 = rob_val_3_1;
      5'b00010:
        casez_tmp_195 = rob_val_3_2;
      5'b00011:
        casez_tmp_195 = rob_val_3_3;
      5'b00100:
        casez_tmp_195 = rob_val_3_4;
      5'b00101:
        casez_tmp_195 = rob_val_3_5;
      5'b00110:
        casez_tmp_195 = rob_val_3_6;
      5'b00111:
        casez_tmp_195 = rob_val_3_7;
      5'b01000:
        casez_tmp_195 = rob_val_3_8;
      5'b01001:
        casez_tmp_195 = rob_val_3_9;
      5'b01010:
        casez_tmp_195 = rob_val_3_10;
      5'b01011:
        casez_tmp_195 = rob_val_3_11;
      5'b01100:
        casez_tmp_195 = rob_val_3_12;
      5'b01101:
        casez_tmp_195 = rob_val_3_13;
      5'b01110:
        casez_tmp_195 = rob_val_3_14;
      5'b01111:
        casez_tmp_195 = rob_val_3_15;
      5'b10000:
        casez_tmp_195 = rob_val_3_16;
      5'b10001:
        casez_tmp_195 = rob_val_3_17;
      5'b10010:
        casez_tmp_195 = rob_val_3_18;
      5'b10011:
        casez_tmp_195 = rob_val_3_19;
      5'b10100:
        casez_tmp_195 = rob_val_3_20;
      5'b10101:
        casez_tmp_195 = rob_val_3_21;
      5'b10110:
        casez_tmp_195 = rob_val_3_22;
      5'b10111:
        casez_tmp_195 = rob_val_3_23;
      5'b11000:
        casez_tmp_195 = rob_val_3_24;
      5'b11001:
        casez_tmp_195 = rob_val_3_25;
      5'b11010:
        casez_tmp_195 = rob_val_3_26;
      5'b11011:
        casez_tmp_195 = rob_val_3_27;
      5'b11100:
        casez_tmp_195 = rob_val_3_28;
      5'b11101:
        casez_tmp_195 = rob_val_3_29;
      5'b11110:
        casez_tmp_195 = rob_val_3_30;
      default:
        casez_tmp_195 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1972 = _GEN_1838 & ~casez_tmp_195;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_196 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_196 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_196 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_196 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_196 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_196 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_196 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_196 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_196 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_196 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_196 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_196 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_196 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_196 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_196 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_196 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_196 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_196 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_196 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_196 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_196 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_196 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_196 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_196 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_196 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_196 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_196 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_196 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_196 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_196 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_196 = rob_bsy_3_30;
      default:
        casez_tmp_196 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1973 = _GEN_1838 & ~casez_tmp_196;
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_197 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_197 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_197 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_197 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_197 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_197 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_197 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_197 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_197 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_197 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_197 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_197 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_197 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_197 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_197 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_197 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_197 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_197 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_197 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_197 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_197 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_197 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_197 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_197 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_197 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_197 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_197 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_197 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_197 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_197 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_197 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_197 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_77)
      5'b00000:
        casez_tmp_198 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_198 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_198 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_198 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_198 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_198 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_198 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_198 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_198 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_198 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_198 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_198 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_198 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_198 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_198 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_198 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_198 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_198 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_198 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_198 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_198 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_198 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_198 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_198 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_198 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_198 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_198 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_198 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_198 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_198 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_198 = rob_uop_3_30_pdst;
      default:
        casez_tmp_198 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1974 = _GEN_1838 & casez_tmp_197 & casez_tmp_198 != io_wb_resps_8_bits_uop_pdst;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_199 = rob_val_3_0;
      5'b00001:
        casez_tmp_199 = rob_val_3_1;
      5'b00010:
        casez_tmp_199 = rob_val_3_2;
      5'b00011:
        casez_tmp_199 = rob_val_3_3;
      5'b00100:
        casez_tmp_199 = rob_val_3_4;
      5'b00101:
        casez_tmp_199 = rob_val_3_5;
      5'b00110:
        casez_tmp_199 = rob_val_3_6;
      5'b00111:
        casez_tmp_199 = rob_val_3_7;
      5'b01000:
        casez_tmp_199 = rob_val_3_8;
      5'b01001:
        casez_tmp_199 = rob_val_3_9;
      5'b01010:
        casez_tmp_199 = rob_val_3_10;
      5'b01011:
        casez_tmp_199 = rob_val_3_11;
      5'b01100:
        casez_tmp_199 = rob_val_3_12;
      5'b01101:
        casez_tmp_199 = rob_val_3_13;
      5'b01110:
        casez_tmp_199 = rob_val_3_14;
      5'b01111:
        casez_tmp_199 = rob_val_3_15;
      5'b10000:
        casez_tmp_199 = rob_val_3_16;
      5'b10001:
        casez_tmp_199 = rob_val_3_17;
      5'b10010:
        casez_tmp_199 = rob_val_3_18;
      5'b10011:
        casez_tmp_199 = rob_val_3_19;
      5'b10100:
        casez_tmp_199 = rob_val_3_20;
      5'b10101:
        casez_tmp_199 = rob_val_3_21;
      5'b10110:
        casez_tmp_199 = rob_val_3_22;
      5'b10111:
        casez_tmp_199 = rob_val_3_23;
      5'b11000:
        casez_tmp_199 = rob_val_3_24;
      5'b11001:
        casez_tmp_199 = rob_val_3_25;
      5'b11010:
        casez_tmp_199 = rob_val_3_26;
      5'b11011:
        casez_tmp_199 = rob_val_3_27;
      5'b11100:
        casez_tmp_199 = rob_val_3_28;
      5'b11101:
        casez_tmp_199 = rob_val_3_29;
      5'b11110:
        casez_tmp_199 = rob_val_3_30;
      default:
        casez_tmp_199 = rob_val_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1975 = _GEN_1381 & ~casez_tmp_199;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_200 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_200 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_200 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_200 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_200 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_200 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_200 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_200 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_200 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_200 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_200 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_200 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_200 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_200 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_200 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_200 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_200 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_200 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_200 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_200 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_200 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_200 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_200 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_200 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_200 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_200 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_200 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_200 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_200 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_200 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_200 = rob_bsy_3_30;
      default:
        casez_tmp_200 = rob_bsy_3_31;
    endcase
  end // always @(*)
  wire       _GEN_1976 = _GEN_1381 & ~casez_tmp_200;
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_201 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_201 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_201 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_201 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_201 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_201 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_201 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_201 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_201 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_201 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_201 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_201 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_201 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_201 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_201 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_201 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_201 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_201 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_201 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_201 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_201 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_201 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_201 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_201 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_201 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_201 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_201 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_201 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_201 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_201 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_201 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_201 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (_temp_uop_T_79)
      5'b00000:
        casez_tmp_202 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_202 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_202 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_202 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_202 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_202 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_202 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_202 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_202 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_202 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_202 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_202 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_202 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_202 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_202 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_202 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_202 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_202 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_202 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_202 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_202 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_202 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_202 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_202 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_202 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_202 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_202 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_202 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_202 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_202 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_202 = rob_uop_3_30_pdst;
      default:
        casez_tmp_202 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  wire       _GEN_1977 = _GEN_1381 & casez_tmp_201 & casez_tmp_202 != io_wb_resps_9_bits_uop_pdst;
  wire [2:0] _GEN_1978 = {1'h0, {1'h0, flush_commit_mask_0} + {1'h0, flush_commit_mask_1}} + {1'h0, {1'h0, flush_commit_mask_2} + {1'h0, flush_commit_mask_3}};
  wire       _GEN_1979 = _io_commit_valids_0_output & ~_rob_uop_com_idx_fp_val & (|rob_head_fflags_0);
  wire       _GEN_1980 = _fflags_val_0_T & (_io_commit_uops_0_uses_ldq_output | _io_commit_uops_0_uses_stq_output) & (|rob_head_fflags_0);
  wire       _GEN_1981 = _io_commit_valids_1_output & ~_rob_uop_1_com_idx_fp_val & (|rob_head_fflags_1);
  wire       _GEN_1982 = _fflags_val_1_T & (_io_commit_uops_1_uses_ldq_output | _io_commit_uops_1_uses_stq_output) & (|rob_head_fflags_1);
  wire       _GEN_1983 = _io_commit_valids_2_output & ~_rob_uop_2_com_idx_fp_val & (|rob_head_fflags_2);
  wire       _GEN_1984 = _fflags_val_2_T & (_io_commit_uops_2_uses_ldq_output | _io_commit_uops_2_uses_stq_output) & (|rob_head_fflags_2);
  wire       _GEN_1985 = _io_commit_valids_3_output & ~_rob_uop_3_com_idx_fp_val & (|rob_head_fflags_3);
  wire       _GEN_1986 = _fflags_val_3_T & (_io_commit_uops_3_uses_ldq_output | _io_commit_uops_3_uses_stq_output) & (|rob_head_fflags_3);
  wire       _GEN_1987 = exception_thrown & _io_ready_T_3;
  wire       _GEN_1988 = empty & r_xcpt_val;
  wire       _GEN_1989 = exception_thrown & r_xcpt_uop_rob_idx[6:2] != rob_head;
  reg        pnr_maybe_at_tail;
  wire       _GEN_1990 = rob_pnr_idx < rob_head_idx;
  wire       _GEN_1991 = _GEN_1990 ^ rob_head_idx < rob_tail_idx ^ rob_pnr_idx >= rob_tail_idx | rob_pnr_idx == rob_tail_idx;
  wire       _GEN_1992 = rob_tail_idx < rob_head_idx ^ _GEN_1990 ^ rob_tail_idx >= rob_pnr_idx | full;
  wire       _GEN_1993 = io_enq_valids_0 & ~reset;
  wire       _GEN_1994 = _GEN_1840 & ~reset;
  wire       _GEN_1995 = _GEN_3 & ~reset;
  wire       _GEN_1996 = _GEN_1841 & ~reset;
  wire       _GEN_1997 = _GEN_1842 & _GEN_1853 & ~reset;
  wire       _GEN_1998 = io_enq_valids_1 & ~reset;
  wire       _GEN_1999 = _GEN_1843 & ~reset;
  wire       _GEN_2000 = _GEN_462 & ~reset;
  wire       _GEN_2001 = _GEN_1844 & ~reset;
  wire       _GEN_2002 = _GEN_1845 & _GEN_1853 & ~reset;
  wire       _GEN_2003 = io_enq_valids_2 & ~reset;
  wire       _GEN_2004 = _GEN_1846 & ~reset;
  wire       _GEN_2005 = _GEN_921 & ~reset;
  wire       _GEN_2006 = _GEN_1847 & ~reset;
  wire       _GEN_2007 = _GEN_1848 & _GEN_1853 & ~reset;
  wire       _GEN_2008 = io_enq_valids_3 & ~reset;
  wire       _GEN_2009 = _GEN_1849 & ~reset;
  wire       _GEN_2010 = _GEN_1380 & ~reset;
  wire       _GEN_2011 = _GEN_1850 & ~reset;
  wire       _GEN_2012 = _GEN_1851 & _GEN_1853 & ~reset;
  `ifndef SYNTHESIS
    wire _GEN_2013 = (`PRINTF_COND_) & ~reset & _GEN_1854;
    always @(posedge clock) begin
      if ((`PRINTF_COND_) & _GEN_1993 & casez_tmp)
        $fwrite(32'h80000002, "Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1993 & ~_GEN_1852)
        $fwrite(32'h80000002, "Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
      if ((`PRINTF_COND_) & _GEN_1994 & ~casez_tmp_0)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1994 & ~casez_tmp_1)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1995 & ~casez_tmp_2)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1995 & ~casez_tmp_3)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1996 & ~casez_tmp_4)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1996 & ~casez_tmp_5)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1997 & ~casez_tmp_6)
        $fwrite(32'h80000002, "Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
      if (_GEN_2013)
        $fwrite(32'h80000002, "Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1855)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1856)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1857)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1858)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1859)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1860)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1861)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1862)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1863)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1864)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1865)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1866)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1867)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1868)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1869)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1870)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1871)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1872)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1873)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1874)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1875)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1876)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1877)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1878)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1879)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1880)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1881)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1882)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1883)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1884)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & _GEN_1998 & casez_tmp_50)
        $fwrite(32'h80000002, "Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1998 & ~_GEN_1885)
        $fwrite(32'h80000002, "Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
      if ((`PRINTF_COND_) & _GEN_1999 & ~casez_tmp_51)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_1999 & ~casez_tmp_52)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2000 & ~casez_tmp_53)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2000 & ~casez_tmp_54)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2001 & ~casez_tmp_55)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2001 & ~casez_tmp_56)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2002 & ~casez_tmp_57)
        $fwrite(32'h80000002, "Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
      if (_GEN_2013)
        $fwrite(32'h80000002, "Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1886)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1887)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1888)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1889)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1890)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1891)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1892)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1893)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1894)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1895)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1896)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1897)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1898)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1899)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1900)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1901)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1902)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1903)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1904)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1905)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1906)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1907)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1908)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1909)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1910)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1911)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1912)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1913)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1914)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1915)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & _GEN_2003 & casez_tmp_101)
        $fwrite(32'h80000002, "Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2003 & ~_GEN_1916)
        $fwrite(32'h80000002, "Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
      if ((`PRINTF_COND_) & _GEN_2004 & ~casez_tmp_102)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2004 & ~casez_tmp_103)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2005 & ~casez_tmp_104)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2005 & ~casez_tmp_105)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2006 & ~casez_tmp_106)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2006 & ~casez_tmp_107)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2007 & ~casez_tmp_108)
        $fwrite(32'h80000002, "Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
      if (_GEN_2013)
        $fwrite(32'h80000002, "Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1917)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1918)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1919)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1920)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1921)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1922)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1923)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1924)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1925)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1926)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1927)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1928)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1929)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1930)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1931)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1932)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1933)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1934)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1935)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1936)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1937)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1938)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1939)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1940)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1941)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1942)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1943)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1944)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1945)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1946)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & _GEN_2008 & casez_tmp_152)
        $fwrite(32'h80000002, "Assertion failed: [rob] overwriting a valid entry.\n    at rob.scala:333 assert (rob_val(rob_tail) === false.B, \"[rob] overwriting a valid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2008 & ~_GEN_1947)
        $fwrite(32'h80000002, "Assertion failed\n    at rob.scala:334 assert ((io.enq_uops(w).rob_idx >> log2Ceil(coreWidth)) === rob_tail)\n");
      if ((`PRINTF_COND_) & _GEN_2009 & ~casez_tmp_153)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2009 & ~casez_tmp_154)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2010 & ~casez_tmp_155)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2010 & ~casez_tmp_156)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2011 & ~casez_tmp_157)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to invalid entry.\n    at rob.scala:365 assert (rob_val(cidx) === true.B, \"[rob] store writing back to invalid entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2011 & ~casez_tmp_158)
        $fwrite(32'h80000002, "Assertion failed: [rob] store writing back to a not-busy entry.\n    at rob.scala:366 assert (rob_bsy(cidx) === true.B, \"[rob] store writing back to a not-busy entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_2012 & ~casez_tmp_159)
        $fwrite(32'h80000002, "Assertion failed: An instruction marked as safe is causing an exception\n    at rob.scala:394 assert(rob_unsafe(GetRowIdx(io.lxcpt.bits.uop.rob_idx)),\n");
      if (_GEN_2013)
        $fwrite(32'h80000002, "Assertion failed: com_valids and rbk_valids are mutually exclusive\n    at rob.scala:434 assert (!(io.commit.valids.reduce(_||_) && io.commit.rbk_valids.reduce(_||_)),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1948)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1949)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1950)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (0) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1951)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1952)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1953)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (1) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1954)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1955)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1956)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (2) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1957)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1958)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1959)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (3) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1960)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1961)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1962)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (4) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1963)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1964)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1965)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (5) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1966)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1967)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1968)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (6) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1969)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1970)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1971)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (7) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1972)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1973)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1974)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (8) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1975)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to an invalid ROB entry.\n    at rob.scala:518 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1976)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to a not-busy ROB entry.\n    at rob.scala:521 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1977)
        $fwrite(32'h80000002, "Assertion failed: [rob] writeback (9) occurred to the wrong pdst.\n    at rob.scala:524 assert (!(io.wb_resps(i).valid && MatchBank(GetBankIdx(rob_idx)) &&\n");
      if ((`PRINTF_COND_) & ~reset & (|(_GEN_1978[2:1])))
        $fwrite(32'h80000002, "Assertion failed: [rob] Can't commit multiple flush_on_commit instructions on one cycle\n    at rob.scala:580 assert(!(PopCount(flush_commit_mask) > 1.U),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1979)
        $fwrite(32'h80000002, "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1980)
        $fwrite(32'h80000002, "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1981)
        $fwrite(32'h80000002, "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1982)
        $fwrite(32'h80000002, "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1983)
        $fwrite(32'h80000002, "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1984)
        $fwrite(32'h80000002, "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1985)
        $fwrite(32'h80000002, "Assertion failed: Committed non-FP instruction has non-zero fflag bits.\n    at rob.scala:613 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1986)
        $fwrite(32'h80000002, "Assertion failed: Committed FP load or store has non-zero fflag bits.\n    at rob.scala:617 assert (!(io.commit.valids(w) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1987)
        $fwrite(32'h80000002, "Assertion failed: ROB trying to throw an exception, but it doesn't have a valid xcpt_cause\n    at rob.scala:667 assert (!(exception_thrown && !r_xcpt_val),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1988)
        $fwrite(32'h80000002, "Assertion failed: ROB is empty, but believes it has an outstanding exception.\n    at rob.scala:670 assert (!(empty && r_xcpt_val),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_1989)
        $fwrite(32'h80000002, "Assertion failed: ROB is throwing an exception, but the stored exception information's rob_idx does not match the rob_head\n    at rob.scala:673 assert (!(will_throw_exception && (GetRowIdx(r_xcpt_uop.rob_idx) =/= rob_head)),\n");
      if ((`PRINTF_COND_) & ~reset & ~_GEN_1991)
        $fwrite(32'h80000002, "Assertion failed\n    at rob.scala:749 assert(!IsOlder(rob_pnr_idx, rob_head_idx, rob_tail_idx) || rob_pnr_idx === rob_tail_idx)\n");
      if ((`PRINTF_COND_) & ~reset & ~_GEN_1992)
        $fwrite(32'h80000002, "Assertion failed\n    at rob.scala:752 assert(!IsOlder(rob_tail_idx, rob_pnr_idx, rob_head_idx) || full)\n");
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire [2:0] _GEN_2014 = {casez_tmp_101, casez_tmp_50, casez_tmp} | {casez_tmp_152, casez_tmp_101, casez_tmp_50};
  wire [1:0] _GEN_2015 = _GEN_2014[1:0] | {casez_tmp_152, casez_tmp_101};
  wire       safe_to_inc = _io_ready_T | (&rob_state);
  wire       rob_pnr_unsafe_0 = casez_tmp_9 & (casez_tmp_7 | casez_tmp_8);
  wire       rob_pnr_unsafe_1 = casez_tmp_60 & (casez_tmp_58 | casez_tmp_59);
  wire       rob_pnr_unsafe_2 = casez_tmp_111 & (casez_tmp_109 | casez_tmp_110);
  wire       _do_inc_row_T_4 = rob_pnr != rob_tail;
  wire       do_inc_row = ~(rob_pnr_unsafe_0 | rob_pnr_unsafe_1 | rob_pnr_unsafe_2 | casez_tmp_162 & (casez_tmp_160 | casez_tmp_161)) & (_do_inc_row_T_4 | full & ~pnr_maybe_at_tail);
  wire [2:0] _rob_pnr_lsb_T_16 = {rob_pnr_unsafe_2, rob_pnr_unsafe_1, rob_pnr_unsafe_0} | ~{_GEN_2014[2], _GEN_2015[1], _GEN_2015[0] | casez_tmp_152};
  wire       _rob_unsafe_rob_tail = io_enq_uops_0_uses_ldq | io_enq_uops_0_uses_stq & ~io_enq_uops_0_is_fence | io_enq_uops_0_is_br | io_enq_uops_0_is_jalr;
  wire       _GEN_2892 = _GEN_9 ? _rob_unsafe_rob_tail : rob_unsafe__0;
  wire       _GEN_2893 = _GEN_23 ? _rob_unsafe_rob_tail : rob_unsafe__1;
  wire       _GEN_2894 = _GEN_37 ? _rob_unsafe_rob_tail : rob_unsafe__2;
  wire       _GEN_2895 = _GEN_51 ? _rob_unsafe_rob_tail : rob_unsafe__3;
  wire       _GEN_2896 = _GEN_65 ? _rob_unsafe_rob_tail : rob_unsafe__4;
  wire       _GEN_2897 = _GEN_79 ? _rob_unsafe_rob_tail : rob_unsafe__5;
  wire       _GEN_2898 = _GEN_93 ? _rob_unsafe_rob_tail : rob_unsafe__6;
  wire       _GEN_2899 = _GEN_107 ? _rob_unsafe_rob_tail : rob_unsafe__7;
  wire       _GEN_2900 = _GEN_121 ? _rob_unsafe_rob_tail : rob_unsafe__8;
  wire       _GEN_2901 = _GEN_135 ? _rob_unsafe_rob_tail : rob_unsafe__9;
  wire       _GEN_2902 = _GEN_149 ? _rob_unsafe_rob_tail : rob_unsafe__10;
  wire       _GEN_2903 = _GEN_163 ? _rob_unsafe_rob_tail : rob_unsafe__11;
  wire       _GEN_2904 = _GEN_177 ? _rob_unsafe_rob_tail : rob_unsafe__12;
  wire       _GEN_2905 = _GEN_191 ? _rob_unsafe_rob_tail : rob_unsafe__13;
  wire       _GEN_2906 = _GEN_205 ? _rob_unsafe_rob_tail : rob_unsafe__14;
  wire       _GEN_2907 = _GEN_219 ? _rob_unsafe_rob_tail : rob_unsafe__15;
  wire       _GEN_2908 = _GEN_233 ? _rob_unsafe_rob_tail : rob_unsafe__16;
  wire       _GEN_2909 = _GEN_247 ? _rob_unsafe_rob_tail : rob_unsafe__17;
  wire       _GEN_2910 = _GEN_261 ? _rob_unsafe_rob_tail : rob_unsafe__18;
  wire       _GEN_2911 = _GEN_275 ? _rob_unsafe_rob_tail : rob_unsafe__19;
  wire       _GEN_2912 = _GEN_289 ? _rob_unsafe_rob_tail : rob_unsafe__20;
  wire       _GEN_2913 = _GEN_303 ? _rob_unsafe_rob_tail : rob_unsafe__21;
  wire       _GEN_2914 = _GEN_317 ? _rob_unsafe_rob_tail : rob_unsafe__22;
  wire       _GEN_2915 = _GEN_331 ? _rob_unsafe_rob_tail : rob_unsafe__23;
  wire       _GEN_2916 = _GEN_345 ? _rob_unsafe_rob_tail : rob_unsafe__24;
  wire       _GEN_2917 = _GEN_359 ? _rob_unsafe_rob_tail : rob_unsafe__25;
  wire       _GEN_2918 = _GEN_373 ? _rob_unsafe_rob_tail : rob_unsafe__26;
  wire       _GEN_2919 = _GEN_387 ? _rob_unsafe_rob_tail : rob_unsafe__27;
  wire       _GEN_2920 = _GEN_401 ? _rob_unsafe_rob_tail : rob_unsafe__28;
  wire       _GEN_2921 = _GEN_415 ? _rob_unsafe_rob_tail : rob_unsafe__29;
  wire       _GEN_2922 = _GEN_429 ? _rob_unsafe_rob_tail : rob_unsafe__30;
  wire       _GEN_2923 = _GEN_443 ? _rob_unsafe_rob_tail : rob_unsafe__31;
  wire       _GEN_5868 = _GEN_8 ? ~_GEN_11 & _GEN_2892 : ~_GEN_10 & _GEN_2892;
  wire       _GEN_5869 = _GEN_8 ? ~_GEN_25 & _GEN_2893 : ~_GEN_24 & _GEN_2893;
  wire       _GEN_5870 = _GEN_8 ? ~_GEN_39 & _GEN_2894 : ~_GEN_38 & _GEN_2894;
  wire       _GEN_5871 = _GEN_8 ? ~_GEN_53 & _GEN_2895 : ~_GEN_52 & _GEN_2895;
  wire       _GEN_5872 = _GEN_8 ? ~_GEN_67 & _GEN_2896 : ~_GEN_66 & _GEN_2896;
  wire       _GEN_5873 = _GEN_8 ? ~_GEN_81 & _GEN_2897 : ~_GEN_80 & _GEN_2897;
  wire       _GEN_5874 = _GEN_8 ? ~_GEN_95 & _GEN_2898 : ~_GEN_94 & _GEN_2898;
  wire       _GEN_5875 = _GEN_8 ? ~_GEN_109 & _GEN_2899 : ~_GEN_108 & _GEN_2899;
  wire       _GEN_5876 = _GEN_8 ? ~_GEN_123 & _GEN_2900 : ~_GEN_122 & _GEN_2900;
  wire       _GEN_5877 = _GEN_8 ? ~_GEN_137 & _GEN_2901 : ~_GEN_136 & _GEN_2901;
  wire       _GEN_5878 = _GEN_8 ? ~_GEN_151 & _GEN_2902 : ~_GEN_150 & _GEN_2902;
  wire       _GEN_5879 = _GEN_8 ? ~_GEN_165 & _GEN_2903 : ~_GEN_164 & _GEN_2903;
  wire       _GEN_5880 = _GEN_8 ? ~_GEN_179 & _GEN_2904 : ~_GEN_178 & _GEN_2904;
  wire       _GEN_5881 = _GEN_8 ? ~_GEN_193 & _GEN_2905 : ~_GEN_192 & _GEN_2905;
  wire       _GEN_5882 = _GEN_8 ? ~_GEN_207 & _GEN_2906 : ~_GEN_206 & _GEN_2906;
  wire       _GEN_5883 = _GEN_8 ? ~_GEN_221 & _GEN_2907 : ~_GEN_220 & _GEN_2907;
  wire       _GEN_5884 = _GEN_8 ? ~_GEN_235 & _GEN_2908 : ~_GEN_234 & _GEN_2908;
  wire       _GEN_5885 = _GEN_8 ? ~_GEN_249 & _GEN_2909 : ~_GEN_248 & _GEN_2909;
  wire       _GEN_5886 = _GEN_8 ? ~_GEN_263 & _GEN_2910 : ~_GEN_262 & _GEN_2910;
  wire       _GEN_5887 = _GEN_8 ? ~_GEN_277 & _GEN_2911 : ~_GEN_276 & _GEN_2911;
  wire       _GEN_5888 = _GEN_8 ? ~_GEN_291 & _GEN_2912 : ~_GEN_290 & _GEN_2912;
  wire       _GEN_5889 = _GEN_8 ? ~_GEN_305 & _GEN_2913 : ~_GEN_304 & _GEN_2913;
  wire       _GEN_5890 = _GEN_8 ? ~_GEN_319 & _GEN_2914 : ~_GEN_318 & _GEN_2914;
  wire       _GEN_5891 = _GEN_8 ? ~_GEN_333 & _GEN_2915 : ~_GEN_332 & _GEN_2915;
  wire       _GEN_5892 = _GEN_8 ? ~_GEN_347 & _GEN_2916 : ~_GEN_346 & _GEN_2916;
  wire       _GEN_5893 = _GEN_8 ? ~_GEN_361 & _GEN_2917 : ~_GEN_360 & _GEN_2917;
  wire       _GEN_5894 = _GEN_8 ? ~_GEN_375 & _GEN_2918 : ~_GEN_374 & _GEN_2918;
  wire       _GEN_5895 = _GEN_8 ? ~_GEN_389 & _GEN_2919 : ~_GEN_388 & _GEN_2919;
  wire       _GEN_5896 = _GEN_8 ? ~_GEN_403 & _GEN_2920 : ~_GEN_402 & _GEN_2920;
  wire       _GEN_5897 = _GEN_8 ? ~_GEN_417 & _GEN_2921 : ~_GEN_416 & _GEN_2921;
  wire       _GEN_5898 = _GEN_8 ? ~_GEN_431 & _GEN_2922 : ~_GEN_430 & _GEN_2922;
  wire       _GEN_5899 = _GEN_8 ? ~_GEN_445 & _GEN_2923 : ~_GEN_444 & _GEN_2923;
  wire       _GEN_6252 = _GEN_7 ? ~_GEN_13 & _GEN_5868 : ~_GEN_12 & _GEN_5868;
  wire       _GEN_6253 = _GEN_7 ? ~_GEN_27 & _GEN_5869 : ~_GEN_26 & _GEN_5869;
  wire       _GEN_6254 = _GEN_7 ? ~_GEN_41 & _GEN_5870 : ~_GEN_40 & _GEN_5870;
  wire       _GEN_6255 = _GEN_7 ? ~_GEN_55 & _GEN_5871 : ~_GEN_54 & _GEN_5871;
  wire       _GEN_6256 = _GEN_7 ? ~_GEN_69 & _GEN_5872 : ~_GEN_68 & _GEN_5872;
  wire       _GEN_6257 = _GEN_7 ? ~_GEN_83 & _GEN_5873 : ~_GEN_82 & _GEN_5873;
  wire       _GEN_6258 = _GEN_7 ? ~_GEN_97 & _GEN_5874 : ~_GEN_96 & _GEN_5874;
  wire       _GEN_6259 = _GEN_7 ? ~_GEN_111 & _GEN_5875 : ~_GEN_110 & _GEN_5875;
  wire       _GEN_6260 = _GEN_7 ? ~_GEN_125 & _GEN_5876 : ~_GEN_124 & _GEN_5876;
  wire       _GEN_6261 = _GEN_7 ? ~_GEN_139 & _GEN_5877 : ~_GEN_138 & _GEN_5877;
  wire       _GEN_6262 = _GEN_7 ? ~_GEN_153 & _GEN_5878 : ~_GEN_152 & _GEN_5878;
  wire       _GEN_6263 = _GEN_7 ? ~_GEN_167 & _GEN_5879 : ~_GEN_166 & _GEN_5879;
  wire       _GEN_6264 = _GEN_7 ? ~_GEN_181 & _GEN_5880 : ~_GEN_180 & _GEN_5880;
  wire       _GEN_6265 = _GEN_7 ? ~_GEN_195 & _GEN_5881 : ~_GEN_194 & _GEN_5881;
  wire       _GEN_6266 = _GEN_7 ? ~_GEN_209 & _GEN_5882 : ~_GEN_208 & _GEN_5882;
  wire       _GEN_6267 = _GEN_7 ? ~_GEN_223 & _GEN_5883 : ~_GEN_222 & _GEN_5883;
  wire       _GEN_6268 = _GEN_7 ? ~_GEN_237 & _GEN_5884 : ~_GEN_236 & _GEN_5884;
  wire       _GEN_6269 = _GEN_7 ? ~_GEN_251 & _GEN_5885 : ~_GEN_250 & _GEN_5885;
  wire       _GEN_6270 = _GEN_7 ? ~_GEN_265 & _GEN_5886 : ~_GEN_264 & _GEN_5886;
  wire       _GEN_6271 = _GEN_7 ? ~_GEN_279 & _GEN_5887 : ~_GEN_278 & _GEN_5887;
  wire       _GEN_6272 = _GEN_7 ? ~_GEN_293 & _GEN_5888 : ~_GEN_292 & _GEN_5888;
  wire       _GEN_6273 = _GEN_7 ? ~_GEN_307 & _GEN_5889 : ~_GEN_306 & _GEN_5889;
  wire       _GEN_6274 = _GEN_7 ? ~_GEN_321 & _GEN_5890 : ~_GEN_320 & _GEN_5890;
  wire       _GEN_6275 = _GEN_7 ? ~_GEN_335 & _GEN_5891 : ~_GEN_334 & _GEN_5891;
  wire       _GEN_6276 = _GEN_7 ? ~_GEN_349 & _GEN_5892 : ~_GEN_348 & _GEN_5892;
  wire       _GEN_6277 = _GEN_7 ? ~_GEN_363 & _GEN_5893 : ~_GEN_362 & _GEN_5893;
  wire       _GEN_6278 = _GEN_7 ? ~_GEN_377 & _GEN_5894 : ~_GEN_376 & _GEN_5894;
  wire       _GEN_6279 = _GEN_7 ? ~_GEN_391 & _GEN_5895 : ~_GEN_390 & _GEN_5895;
  wire       _GEN_6280 = _GEN_7 ? ~_GEN_405 & _GEN_5896 : ~_GEN_404 & _GEN_5896;
  wire       _GEN_6281 = _GEN_7 ? ~_GEN_419 & _GEN_5897 : ~_GEN_418 & _GEN_5897;
  wire       _GEN_6282 = _GEN_7 ? ~_GEN_433 & _GEN_5898 : ~_GEN_432 & _GEN_5898;
  wire       _GEN_6283 = _GEN_7 ? ~_GEN_447 & _GEN_5899 : ~_GEN_446 & _GEN_5899;
  wire       _GEN_6636 = _GEN_6 ? ~_GEN_15 & _GEN_6252 : ~_GEN_14 & _GEN_6252;
  wire       _GEN_6637 = _GEN_6 ? ~_GEN_29 & _GEN_6253 : ~_GEN_28 & _GEN_6253;
  wire       _GEN_6638 = _GEN_6 ? ~_GEN_43 & _GEN_6254 : ~_GEN_42 & _GEN_6254;
  wire       _GEN_6639 = _GEN_6 ? ~_GEN_57 & _GEN_6255 : ~_GEN_56 & _GEN_6255;
  wire       _GEN_6640 = _GEN_6 ? ~_GEN_71 & _GEN_6256 : ~_GEN_70 & _GEN_6256;
  wire       _GEN_6641 = _GEN_6 ? ~_GEN_85 & _GEN_6257 : ~_GEN_84 & _GEN_6257;
  wire       _GEN_6642 = _GEN_6 ? ~_GEN_99 & _GEN_6258 : ~_GEN_98 & _GEN_6258;
  wire       _GEN_6643 = _GEN_6 ? ~_GEN_113 & _GEN_6259 : ~_GEN_112 & _GEN_6259;
  wire       _GEN_6644 = _GEN_6 ? ~_GEN_127 & _GEN_6260 : ~_GEN_126 & _GEN_6260;
  wire       _GEN_6645 = _GEN_6 ? ~_GEN_141 & _GEN_6261 : ~_GEN_140 & _GEN_6261;
  wire       _GEN_6646 = _GEN_6 ? ~_GEN_155 & _GEN_6262 : ~_GEN_154 & _GEN_6262;
  wire       _GEN_6647 = _GEN_6 ? ~_GEN_169 & _GEN_6263 : ~_GEN_168 & _GEN_6263;
  wire       _GEN_6648 = _GEN_6 ? ~_GEN_183 & _GEN_6264 : ~_GEN_182 & _GEN_6264;
  wire       _GEN_6649 = _GEN_6 ? ~_GEN_197 & _GEN_6265 : ~_GEN_196 & _GEN_6265;
  wire       _GEN_6650 = _GEN_6 ? ~_GEN_211 & _GEN_6266 : ~_GEN_210 & _GEN_6266;
  wire       _GEN_6651 = _GEN_6 ? ~_GEN_225 & _GEN_6267 : ~_GEN_224 & _GEN_6267;
  wire       _GEN_6652 = _GEN_6 ? ~_GEN_239 & _GEN_6268 : ~_GEN_238 & _GEN_6268;
  wire       _GEN_6653 = _GEN_6 ? ~_GEN_253 & _GEN_6269 : ~_GEN_252 & _GEN_6269;
  wire       _GEN_6654 = _GEN_6 ? ~_GEN_267 & _GEN_6270 : ~_GEN_266 & _GEN_6270;
  wire       _GEN_6655 = _GEN_6 ? ~_GEN_281 & _GEN_6271 : ~_GEN_280 & _GEN_6271;
  wire       _GEN_6656 = _GEN_6 ? ~_GEN_295 & _GEN_6272 : ~_GEN_294 & _GEN_6272;
  wire       _GEN_6657 = _GEN_6 ? ~_GEN_309 & _GEN_6273 : ~_GEN_308 & _GEN_6273;
  wire       _GEN_6658 = _GEN_6 ? ~_GEN_323 & _GEN_6274 : ~_GEN_322 & _GEN_6274;
  wire       _GEN_6659 = _GEN_6 ? ~_GEN_337 & _GEN_6275 : ~_GEN_336 & _GEN_6275;
  wire       _GEN_6660 = _GEN_6 ? ~_GEN_351 & _GEN_6276 : ~_GEN_350 & _GEN_6276;
  wire       _GEN_6661 = _GEN_6 ? ~_GEN_365 & _GEN_6277 : ~_GEN_364 & _GEN_6277;
  wire       _GEN_6662 = _GEN_6 ? ~_GEN_379 & _GEN_6278 : ~_GEN_378 & _GEN_6278;
  wire       _GEN_6663 = _GEN_6 ? ~_GEN_393 & _GEN_6279 : ~_GEN_392 & _GEN_6279;
  wire       _GEN_6664 = _GEN_6 ? ~_GEN_407 & _GEN_6280 : ~_GEN_406 & _GEN_6280;
  wire       _GEN_6665 = _GEN_6 ? ~_GEN_421 & _GEN_6281 : ~_GEN_420 & _GEN_6281;
  wire       _GEN_6666 = _GEN_6 ? ~_GEN_435 & _GEN_6282 : ~_GEN_434 & _GEN_6282;
  wire       _GEN_6667 = _GEN_6 ? ~_GEN_449 & _GEN_6283 : ~_GEN_448 & _GEN_6283;
  wire       _GEN_7020 = _GEN_5 ? ~_GEN_17 & _GEN_6636 : ~_GEN_16 & _GEN_6636;
  wire       _GEN_7021 = _GEN_5 ? ~_GEN_31 & _GEN_6637 : ~_GEN_30 & _GEN_6637;
  wire       _GEN_7022 = _GEN_5 ? ~_GEN_45 & _GEN_6638 : ~_GEN_44 & _GEN_6638;
  wire       _GEN_7023 = _GEN_5 ? ~_GEN_59 & _GEN_6639 : ~_GEN_58 & _GEN_6639;
  wire       _GEN_7024 = _GEN_5 ? ~_GEN_73 & _GEN_6640 : ~_GEN_72 & _GEN_6640;
  wire       _GEN_7025 = _GEN_5 ? ~_GEN_87 & _GEN_6641 : ~_GEN_86 & _GEN_6641;
  wire       _GEN_7026 = _GEN_5 ? ~_GEN_101 & _GEN_6642 : ~_GEN_100 & _GEN_6642;
  wire       _GEN_7027 = _GEN_5 ? ~_GEN_115 & _GEN_6643 : ~_GEN_114 & _GEN_6643;
  wire       _GEN_7028 = _GEN_5 ? ~_GEN_129 & _GEN_6644 : ~_GEN_128 & _GEN_6644;
  wire       _GEN_7029 = _GEN_5 ? ~_GEN_143 & _GEN_6645 : ~_GEN_142 & _GEN_6645;
  wire       _GEN_7030 = _GEN_5 ? ~_GEN_157 & _GEN_6646 : ~_GEN_156 & _GEN_6646;
  wire       _GEN_7031 = _GEN_5 ? ~_GEN_171 & _GEN_6647 : ~_GEN_170 & _GEN_6647;
  wire       _GEN_7032 = _GEN_5 ? ~_GEN_185 & _GEN_6648 : ~_GEN_184 & _GEN_6648;
  wire       _GEN_7033 = _GEN_5 ? ~_GEN_199 & _GEN_6649 : ~_GEN_198 & _GEN_6649;
  wire       _GEN_7034 = _GEN_5 ? ~_GEN_213 & _GEN_6650 : ~_GEN_212 & _GEN_6650;
  wire       _GEN_7035 = _GEN_5 ? ~_GEN_227 & _GEN_6651 : ~_GEN_226 & _GEN_6651;
  wire       _GEN_7036 = _GEN_5 ? ~_GEN_241 & _GEN_6652 : ~_GEN_240 & _GEN_6652;
  wire       _GEN_7037 = _GEN_5 ? ~_GEN_255 & _GEN_6653 : ~_GEN_254 & _GEN_6653;
  wire       _GEN_7038 = _GEN_5 ? ~_GEN_269 & _GEN_6654 : ~_GEN_268 & _GEN_6654;
  wire       _GEN_7039 = _GEN_5 ? ~_GEN_283 & _GEN_6655 : ~_GEN_282 & _GEN_6655;
  wire       _GEN_7040 = _GEN_5 ? ~_GEN_297 & _GEN_6656 : ~_GEN_296 & _GEN_6656;
  wire       _GEN_7041 = _GEN_5 ? ~_GEN_311 & _GEN_6657 : ~_GEN_310 & _GEN_6657;
  wire       _GEN_7042 = _GEN_5 ? ~_GEN_325 & _GEN_6658 : ~_GEN_324 & _GEN_6658;
  wire       _GEN_7043 = _GEN_5 ? ~_GEN_339 & _GEN_6659 : ~_GEN_338 & _GEN_6659;
  wire       _GEN_7044 = _GEN_5 ? ~_GEN_353 & _GEN_6660 : ~_GEN_352 & _GEN_6660;
  wire       _GEN_7045 = _GEN_5 ? ~_GEN_367 & _GEN_6661 : ~_GEN_366 & _GEN_6661;
  wire       _GEN_7046 = _GEN_5 ? ~_GEN_381 & _GEN_6662 : ~_GEN_380 & _GEN_6662;
  wire       _GEN_7047 = _GEN_5 ? ~_GEN_395 & _GEN_6663 : ~_GEN_394 & _GEN_6663;
  wire       _GEN_7048 = _GEN_5 ? ~_GEN_409 & _GEN_6664 : ~_GEN_408 & _GEN_6664;
  wire       _GEN_7049 = _GEN_5 ? ~_GEN_423 & _GEN_6665 : ~_GEN_422 & _GEN_6665;
  wire       _GEN_7050 = _GEN_5 ? ~_GEN_437 & _GEN_6666 : ~_GEN_436 & _GEN_6666;
  wire       _GEN_7051 = _GEN_5 ? ~_GEN_451 & _GEN_6667 : ~_GEN_450 & _GEN_6667;
  wire       _GEN_7404 = _GEN_4 ? ~_GEN_19 & _GEN_7020 : ~_GEN_18 & _GEN_7020;
  wire       _GEN_7405 = _GEN_4 ? ~_GEN_33 & _GEN_7021 : ~_GEN_32 & _GEN_7021;
  wire       _GEN_7406 = _GEN_4 ? ~_GEN_47 & _GEN_7022 : ~_GEN_46 & _GEN_7022;
  wire       _GEN_7407 = _GEN_4 ? ~_GEN_61 & _GEN_7023 : ~_GEN_60 & _GEN_7023;
  wire       _GEN_7408 = _GEN_4 ? ~_GEN_75 & _GEN_7024 : ~_GEN_74 & _GEN_7024;
  wire       _GEN_7409 = _GEN_4 ? ~_GEN_89 & _GEN_7025 : ~_GEN_88 & _GEN_7025;
  wire       _GEN_7410 = _GEN_4 ? ~_GEN_103 & _GEN_7026 : ~_GEN_102 & _GEN_7026;
  wire       _GEN_7411 = _GEN_4 ? ~_GEN_117 & _GEN_7027 : ~_GEN_116 & _GEN_7027;
  wire       _GEN_7412 = _GEN_4 ? ~_GEN_131 & _GEN_7028 : ~_GEN_130 & _GEN_7028;
  wire       _GEN_7413 = _GEN_4 ? ~_GEN_145 & _GEN_7029 : ~_GEN_144 & _GEN_7029;
  wire       _GEN_7414 = _GEN_4 ? ~_GEN_159 & _GEN_7030 : ~_GEN_158 & _GEN_7030;
  wire       _GEN_7415 = _GEN_4 ? ~_GEN_173 & _GEN_7031 : ~_GEN_172 & _GEN_7031;
  wire       _GEN_7416 = _GEN_4 ? ~_GEN_187 & _GEN_7032 : ~_GEN_186 & _GEN_7032;
  wire       _GEN_7417 = _GEN_4 ? ~_GEN_201 & _GEN_7033 : ~_GEN_200 & _GEN_7033;
  wire       _GEN_7418 = _GEN_4 ? ~_GEN_215 & _GEN_7034 : ~_GEN_214 & _GEN_7034;
  wire       _GEN_7419 = _GEN_4 ? ~_GEN_229 & _GEN_7035 : ~_GEN_228 & _GEN_7035;
  wire       _GEN_7420 = _GEN_4 ? ~_GEN_243 & _GEN_7036 : ~_GEN_242 & _GEN_7036;
  wire       _GEN_7421 = _GEN_4 ? ~_GEN_257 & _GEN_7037 : ~_GEN_256 & _GEN_7037;
  wire       _GEN_7422 = _GEN_4 ? ~_GEN_271 & _GEN_7038 : ~_GEN_270 & _GEN_7038;
  wire       _GEN_7423 = _GEN_4 ? ~_GEN_285 & _GEN_7039 : ~_GEN_284 & _GEN_7039;
  wire       _GEN_7424 = _GEN_4 ? ~_GEN_299 & _GEN_7040 : ~_GEN_298 & _GEN_7040;
  wire       _GEN_7425 = _GEN_4 ? ~_GEN_313 & _GEN_7041 : ~_GEN_312 & _GEN_7041;
  wire       _GEN_7426 = _GEN_4 ? ~_GEN_327 & _GEN_7042 : ~_GEN_326 & _GEN_7042;
  wire       _GEN_7427 = _GEN_4 ? ~_GEN_341 & _GEN_7043 : ~_GEN_340 & _GEN_7043;
  wire       _GEN_7428 = _GEN_4 ? ~_GEN_355 & _GEN_7044 : ~_GEN_354 & _GEN_7044;
  wire       _GEN_7429 = _GEN_4 ? ~_GEN_369 & _GEN_7045 : ~_GEN_368 & _GEN_7045;
  wire       _GEN_7430 = _GEN_4 ? ~_GEN_383 & _GEN_7046 : ~_GEN_382 & _GEN_7046;
  wire       _GEN_7431 = _GEN_4 ? ~_GEN_397 & _GEN_7047 : ~_GEN_396 & _GEN_7047;
  wire       _GEN_7432 = _GEN_4 ? ~_GEN_411 & _GEN_7048 : ~_GEN_410 & _GEN_7048;
  wire       _GEN_7433 = _GEN_4 ? ~_GEN_425 & _GEN_7049 : ~_GEN_424 & _GEN_7049;
  wire       _GEN_7434 = _GEN_4 ? ~_GEN_439 & _GEN_7050 : ~_GEN_438 & _GEN_7050;
  wire       _GEN_7435 = _GEN_4 ? ~_GEN_453 & _GEN_7051 : ~_GEN_452 & _GEN_7051;
  wire       _rob_unsafe_1_rob_tail = io_enq_uops_1_uses_ldq | io_enq_uops_1_uses_stq & ~io_enq_uops_1_is_fence | io_enq_uops_1_is_br | io_enq_uops_1_is_jalr;
  wire       _GEN_16256 = _GEN_468 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_0;
  wire       _GEN_16257 = _GEN_482 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_1;
  wire       _GEN_16258 = _GEN_496 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_2;
  wire       _GEN_16259 = _GEN_510 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_3;
  wire       _GEN_16260 = _GEN_524 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_4;
  wire       _GEN_16261 = _GEN_538 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_5;
  wire       _GEN_16262 = _GEN_552 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_6;
  wire       _GEN_16263 = _GEN_566 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_7;
  wire       _GEN_16264 = _GEN_580 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_8;
  wire       _GEN_16265 = _GEN_594 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_9;
  wire       _GEN_16266 = _GEN_608 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_10;
  wire       _GEN_16267 = _GEN_622 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_11;
  wire       _GEN_16268 = _GEN_636 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_12;
  wire       _GEN_16269 = _GEN_650 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_13;
  wire       _GEN_16270 = _GEN_664 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_14;
  wire       _GEN_16271 = _GEN_678 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_15;
  wire       _GEN_16272 = _GEN_692 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_16;
  wire       _GEN_16273 = _GEN_706 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_17;
  wire       _GEN_16274 = _GEN_720 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_18;
  wire       _GEN_16275 = _GEN_734 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_19;
  wire       _GEN_16276 = _GEN_748 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_20;
  wire       _GEN_16277 = _GEN_762 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_21;
  wire       _GEN_16278 = _GEN_776 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_22;
  wire       _GEN_16279 = _GEN_790 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_23;
  wire       _GEN_16280 = _GEN_804 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_24;
  wire       _GEN_16281 = _GEN_818 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_25;
  wire       _GEN_16282 = _GEN_832 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_26;
  wire       _GEN_16283 = _GEN_846 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_27;
  wire       _GEN_16284 = _GEN_860 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_28;
  wire       _GEN_16285 = _GEN_874 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_29;
  wire       _GEN_16286 = _GEN_888 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_30;
  wire       _GEN_16287 = _GEN_902 ? _rob_unsafe_1_rob_tail : rob_unsafe_1_31;
  wire       _GEN_19232 = _GEN_467 ? ~_GEN_470 & _GEN_16256 : ~_GEN_469 & _GEN_16256;
  wire       _GEN_19233 = _GEN_467 ? ~_GEN_484 & _GEN_16257 : ~_GEN_483 & _GEN_16257;
  wire       _GEN_19234 = _GEN_467 ? ~_GEN_498 & _GEN_16258 : ~_GEN_497 & _GEN_16258;
  wire       _GEN_19235 = _GEN_467 ? ~_GEN_512 & _GEN_16259 : ~_GEN_511 & _GEN_16259;
  wire       _GEN_19236 = _GEN_467 ? ~_GEN_526 & _GEN_16260 : ~_GEN_525 & _GEN_16260;
  wire       _GEN_19237 = _GEN_467 ? ~_GEN_540 & _GEN_16261 : ~_GEN_539 & _GEN_16261;
  wire       _GEN_19238 = _GEN_467 ? ~_GEN_554 & _GEN_16262 : ~_GEN_553 & _GEN_16262;
  wire       _GEN_19239 = _GEN_467 ? ~_GEN_568 & _GEN_16263 : ~_GEN_567 & _GEN_16263;
  wire       _GEN_19240 = _GEN_467 ? ~_GEN_582 & _GEN_16264 : ~_GEN_581 & _GEN_16264;
  wire       _GEN_19241 = _GEN_467 ? ~_GEN_596 & _GEN_16265 : ~_GEN_595 & _GEN_16265;
  wire       _GEN_19242 = _GEN_467 ? ~_GEN_610 & _GEN_16266 : ~_GEN_609 & _GEN_16266;
  wire       _GEN_19243 = _GEN_467 ? ~_GEN_624 & _GEN_16267 : ~_GEN_623 & _GEN_16267;
  wire       _GEN_19244 = _GEN_467 ? ~_GEN_638 & _GEN_16268 : ~_GEN_637 & _GEN_16268;
  wire       _GEN_19245 = _GEN_467 ? ~_GEN_652 & _GEN_16269 : ~_GEN_651 & _GEN_16269;
  wire       _GEN_19246 = _GEN_467 ? ~_GEN_666 & _GEN_16270 : ~_GEN_665 & _GEN_16270;
  wire       _GEN_19247 = _GEN_467 ? ~_GEN_680 & _GEN_16271 : ~_GEN_679 & _GEN_16271;
  wire       _GEN_19248 = _GEN_467 ? ~_GEN_694 & _GEN_16272 : ~_GEN_693 & _GEN_16272;
  wire       _GEN_19249 = _GEN_467 ? ~_GEN_708 & _GEN_16273 : ~_GEN_707 & _GEN_16273;
  wire       _GEN_19250 = _GEN_467 ? ~_GEN_722 & _GEN_16274 : ~_GEN_721 & _GEN_16274;
  wire       _GEN_19251 = _GEN_467 ? ~_GEN_736 & _GEN_16275 : ~_GEN_735 & _GEN_16275;
  wire       _GEN_19252 = _GEN_467 ? ~_GEN_750 & _GEN_16276 : ~_GEN_749 & _GEN_16276;
  wire       _GEN_19253 = _GEN_467 ? ~_GEN_764 & _GEN_16277 : ~_GEN_763 & _GEN_16277;
  wire       _GEN_19254 = _GEN_467 ? ~_GEN_778 & _GEN_16278 : ~_GEN_777 & _GEN_16278;
  wire       _GEN_19255 = _GEN_467 ? ~_GEN_792 & _GEN_16279 : ~_GEN_791 & _GEN_16279;
  wire       _GEN_19256 = _GEN_467 ? ~_GEN_806 & _GEN_16280 : ~_GEN_805 & _GEN_16280;
  wire       _GEN_19257 = _GEN_467 ? ~_GEN_820 & _GEN_16281 : ~_GEN_819 & _GEN_16281;
  wire       _GEN_19258 = _GEN_467 ? ~_GEN_834 & _GEN_16282 : ~_GEN_833 & _GEN_16282;
  wire       _GEN_19259 = _GEN_467 ? ~_GEN_848 & _GEN_16283 : ~_GEN_847 & _GEN_16283;
  wire       _GEN_19260 = _GEN_467 ? ~_GEN_862 & _GEN_16284 : ~_GEN_861 & _GEN_16284;
  wire       _GEN_19261 = _GEN_467 ? ~_GEN_876 & _GEN_16285 : ~_GEN_875 & _GEN_16285;
  wire       _GEN_19262 = _GEN_467 ? ~_GEN_890 & _GEN_16286 : ~_GEN_889 & _GEN_16286;
  wire       _GEN_19263 = _GEN_467 ? ~_GEN_904 & _GEN_16287 : ~_GEN_903 & _GEN_16287;
  wire       _GEN_19616 = _GEN_466 ? ~_GEN_472 & _GEN_19232 : ~_GEN_471 & _GEN_19232;
  wire       _GEN_19617 = _GEN_466 ? ~_GEN_486 & _GEN_19233 : ~_GEN_485 & _GEN_19233;
  wire       _GEN_19618 = _GEN_466 ? ~_GEN_500 & _GEN_19234 : ~_GEN_499 & _GEN_19234;
  wire       _GEN_19619 = _GEN_466 ? ~_GEN_514 & _GEN_19235 : ~_GEN_513 & _GEN_19235;
  wire       _GEN_19620 = _GEN_466 ? ~_GEN_528 & _GEN_19236 : ~_GEN_527 & _GEN_19236;
  wire       _GEN_19621 = _GEN_466 ? ~_GEN_542 & _GEN_19237 : ~_GEN_541 & _GEN_19237;
  wire       _GEN_19622 = _GEN_466 ? ~_GEN_556 & _GEN_19238 : ~_GEN_555 & _GEN_19238;
  wire       _GEN_19623 = _GEN_466 ? ~_GEN_570 & _GEN_19239 : ~_GEN_569 & _GEN_19239;
  wire       _GEN_19624 = _GEN_466 ? ~_GEN_584 & _GEN_19240 : ~_GEN_583 & _GEN_19240;
  wire       _GEN_19625 = _GEN_466 ? ~_GEN_598 & _GEN_19241 : ~_GEN_597 & _GEN_19241;
  wire       _GEN_19626 = _GEN_466 ? ~_GEN_612 & _GEN_19242 : ~_GEN_611 & _GEN_19242;
  wire       _GEN_19627 = _GEN_466 ? ~_GEN_626 & _GEN_19243 : ~_GEN_625 & _GEN_19243;
  wire       _GEN_19628 = _GEN_466 ? ~_GEN_640 & _GEN_19244 : ~_GEN_639 & _GEN_19244;
  wire       _GEN_19629 = _GEN_466 ? ~_GEN_654 & _GEN_19245 : ~_GEN_653 & _GEN_19245;
  wire       _GEN_19630 = _GEN_466 ? ~_GEN_668 & _GEN_19246 : ~_GEN_667 & _GEN_19246;
  wire       _GEN_19631 = _GEN_466 ? ~_GEN_682 & _GEN_19247 : ~_GEN_681 & _GEN_19247;
  wire       _GEN_19632 = _GEN_466 ? ~_GEN_696 & _GEN_19248 : ~_GEN_695 & _GEN_19248;
  wire       _GEN_19633 = _GEN_466 ? ~_GEN_710 & _GEN_19249 : ~_GEN_709 & _GEN_19249;
  wire       _GEN_19634 = _GEN_466 ? ~_GEN_724 & _GEN_19250 : ~_GEN_723 & _GEN_19250;
  wire       _GEN_19635 = _GEN_466 ? ~_GEN_738 & _GEN_19251 : ~_GEN_737 & _GEN_19251;
  wire       _GEN_19636 = _GEN_466 ? ~_GEN_752 & _GEN_19252 : ~_GEN_751 & _GEN_19252;
  wire       _GEN_19637 = _GEN_466 ? ~_GEN_766 & _GEN_19253 : ~_GEN_765 & _GEN_19253;
  wire       _GEN_19638 = _GEN_466 ? ~_GEN_780 & _GEN_19254 : ~_GEN_779 & _GEN_19254;
  wire       _GEN_19639 = _GEN_466 ? ~_GEN_794 & _GEN_19255 : ~_GEN_793 & _GEN_19255;
  wire       _GEN_19640 = _GEN_466 ? ~_GEN_808 & _GEN_19256 : ~_GEN_807 & _GEN_19256;
  wire       _GEN_19641 = _GEN_466 ? ~_GEN_822 & _GEN_19257 : ~_GEN_821 & _GEN_19257;
  wire       _GEN_19642 = _GEN_466 ? ~_GEN_836 & _GEN_19258 : ~_GEN_835 & _GEN_19258;
  wire       _GEN_19643 = _GEN_466 ? ~_GEN_850 & _GEN_19259 : ~_GEN_849 & _GEN_19259;
  wire       _GEN_19644 = _GEN_466 ? ~_GEN_864 & _GEN_19260 : ~_GEN_863 & _GEN_19260;
  wire       _GEN_19645 = _GEN_466 ? ~_GEN_878 & _GEN_19261 : ~_GEN_877 & _GEN_19261;
  wire       _GEN_19646 = _GEN_466 ? ~_GEN_892 & _GEN_19262 : ~_GEN_891 & _GEN_19262;
  wire       _GEN_19647 = _GEN_466 ? ~_GEN_906 & _GEN_19263 : ~_GEN_905 & _GEN_19263;
  wire       _GEN_20000 = _GEN_465 ? ~_GEN_474 & _GEN_19616 : ~_GEN_473 & _GEN_19616;
  wire       _GEN_20001 = _GEN_465 ? ~_GEN_488 & _GEN_19617 : ~_GEN_487 & _GEN_19617;
  wire       _GEN_20002 = _GEN_465 ? ~_GEN_502 & _GEN_19618 : ~_GEN_501 & _GEN_19618;
  wire       _GEN_20003 = _GEN_465 ? ~_GEN_516 & _GEN_19619 : ~_GEN_515 & _GEN_19619;
  wire       _GEN_20004 = _GEN_465 ? ~_GEN_530 & _GEN_19620 : ~_GEN_529 & _GEN_19620;
  wire       _GEN_20005 = _GEN_465 ? ~_GEN_544 & _GEN_19621 : ~_GEN_543 & _GEN_19621;
  wire       _GEN_20006 = _GEN_465 ? ~_GEN_558 & _GEN_19622 : ~_GEN_557 & _GEN_19622;
  wire       _GEN_20007 = _GEN_465 ? ~_GEN_572 & _GEN_19623 : ~_GEN_571 & _GEN_19623;
  wire       _GEN_20008 = _GEN_465 ? ~_GEN_586 & _GEN_19624 : ~_GEN_585 & _GEN_19624;
  wire       _GEN_20009 = _GEN_465 ? ~_GEN_600 & _GEN_19625 : ~_GEN_599 & _GEN_19625;
  wire       _GEN_20010 = _GEN_465 ? ~_GEN_614 & _GEN_19626 : ~_GEN_613 & _GEN_19626;
  wire       _GEN_20011 = _GEN_465 ? ~_GEN_628 & _GEN_19627 : ~_GEN_627 & _GEN_19627;
  wire       _GEN_20012 = _GEN_465 ? ~_GEN_642 & _GEN_19628 : ~_GEN_641 & _GEN_19628;
  wire       _GEN_20013 = _GEN_465 ? ~_GEN_656 & _GEN_19629 : ~_GEN_655 & _GEN_19629;
  wire       _GEN_20014 = _GEN_465 ? ~_GEN_670 & _GEN_19630 : ~_GEN_669 & _GEN_19630;
  wire       _GEN_20015 = _GEN_465 ? ~_GEN_684 & _GEN_19631 : ~_GEN_683 & _GEN_19631;
  wire       _GEN_20016 = _GEN_465 ? ~_GEN_698 & _GEN_19632 : ~_GEN_697 & _GEN_19632;
  wire       _GEN_20017 = _GEN_465 ? ~_GEN_712 & _GEN_19633 : ~_GEN_711 & _GEN_19633;
  wire       _GEN_20018 = _GEN_465 ? ~_GEN_726 & _GEN_19634 : ~_GEN_725 & _GEN_19634;
  wire       _GEN_20019 = _GEN_465 ? ~_GEN_740 & _GEN_19635 : ~_GEN_739 & _GEN_19635;
  wire       _GEN_20020 = _GEN_465 ? ~_GEN_754 & _GEN_19636 : ~_GEN_753 & _GEN_19636;
  wire       _GEN_20021 = _GEN_465 ? ~_GEN_768 & _GEN_19637 : ~_GEN_767 & _GEN_19637;
  wire       _GEN_20022 = _GEN_465 ? ~_GEN_782 & _GEN_19638 : ~_GEN_781 & _GEN_19638;
  wire       _GEN_20023 = _GEN_465 ? ~_GEN_796 & _GEN_19639 : ~_GEN_795 & _GEN_19639;
  wire       _GEN_20024 = _GEN_465 ? ~_GEN_810 & _GEN_19640 : ~_GEN_809 & _GEN_19640;
  wire       _GEN_20025 = _GEN_465 ? ~_GEN_824 & _GEN_19641 : ~_GEN_823 & _GEN_19641;
  wire       _GEN_20026 = _GEN_465 ? ~_GEN_838 & _GEN_19642 : ~_GEN_837 & _GEN_19642;
  wire       _GEN_20027 = _GEN_465 ? ~_GEN_852 & _GEN_19643 : ~_GEN_851 & _GEN_19643;
  wire       _GEN_20028 = _GEN_465 ? ~_GEN_866 & _GEN_19644 : ~_GEN_865 & _GEN_19644;
  wire       _GEN_20029 = _GEN_465 ? ~_GEN_880 & _GEN_19645 : ~_GEN_879 & _GEN_19645;
  wire       _GEN_20030 = _GEN_465 ? ~_GEN_894 & _GEN_19646 : ~_GEN_893 & _GEN_19646;
  wire       _GEN_20031 = _GEN_465 ? ~_GEN_908 & _GEN_19647 : ~_GEN_907 & _GEN_19647;
  wire       _GEN_20384 = _GEN_464 ? ~_GEN_476 & _GEN_20000 : ~_GEN_475 & _GEN_20000;
  wire       _GEN_20385 = _GEN_464 ? ~_GEN_490 & _GEN_20001 : ~_GEN_489 & _GEN_20001;
  wire       _GEN_20386 = _GEN_464 ? ~_GEN_504 & _GEN_20002 : ~_GEN_503 & _GEN_20002;
  wire       _GEN_20387 = _GEN_464 ? ~_GEN_518 & _GEN_20003 : ~_GEN_517 & _GEN_20003;
  wire       _GEN_20388 = _GEN_464 ? ~_GEN_532 & _GEN_20004 : ~_GEN_531 & _GEN_20004;
  wire       _GEN_20389 = _GEN_464 ? ~_GEN_546 & _GEN_20005 : ~_GEN_545 & _GEN_20005;
  wire       _GEN_20390 = _GEN_464 ? ~_GEN_560 & _GEN_20006 : ~_GEN_559 & _GEN_20006;
  wire       _GEN_20391 = _GEN_464 ? ~_GEN_574 & _GEN_20007 : ~_GEN_573 & _GEN_20007;
  wire       _GEN_20392 = _GEN_464 ? ~_GEN_588 & _GEN_20008 : ~_GEN_587 & _GEN_20008;
  wire       _GEN_20393 = _GEN_464 ? ~_GEN_602 & _GEN_20009 : ~_GEN_601 & _GEN_20009;
  wire       _GEN_20394 = _GEN_464 ? ~_GEN_616 & _GEN_20010 : ~_GEN_615 & _GEN_20010;
  wire       _GEN_20395 = _GEN_464 ? ~_GEN_630 & _GEN_20011 : ~_GEN_629 & _GEN_20011;
  wire       _GEN_20396 = _GEN_464 ? ~_GEN_644 & _GEN_20012 : ~_GEN_643 & _GEN_20012;
  wire       _GEN_20397 = _GEN_464 ? ~_GEN_658 & _GEN_20013 : ~_GEN_657 & _GEN_20013;
  wire       _GEN_20398 = _GEN_464 ? ~_GEN_672 & _GEN_20014 : ~_GEN_671 & _GEN_20014;
  wire       _GEN_20399 = _GEN_464 ? ~_GEN_686 & _GEN_20015 : ~_GEN_685 & _GEN_20015;
  wire       _GEN_20400 = _GEN_464 ? ~_GEN_700 & _GEN_20016 : ~_GEN_699 & _GEN_20016;
  wire       _GEN_20401 = _GEN_464 ? ~_GEN_714 & _GEN_20017 : ~_GEN_713 & _GEN_20017;
  wire       _GEN_20402 = _GEN_464 ? ~_GEN_728 & _GEN_20018 : ~_GEN_727 & _GEN_20018;
  wire       _GEN_20403 = _GEN_464 ? ~_GEN_742 & _GEN_20019 : ~_GEN_741 & _GEN_20019;
  wire       _GEN_20404 = _GEN_464 ? ~_GEN_756 & _GEN_20020 : ~_GEN_755 & _GEN_20020;
  wire       _GEN_20405 = _GEN_464 ? ~_GEN_770 & _GEN_20021 : ~_GEN_769 & _GEN_20021;
  wire       _GEN_20406 = _GEN_464 ? ~_GEN_784 & _GEN_20022 : ~_GEN_783 & _GEN_20022;
  wire       _GEN_20407 = _GEN_464 ? ~_GEN_798 & _GEN_20023 : ~_GEN_797 & _GEN_20023;
  wire       _GEN_20408 = _GEN_464 ? ~_GEN_812 & _GEN_20024 : ~_GEN_811 & _GEN_20024;
  wire       _GEN_20409 = _GEN_464 ? ~_GEN_826 & _GEN_20025 : ~_GEN_825 & _GEN_20025;
  wire       _GEN_20410 = _GEN_464 ? ~_GEN_840 & _GEN_20026 : ~_GEN_839 & _GEN_20026;
  wire       _GEN_20411 = _GEN_464 ? ~_GEN_854 & _GEN_20027 : ~_GEN_853 & _GEN_20027;
  wire       _GEN_20412 = _GEN_464 ? ~_GEN_868 & _GEN_20028 : ~_GEN_867 & _GEN_20028;
  wire       _GEN_20413 = _GEN_464 ? ~_GEN_882 & _GEN_20029 : ~_GEN_881 & _GEN_20029;
  wire       _GEN_20414 = _GEN_464 ? ~_GEN_896 & _GEN_20030 : ~_GEN_895 & _GEN_20030;
  wire       _GEN_20415 = _GEN_464 ? ~_GEN_910 & _GEN_20031 : ~_GEN_909 & _GEN_20031;
  wire       _GEN_20768 = _GEN_463 ? ~_GEN_478 & _GEN_20384 : ~_GEN_477 & _GEN_20384;
  wire       _GEN_20769 = _GEN_463 ? ~_GEN_492 & _GEN_20385 : ~_GEN_491 & _GEN_20385;
  wire       _GEN_20770 = _GEN_463 ? ~_GEN_506 & _GEN_20386 : ~_GEN_505 & _GEN_20386;
  wire       _GEN_20771 = _GEN_463 ? ~_GEN_520 & _GEN_20387 : ~_GEN_519 & _GEN_20387;
  wire       _GEN_20772 = _GEN_463 ? ~_GEN_534 & _GEN_20388 : ~_GEN_533 & _GEN_20388;
  wire       _GEN_20773 = _GEN_463 ? ~_GEN_548 & _GEN_20389 : ~_GEN_547 & _GEN_20389;
  wire       _GEN_20774 = _GEN_463 ? ~_GEN_562 & _GEN_20390 : ~_GEN_561 & _GEN_20390;
  wire       _GEN_20775 = _GEN_463 ? ~_GEN_576 & _GEN_20391 : ~_GEN_575 & _GEN_20391;
  wire       _GEN_20776 = _GEN_463 ? ~_GEN_590 & _GEN_20392 : ~_GEN_589 & _GEN_20392;
  wire       _GEN_20777 = _GEN_463 ? ~_GEN_604 & _GEN_20393 : ~_GEN_603 & _GEN_20393;
  wire       _GEN_20778 = _GEN_463 ? ~_GEN_618 & _GEN_20394 : ~_GEN_617 & _GEN_20394;
  wire       _GEN_20779 = _GEN_463 ? ~_GEN_632 & _GEN_20395 : ~_GEN_631 & _GEN_20395;
  wire       _GEN_20780 = _GEN_463 ? ~_GEN_646 & _GEN_20396 : ~_GEN_645 & _GEN_20396;
  wire       _GEN_20781 = _GEN_463 ? ~_GEN_660 & _GEN_20397 : ~_GEN_659 & _GEN_20397;
  wire       _GEN_20782 = _GEN_463 ? ~_GEN_674 & _GEN_20398 : ~_GEN_673 & _GEN_20398;
  wire       _GEN_20783 = _GEN_463 ? ~_GEN_688 & _GEN_20399 : ~_GEN_687 & _GEN_20399;
  wire       _GEN_20784 = _GEN_463 ? ~_GEN_702 & _GEN_20400 : ~_GEN_701 & _GEN_20400;
  wire       _GEN_20785 = _GEN_463 ? ~_GEN_716 & _GEN_20401 : ~_GEN_715 & _GEN_20401;
  wire       _GEN_20786 = _GEN_463 ? ~_GEN_730 & _GEN_20402 : ~_GEN_729 & _GEN_20402;
  wire       _GEN_20787 = _GEN_463 ? ~_GEN_744 & _GEN_20403 : ~_GEN_743 & _GEN_20403;
  wire       _GEN_20788 = _GEN_463 ? ~_GEN_758 & _GEN_20404 : ~_GEN_757 & _GEN_20404;
  wire       _GEN_20789 = _GEN_463 ? ~_GEN_772 & _GEN_20405 : ~_GEN_771 & _GEN_20405;
  wire       _GEN_20790 = _GEN_463 ? ~_GEN_786 & _GEN_20406 : ~_GEN_785 & _GEN_20406;
  wire       _GEN_20791 = _GEN_463 ? ~_GEN_800 & _GEN_20407 : ~_GEN_799 & _GEN_20407;
  wire       _GEN_20792 = _GEN_463 ? ~_GEN_814 & _GEN_20408 : ~_GEN_813 & _GEN_20408;
  wire       _GEN_20793 = _GEN_463 ? ~_GEN_828 & _GEN_20409 : ~_GEN_827 & _GEN_20409;
  wire       _GEN_20794 = _GEN_463 ? ~_GEN_842 & _GEN_20410 : ~_GEN_841 & _GEN_20410;
  wire       _GEN_20795 = _GEN_463 ? ~_GEN_856 & _GEN_20411 : ~_GEN_855 & _GEN_20411;
  wire       _GEN_20796 = _GEN_463 ? ~_GEN_870 & _GEN_20412 : ~_GEN_869 & _GEN_20412;
  wire       _GEN_20797 = _GEN_463 ? ~_GEN_884 & _GEN_20413 : ~_GEN_883 & _GEN_20413;
  wire       _GEN_20798 = _GEN_463 ? ~_GEN_898 & _GEN_20414 : ~_GEN_897 & _GEN_20414;
  wire       _GEN_20799 = _GEN_463 ? ~_GEN_912 & _GEN_20415 : ~_GEN_911 & _GEN_20415;
  wire       _rob_unsafe_2_rob_tail = io_enq_uops_2_uses_ldq | io_enq_uops_2_uses_stq & ~io_enq_uops_2_is_fence | io_enq_uops_2_is_br | io_enq_uops_2_is_jalr;
  wire       _GEN_29620 = _GEN_927 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_0;
  wire       _GEN_29621 = _GEN_941 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_1;
  wire       _GEN_29622 = _GEN_955 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_2;
  wire       _GEN_29623 = _GEN_969 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_3;
  wire       _GEN_29624 = _GEN_983 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_4;
  wire       _GEN_29625 = _GEN_997 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_5;
  wire       _GEN_29626 = _GEN_1011 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_6;
  wire       _GEN_29627 = _GEN_1025 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_7;
  wire       _GEN_29628 = _GEN_1039 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_8;
  wire       _GEN_29629 = _GEN_1053 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_9;
  wire       _GEN_29630 = _GEN_1067 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_10;
  wire       _GEN_29631 = _GEN_1081 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_11;
  wire       _GEN_29632 = _GEN_1095 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_12;
  wire       _GEN_29633 = _GEN_1109 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_13;
  wire       _GEN_29634 = _GEN_1123 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_14;
  wire       _GEN_29635 = _GEN_1137 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_15;
  wire       _GEN_29636 = _GEN_1151 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_16;
  wire       _GEN_29637 = _GEN_1165 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_17;
  wire       _GEN_29638 = _GEN_1179 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_18;
  wire       _GEN_29639 = _GEN_1193 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_19;
  wire       _GEN_29640 = _GEN_1207 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_20;
  wire       _GEN_29641 = _GEN_1221 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_21;
  wire       _GEN_29642 = _GEN_1235 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_22;
  wire       _GEN_29643 = _GEN_1249 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_23;
  wire       _GEN_29644 = _GEN_1263 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_24;
  wire       _GEN_29645 = _GEN_1277 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_25;
  wire       _GEN_29646 = _GEN_1291 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_26;
  wire       _GEN_29647 = _GEN_1305 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_27;
  wire       _GEN_29648 = _GEN_1319 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_28;
  wire       _GEN_29649 = _GEN_1333 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_29;
  wire       _GEN_29650 = _GEN_1347 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_30;
  wire       _GEN_29651 = _GEN_1361 ? _rob_unsafe_2_rob_tail : rob_unsafe_2_31;
  wire       _GEN_32596 = _GEN_926 ? ~_GEN_929 & _GEN_29620 : ~_GEN_928 & _GEN_29620;
  wire       _GEN_32597 = _GEN_926 ? ~_GEN_943 & _GEN_29621 : ~_GEN_942 & _GEN_29621;
  wire       _GEN_32598 = _GEN_926 ? ~_GEN_957 & _GEN_29622 : ~_GEN_956 & _GEN_29622;
  wire       _GEN_32599 = _GEN_926 ? ~_GEN_971 & _GEN_29623 : ~_GEN_970 & _GEN_29623;
  wire       _GEN_32600 = _GEN_926 ? ~_GEN_985 & _GEN_29624 : ~_GEN_984 & _GEN_29624;
  wire       _GEN_32601 = _GEN_926 ? ~_GEN_999 & _GEN_29625 : ~_GEN_998 & _GEN_29625;
  wire       _GEN_32602 = _GEN_926 ? ~_GEN_1013 & _GEN_29626 : ~_GEN_1012 & _GEN_29626;
  wire       _GEN_32603 = _GEN_926 ? ~_GEN_1027 & _GEN_29627 : ~_GEN_1026 & _GEN_29627;
  wire       _GEN_32604 = _GEN_926 ? ~_GEN_1041 & _GEN_29628 : ~_GEN_1040 & _GEN_29628;
  wire       _GEN_32605 = _GEN_926 ? ~_GEN_1055 & _GEN_29629 : ~_GEN_1054 & _GEN_29629;
  wire       _GEN_32606 = _GEN_926 ? ~_GEN_1069 & _GEN_29630 : ~_GEN_1068 & _GEN_29630;
  wire       _GEN_32607 = _GEN_926 ? ~_GEN_1083 & _GEN_29631 : ~_GEN_1082 & _GEN_29631;
  wire       _GEN_32608 = _GEN_926 ? ~_GEN_1097 & _GEN_29632 : ~_GEN_1096 & _GEN_29632;
  wire       _GEN_32609 = _GEN_926 ? ~_GEN_1111 & _GEN_29633 : ~_GEN_1110 & _GEN_29633;
  wire       _GEN_32610 = _GEN_926 ? ~_GEN_1125 & _GEN_29634 : ~_GEN_1124 & _GEN_29634;
  wire       _GEN_32611 = _GEN_926 ? ~_GEN_1139 & _GEN_29635 : ~_GEN_1138 & _GEN_29635;
  wire       _GEN_32612 = _GEN_926 ? ~_GEN_1153 & _GEN_29636 : ~_GEN_1152 & _GEN_29636;
  wire       _GEN_32613 = _GEN_926 ? ~_GEN_1167 & _GEN_29637 : ~_GEN_1166 & _GEN_29637;
  wire       _GEN_32614 = _GEN_926 ? ~_GEN_1181 & _GEN_29638 : ~_GEN_1180 & _GEN_29638;
  wire       _GEN_32615 = _GEN_926 ? ~_GEN_1195 & _GEN_29639 : ~_GEN_1194 & _GEN_29639;
  wire       _GEN_32616 = _GEN_926 ? ~_GEN_1209 & _GEN_29640 : ~_GEN_1208 & _GEN_29640;
  wire       _GEN_32617 = _GEN_926 ? ~_GEN_1223 & _GEN_29641 : ~_GEN_1222 & _GEN_29641;
  wire       _GEN_32618 = _GEN_926 ? ~_GEN_1237 & _GEN_29642 : ~_GEN_1236 & _GEN_29642;
  wire       _GEN_32619 = _GEN_926 ? ~_GEN_1251 & _GEN_29643 : ~_GEN_1250 & _GEN_29643;
  wire       _GEN_32620 = _GEN_926 ? ~_GEN_1265 & _GEN_29644 : ~_GEN_1264 & _GEN_29644;
  wire       _GEN_32621 = _GEN_926 ? ~_GEN_1279 & _GEN_29645 : ~_GEN_1278 & _GEN_29645;
  wire       _GEN_32622 = _GEN_926 ? ~_GEN_1293 & _GEN_29646 : ~_GEN_1292 & _GEN_29646;
  wire       _GEN_32623 = _GEN_926 ? ~_GEN_1307 & _GEN_29647 : ~_GEN_1306 & _GEN_29647;
  wire       _GEN_32624 = _GEN_926 ? ~_GEN_1321 & _GEN_29648 : ~_GEN_1320 & _GEN_29648;
  wire       _GEN_32625 = _GEN_926 ? ~_GEN_1335 & _GEN_29649 : ~_GEN_1334 & _GEN_29649;
  wire       _GEN_32626 = _GEN_926 ? ~_GEN_1349 & _GEN_29650 : ~_GEN_1348 & _GEN_29650;
  wire       _GEN_32627 = _GEN_926 ? ~_GEN_1363 & _GEN_29651 : ~_GEN_1362 & _GEN_29651;
  wire       _GEN_32980 = _GEN_925 ? ~_GEN_931 & _GEN_32596 : ~_GEN_930 & _GEN_32596;
  wire       _GEN_32981 = _GEN_925 ? ~_GEN_945 & _GEN_32597 : ~_GEN_944 & _GEN_32597;
  wire       _GEN_32982 = _GEN_925 ? ~_GEN_959 & _GEN_32598 : ~_GEN_958 & _GEN_32598;
  wire       _GEN_32983 = _GEN_925 ? ~_GEN_973 & _GEN_32599 : ~_GEN_972 & _GEN_32599;
  wire       _GEN_32984 = _GEN_925 ? ~_GEN_987 & _GEN_32600 : ~_GEN_986 & _GEN_32600;
  wire       _GEN_32985 = _GEN_925 ? ~_GEN_1001 & _GEN_32601 : ~_GEN_1000 & _GEN_32601;
  wire       _GEN_32986 = _GEN_925 ? ~_GEN_1015 & _GEN_32602 : ~_GEN_1014 & _GEN_32602;
  wire       _GEN_32987 = _GEN_925 ? ~_GEN_1029 & _GEN_32603 : ~_GEN_1028 & _GEN_32603;
  wire       _GEN_32988 = _GEN_925 ? ~_GEN_1043 & _GEN_32604 : ~_GEN_1042 & _GEN_32604;
  wire       _GEN_32989 = _GEN_925 ? ~_GEN_1057 & _GEN_32605 : ~_GEN_1056 & _GEN_32605;
  wire       _GEN_32990 = _GEN_925 ? ~_GEN_1071 & _GEN_32606 : ~_GEN_1070 & _GEN_32606;
  wire       _GEN_32991 = _GEN_925 ? ~_GEN_1085 & _GEN_32607 : ~_GEN_1084 & _GEN_32607;
  wire       _GEN_32992 = _GEN_925 ? ~_GEN_1099 & _GEN_32608 : ~_GEN_1098 & _GEN_32608;
  wire       _GEN_32993 = _GEN_925 ? ~_GEN_1113 & _GEN_32609 : ~_GEN_1112 & _GEN_32609;
  wire       _GEN_32994 = _GEN_925 ? ~_GEN_1127 & _GEN_32610 : ~_GEN_1126 & _GEN_32610;
  wire       _GEN_32995 = _GEN_925 ? ~_GEN_1141 & _GEN_32611 : ~_GEN_1140 & _GEN_32611;
  wire       _GEN_32996 = _GEN_925 ? ~_GEN_1155 & _GEN_32612 : ~_GEN_1154 & _GEN_32612;
  wire       _GEN_32997 = _GEN_925 ? ~_GEN_1169 & _GEN_32613 : ~_GEN_1168 & _GEN_32613;
  wire       _GEN_32998 = _GEN_925 ? ~_GEN_1183 & _GEN_32614 : ~_GEN_1182 & _GEN_32614;
  wire       _GEN_32999 = _GEN_925 ? ~_GEN_1197 & _GEN_32615 : ~_GEN_1196 & _GEN_32615;
  wire       _GEN_33000 = _GEN_925 ? ~_GEN_1211 & _GEN_32616 : ~_GEN_1210 & _GEN_32616;
  wire       _GEN_33001 = _GEN_925 ? ~_GEN_1225 & _GEN_32617 : ~_GEN_1224 & _GEN_32617;
  wire       _GEN_33002 = _GEN_925 ? ~_GEN_1239 & _GEN_32618 : ~_GEN_1238 & _GEN_32618;
  wire       _GEN_33003 = _GEN_925 ? ~_GEN_1253 & _GEN_32619 : ~_GEN_1252 & _GEN_32619;
  wire       _GEN_33004 = _GEN_925 ? ~_GEN_1267 & _GEN_32620 : ~_GEN_1266 & _GEN_32620;
  wire       _GEN_33005 = _GEN_925 ? ~_GEN_1281 & _GEN_32621 : ~_GEN_1280 & _GEN_32621;
  wire       _GEN_33006 = _GEN_925 ? ~_GEN_1295 & _GEN_32622 : ~_GEN_1294 & _GEN_32622;
  wire       _GEN_33007 = _GEN_925 ? ~_GEN_1309 & _GEN_32623 : ~_GEN_1308 & _GEN_32623;
  wire       _GEN_33008 = _GEN_925 ? ~_GEN_1323 & _GEN_32624 : ~_GEN_1322 & _GEN_32624;
  wire       _GEN_33009 = _GEN_925 ? ~_GEN_1337 & _GEN_32625 : ~_GEN_1336 & _GEN_32625;
  wire       _GEN_33010 = _GEN_925 ? ~_GEN_1351 & _GEN_32626 : ~_GEN_1350 & _GEN_32626;
  wire       _GEN_33011 = _GEN_925 ? ~_GEN_1365 & _GEN_32627 : ~_GEN_1364 & _GEN_32627;
  wire       _GEN_33364 = _GEN_924 ? ~_GEN_933 & _GEN_32980 : ~_GEN_932 & _GEN_32980;
  wire       _GEN_33365 = _GEN_924 ? ~_GEN_947 & _GEN_32981 : ~_GEN_946 & _GEN_32981;
  wire       _GEN_33366 = _GEN_924 ? ~_GEN_961 & _GEN_32982 : ~_GEN_960 & _GEN_32982;
  wire       _GEN_33367 = _GEN_924 ? ~_GEN_975 & _GEN_32983 : ~_GEN_974 & _GEN_32983;
  wire       _GEN_33368 = _GEN_924 ? ~_GEN_989 & _GEN_32984 : ~_GEN_988 & _GEN_32984;
  wire       _GEN_33369 = _GEN_924 ? ~_GEN_1003 & _GEN_32985 : ~_GEN_1002 & _GEN_32985;
  wire       _GEN_33370 = _GEN_924 ? ~_GEN_1017 & _GEN_32986 : ~_GEN_1016 & _GEN_32986;
  wire       _GEN_33371 = _GEN_924 ? ~_GEN_1031 & _GEN_32987 : ~_GEN_1030 & _GEN_32987;
  wire       _GEN_33372 = _GEN_924 ? ~_GEN_1045 & _GEN_32988 : ~_GEN_1044 & _GEN_32988;
  wire       _GEN_33373 = _GEN_924 ? ~_GEN_1059 & _GEN_32989 : ~_GEN_1058 & _GEN_32989;
  wire       _GEN_33374 = _GEN_924 ? ~_GEN_1073 & _GEN_32990 : ~_GEN_1072 & _GEN_32990;
  wire       _GEN_33375 = _GEN_924 ? ~_GEN_1087 & _GEN_32991 : ~_GEN_1086 & _GEN_32991;
  wire       _GEN_33376 = _GEN_924 ? ~_GEN_1101 & _GEN_32992 : ~_GEN_1100 & _GEN_32992;
  wire       _GEN_33377 = _GEN_924 ? ~_GEN_1115 & _GEN_32993 : ~_GEN_1114 & _GEN_32993;
  wire       _GEN_33378 = _GEN_924 ? ~_GEN_1129 & _GEN_32994 : ~_GEN_1128 & _GEN_32994;
  wire       _GEN_33379 = _GEN_924 ? ~_GEN_1143 & _GEN_32995 : ~_GEN_1142 & _GEN_32995;
  wire       _GEN_33380 = _GEN_924 ? ~_GEN_1157 & _GEN_32996 : ~_GEN_1156 & _GEN_32996;
  wire       _GEN_33381 = _GEN_924 ? ~_GEN_1171 & _GEN_32997 : ~_GEN_1170 & _GEN_32997;
  wire       _GEN_33382 = _GEN_924 ? ~_GEN_1185 & _GEN_32998 : ~_GEN_1184 & _GEN_32998;
  wire       _GEN_33383 = _GEN_924 ? ~_GEN_1199 & _GEN_32999 : ~_GEN_1198 & _GEN_32999;
  wire       _GEN_33384 = _GEN_924 ? ~_GEN_1213 & _GEN_33000 : ~_GEN_1212 & _GEN_33000;
  wire       _GEN_33385 = _GEN_924 ? ~_GEN_1227 & _GEN_33001 : ~_GEN_1226 & _GEN_33001;
  wire       _GEN_33386 = _GEN_924 ? ~_GEN_1241 & _GEN_33002 : ~_GEN_1240 & _GEN_33002;
  wire       _GEN_33387 = _GEN_924 ? ~_GEN_1255 & _GEN_33003 : ~_GEN_1254 & _GEN_33003;
  wire       _GEN_33388 = _GEN_924 ? ~_GEN_1269 & _GEN_33004 : ~_GEN_1268 & _GEN_33004;
  wire       _GEN_33389 = _GEN_924 ? ~_GEN_1283 & _GEN_33005 : ~_GEN_1282 & _GEN_33005;
  wire       _GEN_33390 = _GEN_924 ? ~_GEN_1297 & _GEN_33006 : ~_GEN_1296 & _GEN_33006;
  wire       _GEN_33391 = _GEN_924 ? ~_GEN_1311 & _GEN_33007 : ~_GEN_1310 & _GEN_33007;
  wire       _GEN_33392 = _GEN_924 ? ~_GEN_1325 & _GEN_33008 : ~_GEN_1324 & _GEN_33008;
  wire       _GEN_33393 = _GEN_924 ? ~_GEN_1339 & _GEN_33009 : ~_GEN_1338 & _GEN_33009;
  wire       _GEN_33394 = _GEN_924 ? ~_GEN_1353 & _GEN_33010 : ~_GEN_1352 & _GEN_33010;
  wire       _GEN_33395 = _GEN_924 ? ~_GEN_1367 & _GEN_33011 : ~_GEN_1366 & _GEN_33011;
  wire       _GEN_33748 = _GEN_923 ? ~_GEN_935 & _GEN_33364 : ~_GEN_934 & _GEN_33364;
  wire       _GEN_33749 = _GEN_923 ? ~_GEN_949 & _GEN_33365 : ~_GEN_948 & _GEN_33365;
  wire       _GEN_33750 = _GEN_923 ? ~_GEN_963 & _GEN_33366 : ~_GEN_962 & _GEN_33366;
  wire       _GEN_33751 = _GEN_923 ? ~_GEN_977 & _GEN_33367 : ~_GEN_976 & _GEN_33367;
  wire       _GEN_33752 = _GEN_923 ? ~_GEN_991 & _GEN_33368 : ~_GEN_990 & _GEN_33368;
  wire       _GEN_33753 = _GEN_923 ? ~_GEN_1005 & _GEN_33369 : ~_GEN_1004 & _GEN_33369;
  wire       _GEN_33754 = _GEN_923 ? ~_GEN_1019 & _GEN_33370 : ~_GEN_1018 & _GEN_33370;
  wire       _GEN_33755 = _GEN_923 ? ~_GEN_1033 & _GEN_33371 : ~_GEN_1032 & _GEN_33371;
  wire       _GEN_33756 = _GEN_923 ? ~_GEN_1047 & _GEN_33372 : ~_GEN_1046 & _GEN_33372;
  wire       _GEN_33757 = _GEN_923 ? ~_GEN_1061 & _GEN_33373 : ~_GEN_1060 & _GEN_33373;
  wire       _GEN_33758 = _GEN_923 ? ~_GEN_1075 & _GEN_33374 : ~_GEN_1074 & _GEN_33374;
  wire       _GEN_33759 = _GEN_923 ? ~_GEN_1089 & _GEN_33375 : ~_GEN_1088 & _GEN_33375;
  wire       _GEN_33760 = _GEN_923 ? ~_GEN_1103 & _GEN_33376 : ~_GEN_1102 & _GEN_33376;
  wire       _GEN_33761 = _GEN_923 ? ~_GEN_1117 & _GEN_33377 : ~_GEN_1116 & _GEN_33377;
  wire       _GEN_33762 = _GEN_923 ? ~_GEN_1131 & _GEN_33378 : ~_GEN_1130 & _GEN_33378;
  wire       _GEN_33763 = _GEN_923 ? ~_GEN_1145 & _GEN_33379 : ~_GEN_1144 & _GEN_33379;
  wire       _GEN_33764 = _GEN_923 ? ~_GEN_1159 & _GEN_33380 : ~_GEN_1158 & _GEN_33380;
  wire       _GEN_33765 = _GEN_923 ? ~_GEN_1173 & _GEN_33381 : ~_GEN_1172 & _GEN_33381;
  wire       _GEN_33766 = _GEN_923 ? ~_GEN_1187 & _GEN_33382 : ~_GEN_1186 & _GEN_33382;
  wire       _GEN_33767 = _GEN_923 ? ~_GEN_1201 & _GEN_33383 : ~_GEN_1200 & _GEN_33383;
  wire       _GEN_33768 = _GEN_923 ? ~_GEN_1215 & _GEN_33384 : ~_GEN_1214 & _GEN_33384;
  wire       _GEN_33769 = _GEN_923 ? ~_GEN_1229 & _GEN_33385 : ~_GEN_1228 & _GEN_33385;
  wire       _GEN_33770 = _GEN_923 ? ~_GEN_1243 & _GEN_33386 : ~_GEN_1242 & _GEN_33386;
  wire       _GEN_33771 = _GEN_923 ? ~_GEN_1257 & _GEN_33387 : ~_GEN_1256 & _GEN_33387;
  wire       _GEN_33772 = _GEN_923 ? ~_GEN_1271 & _GEN_33388 : ~_GEN_1270 & _GEN_33388;
  wire       _GEN_33773 = _GEN_923 ? ~_GEN_1285 & _GEN_33389 : ~_GEN_1284 & _GEN_33389;
  wire       _GEN_33774 = _GEN_923 ? ~_GEN_1299 & _GEN_33390 : ~_GEN_1298 & _GEN_33390;
  wire       _GEN_33775 = _GEN_923 ? ~_GEN_1313 & _GEN_33391 : ~_GEN_1312 & _GEN_33391;
  wire       _GEN_33776 = _GEN_923 ? ~_GEN_1327 & _GEN_33392 : ~_GEN_1326 & _GEN_33392;
  wire       _GEN_33777 = _GEN_923 ? ~_GEN_1341 & _GEN_33393 : ~_GEN_1340 & _GEN_33393;
  wire       _GEN_33778 = _GEN_923 ? ~_GEN_1355 & _GEN_33394 : ~_GEN_1354 & _GEN_33394;
  wire       _GEN_33779 = _GEN_923 ? ~_GEN_1369 & _GEN_33395 : ~_GEN_1368 & _GEN_33395;
  wire       _GEN_34132 = _GEN_922 ? ~_GEN_937 & _GEN_33748 : ~_GEN_936 & _GEN_33748;
  wire       _GEN_34133 = _GEN_922 ? ~_GEN_951 & _GEN_33749 : ~_GEN_950 & _GEN_33749;
  wire       _GEN_34134 = _GEN_922 ? ~_GEN_965 & _GEN_33750 : ~_GEN_964 & _GEN_33750;
  wire       _GEN_34135 = _GEN_922 ? ~_GEN_979 & _GEN_33751 : ~_GEN_978 & _GEN_33751;
  wire       _GEN_34136 = _GEN_922 ? ~_GEN_993 & _GEN_33752 : ~_GEN_992 & _GEN_33752;
  wire       _GEN_34137 = _GEN_922 ? ~_GEN_1007 & _GEN_33753 : ~_GEN_1006 & _GEN_33753;
  wire       _GEN_34138 = _GEN_922 ? ~_GEN_1021 & _GEN_33754 : ~_GEN_1020 & _GEN_33754;
  wire       _GEN_34139 = _GEN_922 ? ~_GEN_1035 & _GEN_33755 : ~_GEN_1034 & _GEN_33755;
  wire       _GEN_34140 = _GEN_922 ? ~_GEN_1049 & _GEN_33756 : ~_GEN_1048 & _GEN_33756;
  wire       _GEN_34141 = _GEN_922 ? ~_GEN_1063 & _GEN_33757 : ~_GEN_1062 & _GEN_33757;
  wire       _GEN_34142 = _GEN_922 ? ~_GEN_1077 & _GEN_33758 : ~_GEN_1076 & _GEN_33758;
  wire       _GEN_34143 = _GEN_922 ? ~_GEN_1091 & _GEN_33759 : ~_GEN_1090 & _GEN_33759;
  wire       _GEN_34144 = _GEN_922 ? ~_GEN_1105 & _GEN_33760 : ~_GEN_1104 & _GEN_33760;
  wire       _GEN_34145 = _GEN_922 ? ~_GEN_1119 & _GEN_33761 : ~_GEN_1118 & _GEN_33761;
  wire       _GEN_34146 = _GEN_922 ? ~_GEN_1133 & _GEN_33762 : ~_GEN_1132 & _GEN_33762;
  wire       _GEN_34147 = _GEN_922 ? ~_GEN_1147 & _GEN_33763 : ~_GEN_1146 & _GEN_33763;
  wire       _GEN_34148 = _GEN_922 ? ~_GEN_1161 & _GEN_33764 : ~_GEN_1160 & _GEN_33764;
  wire       _GEN_34149 = _GEN_922 ? ~_GEN_1175 & _GEN_33765 : ~_GEN_1174 & _GEN_33765;
  wire       _GEN_34150 = _GEN_922 ? ~_GEN_1189 & _GEN_33766 : ~_GEN_1188 & _GEN_33766;
  wire       _GEN_34151 = _GEN_922 ? ~_GEN_1203 & _GEN_33767 : ~_GEN_1202 & _GEN_33767;
  wire       _GEN_34152 = _GEN_922 ? ~_GEN_1217 & _GEN_33768 : ~_GEN_1216 & _GEN_33768;
  wire       _GEN_34153 = _GEN_922 ? ~_GEN_1231 & _GEN_33769 : ~_GEN_1230 & _GEN_33769;
  wire       _GEN_34154 = _GEN_922 ? ~_GEN_1245 & _GEN_33770 : ~_GEN_1244 & _GEN_33770;
  wire       _GEN_34155 = _GEN_922 ? ~_GEN_1259 & _GEN_33771 : ~_GEN_1258 & _GEN_33771;
  wire       _GEN_34156 = _GEN_922 ? ~_GEN_1273 & _GEN_33772 : ~_GEN_1272 & _GEN_33772;
  wire       _GEN_34157 = _GEN_922 ? ~_GEN_1287 & _GEN_33773 : ~_GEN_1286 & _GEN_33773;
  wire       _GEN_34158 = _GEN_922 ? ~_GEN_1301 & _GEN_33774 : ~_GEN_1300 & _GEN_33774;
  wire       _GEN_34159 = _GEN_922 ? ~_GEN_1315 & _GEN_33775 : ~_GEN_1314 & _GEN_33775;
  wire       _GEN_34160 = _GEN_922 ? ~_GEN_1329 & _GEN_33776 : ~_GEN_1328 & _GEN_33776;
  wire       _GEN_34161 = _GEN_922 ? ~_GEN_1343 & _GEN_33777 : ~_GEN_1342 & _GEN_33777;
  wire       _GEN_34162 = _GEN_922 ? ~_GEN_1357 & _GEN_33778 : ~_GEN_1356 & _GEN_33778;
  wire       _GEN_34163 = _GEN_922 ? ~_GEN_1371 & _GEN_33779 : ~_GEN_1370 & _GEN_33779;
  wire       _rob_unsafe_3_rob_tail = io_enq_uops_3_uses_ldq | io_enq_uops_3_uses_stq & ~io_enq_uops_3_is_fence | io_enq_uops_3_is_br | io_enq_uops_3_is_jalr;
  wire       _GEN_42984 = _GEN_1386 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_0;
  wire       _GEN_42985 = _GEN_1400 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_1;
  wire       _GEN_42986 = _GEN_1414 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_2;
  wire       _GEN_42987 = _GEN_1428 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_3;
  wire       _GEN_42988 = _GEN_1442 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_4;
  wire       _GEN_42989 = _GEN_1456 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_5;
  wire       _GEN_42990 = _GEN_1470 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_6;
  wire       _GEN_42991 = _GEN_1484 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_7;
  wire       _GEN_42992 = _GEN_1498 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_8;
  wire       _GEN_42993 = _GEN_1512 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_9;
  wire       _GEN_42994 = _GEN_1526 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_10;
  wire       _GEN_42995 = _GEN_1540 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_11;
  wire       _GEN_42996 = _GEN_1554 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_12;
  wire       _GEN_42997 = _GEN_1568 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_13;
  wire       _GEN_42998 = _GEN_1582 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_14;
  wire       _GEN_42999 = _GEN_1596 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_15;
  wire       _GEN_43000 = _GEN_1610 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_16;
  wire       _GEN_43001 = _GEN_1624 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_17;
  wire       _GEN_43002 = _GEN_1638 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_18;
  wire       _GEN_43003 = _GEN_1652 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_19;
  wire       _GEN_43004 = _GEN_1666 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_20;
  wire       _GEN_43005 = _GEN_1680 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_21;
  wire       _GEN_43006 = _GEN_1694 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_22;
  wire       _GEN_43007 = _GEN_1708 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_23;
  wire       _GEN_43008 = _GEN_1722 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_24;
  wire       _GEN_43009 = _GEN_1736 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_25;
  wire       _GEN_43010 = _GEN_1750 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_26;
  wire       _GEN_43011 = _GEN_1764 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_27;
  wire       _GEN_43012 = _GEN_1778 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_28;
  wire       _GEN_43013 = _GEN_1792 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_29;
  wire       _GEN_43014 = _GEN_1806 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_30;
  wire       _GEN_43015 = _GEN_1820 ? _rob_unsafe_3_rob_tail : rob_unsafe_3_31;
  wire       _GEN_45960 = _GEN_1385 ? ~_GEN_1388 & _GEN_42984 : ~_GEN_1387 & _GEN_42984;
  wire       _GEN_45961 = _GEN_1385 ? ~_GEN_1402 & _GEN_42985 : ~_GEN_1401 & _GEN_42985;
  wire       _GEN_45962 = _GEN_1385 ? ~_GEN_1416 & _GEN_42986 : ~_GEN_1415 & _GEN_42986;
  wire       _GEN_45963 = _GEN_1385 ? ~_GEN_1430 & _GEN_42987 : ~_GEN_1429 & _GEN_42987;
  wire       _GEN_45964 = _GEN_1385 ? ~_GEN_1444 & _GEN_42988 : ~_GEN_1443 & _GEN_42988;
  wire       _GEN_45965 = _GEN_1385 ? ~_GEN_1458 & _GEN_42989 : ~_GEN_1457 & _GEN_42989;
  wire       _GEN_45966 = _GEN_1385 ? ~_GEN_1472 & _GEN_42990 : ~_GEN_1471 & _GEN_42990;
  wire       _GEN_45967 = _GEN_1385 ? ~_GEN_1486 & _GEN_42991 : ~_GEN_1485 & _GEN_42991;
  wire       _GEN_45968 = _GEN_1385 ? ~_GEN_1500 & _GEN_42992 : ~_GEN_1499 & _GEN_42992;
  wire       _GEN_45969 = _GEN_1385 ? ~_GEN_1514 & _GEN_42993 : ~_GEN_1513 & _GEN_42993;
  wire       _GEN_45970 = _GEN_1385 ? ~_GEN_1528 & _GEN_42994 : ~_GEN_1527 & _GEN_42994;
  wire       _GEN_45971 = _GEN_1385 ? ~_GEN_1542 & _GEN_42995 : ~_GEN_1541 & _GEN_42995;
  wire       _GEN_45972 = _GEN_1385 ? ~_GEN_1556 & _GEN_42996 : ~_GEN_1555 & _GEN_42996;
  wire       _GEN_45973 = _GEN_1385 ? ~_GEN_1570 & _GEN_42997 : ~_GEN_1569 & _GEN_42997;
  wire       _GEN_45974 = _GEN_1385 ? ~_GEN_1584 & _GEN_42998 : ~_GEN_1583 & _GEN_42998;
  wire       _GEN_45975 = _GEN_1385 ? ~_GEN_1598 & _GEN_42999 : ~_GEN_1597 & _GEN_42999;
  wire       _GEN_45976 = _GEN_1385 ? ~_GEN_1612 & _GEN_43000 : ~_GEN_1611 & _GEN_43000;
  wire       _GEN_45977 = _GEN_1385 ? ~_GEN_1626 & _GEN_43001 : ~_GEN_1625 & _GEN_43001;
  wire       _GEN_45978 = _GEN_1385 ? ~_GEN_1640 & _GEN_43002 : ~_GEN_1639 & _GEN_43002;
  wire       _GEN_45979 = _GEN_1385 ? ~_GEN_1654 & _GEN_43003 : ~_GEN_1653 & _GEN_43003;
  wire       _GEN_45980 = _GEN_1385 ? ~_GEN_1668 & _GEN_43004 : ~_GEN_1667 & _GEN_43004;
  wire       _GEN_45981 = _GEN_1385 ? ~_GEN_1682 & _GEN_43005 : ~_GEN_1681 & _GEN_43005;
  wire       _GEN_45982 = _GEN_1385 ? ~_GEN_1696 & _GEN_43006 : ~_GEN_1695 & _GEN_43006;
  wire       _GEN_45983 = _GEN_1385 ? ~_GEN_1710 & _GEN_43007 : ~_GEN_1709 & _GEN_43007;
  wire       _GEN_45984 = _GEN_1385 ? ~_GEN_1724 & _GEN_43008 : ~_GEN_1723 & _GEN_43008;
  wire       _GEN_45985 = _GEN_1385 ? ~_GEN_1738 & _GEN_43009 : ~_GEN_1737 & _GEN_43009;
  wire       _GEN_45986 = _GEN_1385 ? ~_GEN_1752 & _GEN_43010 : ~_GEN_1751 & _GEN_43010;
  wire       _GEN_45987 = _GEN_1385 ? ~_GEN_1766 & _GEN_43011 : ~_GEN_1765 & _GEN_43011;
  wire       _GEN_45988 = _GEN_1385 ? ~_GEN_1780 & _GEN_43012 : ~_GEN_1779 & _GEN_43012;
  wire       _GEN_45989 = _GEN_1385 ? ~_GEN_1794 & _GEN_43013 : ~_GEN_1793 & _GEN_43013;
  wire       _GEN_45990 = _GEN_1385 ? ~_GEN_1808 & _GEN_43014 : ~_GEN_1807 & _GEN_43014;
  wire       _GEN_45991 = _GEN_1385 ? ~_GEN_1822 & _GEN_43015 : ~_GEN_1821 & _GEN_43015;
  wire       _GEN_46344 = _GEN_1384 ? ~_GEN_1390 & _GEN_45960 : ~_GEN_1389 & _GEN_45960;
  wire       _GEN_46345 = _GEN_1384 ? ~_GEN_1404 & _GEN_45961 : ~_GEN_1403 & _GEN_45961;
  wire       _GEN_46346 = _GEN_1384 ? ~_GEN_1418 & _GEN_45962 : ~_GEN_1417 & _GEN_45962;
  wire       _GEN_46347 = _GEN_1384 ? ~_GEN_1432 & _GEN_45963 : ~_GEN_1431 & _GEN_45963;
  wire       _GEN_46348 = _GEN_1384 ? ~_GEN_1446 & _GEN_45964 : ~_GEN_1445 & _GEN_45964;
  wire       _GEN_46349 = _GEN_1384 ? ~_GEN_1460 & _GEN_45965 : ~_GEN_1459 & _GEN_45965;
  wire       _GEN_46350 = _GEN_1384 ? ~_GEN_1474 & _GEN_45966 : ~_GEN_1473 & _GEN_45966;
  wire       _GEN_46351 = _GEN_1384 ? ~_GEN_1488 & _GEN_45967 : ~_GEN_1487 & _GEN_45967;
  wire       _GEN_46352 = _GEN_1384 ? ~_GEN_1502 & _GEN_45968 : ~_GEN_1501 & _GEN_45968;
  wire       _GEN_46353 = _GEN_1384 ? ~_GEN_1516 & _GEN_45969 : ~_GEN_1515 & _GEN_45969;
  wire       _GEN_46354 = _GEN_1384 ? ~_GEN_1530 & _GEN_45970 : ~_GEN_1529 & _GEN_45970;
  wire       _GEN_46355 = _GEN_1384 ? ~_GEN_1544 & _GEN_45971 : ~_GEN_1543 & _GEN_45971;
  wire       _GEN_46356 = _GEN_1384 ? ~_GEN_1558 & _GEN_45972 : ~_GEN_1557 & _GEN_45972;
  wire       _GEN_46357 = _GEN_1384 ? ~_GEN_1572 & _GEN_45973 : ~_GEN_1571 & _GEN_45973;
  wire       _GEN_46358 = _GEN_1384 ? ~_GEN_1586 & _GEN_45974 : ~_GEN_1585 & _GEN_45974;
  wire       _GEN_46359 = _GEN_1384 ? ~_GEN_1600 & _GEN_45975 : ~_GEN_1599 & _GEN_45975;
  wire       _GEN_46360 = _GEN_1384 ? ~_GEN_1614 & _GEN_45976 : ~_GEN_1613 & _GEN_45976;
  wire       _GEN_46361 = _GEN_1384 ? ~_GEN_1628 & _GEN_45977 : ~_GEN_1627 & _GEN_45977;
  wire       _GEN_46362 = _GEN_1384 ? ~_GEN_1642 & _GEN_45978 : ~_GEN_1641 & _GEN_45978;
  wire       _GEN_46363 = _GEN_1384 ? ~_GEN_1656 & _GEN_45979 : ~_GEN_1655 & _GEN_45979;
  wire       _GEN_46364 = _GEN_1384 ? ~_GEN_1670 & _GEN_45980 : ~_GEN_1669 & _GEN_45980;
  wire       _GEN_46365 = _GEN_1384 ? ~_GEN_1684 & _GEN_45981 : ~_GEN_1683 & _GEN_45981;
  wire       _GEN_46366 = _GEN_1384 ? ~_GEN_1698 & _GEN_45982 : ~_GEN_1697 & _GEN_45982;
  wire       _GEN_46367 = _GEN_1384 ? ~_GEN_1712 & _GEN_45983 : ~_GEN_1711 & _GEN_45983;
  wire       _GEN_46368 = _GEN_1384 ? ~_GEN_1726 & _GEN_45984 : ~_GEN_1725 & _GEN_45984;
  wire       _GEN_46369 = _GEN_1384 ? ~_GEN_1740 & _GEN_45985 : ~_GEN_1739 & _GEN_45985;
  wire       _GEN_46370 = _GEN_1384 ? ~_GEN_1754 & _GEN_45986 : ~_GEN_1753 & _GEN_45986;
  wire       _GEN_46371 = _GEN_1384 ? ~_GEN_1768 & _GEN_45987 : ~_GEN_1767 & _GEN_45987;
  wire       _GEN_46372 = _GEN_1384 ? ~_GEN_1782 & _GEN_45988 : ~_GEN_1781 & _GEN_45988;
  wire       _GEN_46373 = _GEN_1384 ? ~_GEN_1796 & _GEN_45989 : ~_GEN_1795 & _GEN_45989;
  wire       _GEN_46374 = _GEN_1384 ? ~_GEN_1810 & _GEN_45990 : ~_GEN_1809 & _GEN_45990;
  wire       _GEN_46375 = _GEN_1384 ? ~_GEN_1824 & _GEN_45991 : ~_GEN_1823 & _GEN_45991;
  wire       _GEN_46728 = _GEN_1383 ? ~_GEN_1392 & _GEN_46344 : ~_GEN_1391 & _GEN_46344;
  wire       _GEN_46729 = _GEN_1383 ? ~_GEN_1406 & _GEN_46345 : ~_GEN_1405 & _GEN_46345;
  wire       _GEN_46730 = _GEN_1383 ? ~_GEN_1420 & _GEN_46346 : ~_GEN_1419 & _GEN_46346;
  wire       _GEN_46731 = _GEN_1383 ? ~_GEN_1434 & _GEN_46347 : ~_GEN_1433 & _GEN_46347;
  wire       _GEN_46732 = _GEN_1383 ? ~_GEN_1448 & _GEN_46348 : ~_GEN_1447 & _GEN_46348;
  wire       _GEN_46733 = _GEN_1383 ? ~_GEN_1462 & _GEN_46349 : ~_GEN_1461 & _GEN_46349;
  wire       _GEN_46734 = _GEN_1383 ? ~_GEN_1476 & _GEN_46350 : ~_GEN_1475 & _GEN_46350;
  wire       _GEN_46735 = _GEN_1383 ? ~_GEN_1490 & _GEN_46351 : ~_GEN_1489 & _GEN_46351;
  wire       _GEN_46736 = _GEN_1383 ? ~_GEN_1504 & _GEN_46352 : ~_GEN_1503 & _GEN_46352;
  wire       _GEN_46737 = _GEN_1383 ? ~_GEN_1518 & _GEN_46353 : ~_GEN_1517 & _GEN_46353;
  wire       _GEN_46738 = _GEN_1383 ? ~_GEN_1532 & _GEN_46354 : ~_GEN_1531 & _GEN_46354;
  wire       _GEN_46739 = _GEN_1383 ? ~_GEN_1546 & _GEN_46355 : ~_GEN_1545 & _GEN_46355;
  wire       _GEN_46740 = _GEN_1383 ? ~_GEN_1560 & _GEN_46356 : ~_GEN_1559 & _GEN_46356;
  wire       _GEN_46741 = _GEN_1383 ? ~_GEN_1574 & _GEN_46357 : ~_GEN_1573 & _GEN_46357;
  wire       _GEN_46742 = _GEN_1383 ? ~_GEN_1588 & _GEN_46358 : ~_GEN_1587 & _GEN_46358;
  wire       _GEN_46743 = _GEN_1383 ? ~_GEN_1602 & _GEN_46359 : ~_GEN_1601 & _GEN_46359;
  wire       _GEN_46744 = _GEN_1383 ? ~_GEN_1616 & _GEN_46360 : ~_GEN_1615 & _GEN_46360;
  wire       _GEN_46745 = _GEN_1383 ? ~_GEN_1630 & _GEN_46361 : ~_GEN_1629 & _GEN_46361;
  wire       _GEN_46746 = _GEN_1383 ? ~_GEN_1644 & _GEN_46362 : ~_GEN_1643 & _GEN_46362;
  wire       _GEN_46747 = _GEN_1383 ? ~_GEN_1658 & _GEN_46363 : ~_GEN_1657 & _GEN_46363;
  wire       _GEN_46748 = _GEN_1383 ? ~_GEN_1672 & _GEN_46364 : ~_GEN_1671 & _GEN_46364;
  wire       _GEN_46749 = _GEN_1383 ? ~_GEN_1686 & _GEN_46365 : ~_GEN_1685 & _GEN_46365;
  wire       _GEN_46750 = _GEN_1383 ? ~_GEN_1700 & _GEN_46366 : ~_GEN_1699 & _GEN_46366;
  wire       _GEN_46751 = _GEN_1383 ? ~_GEN_1714 & _GEN_46367 : ~_GEN_1713 & _GEN_46367;
  wire       _GEN_46752 = _GEN_1383 ? ~_GEN_1728 & _GEN_46368 : ~_GEN_1727 & _GEN_46368;
  wire       _GEN_46753 = _GEN_1383 ? ~_GEN_1742 & _GEN_46369 : ~_GEN_1741 & _GEN_46369;
  wire       _GEN_46754 = _GEN_1383 ? ~_GEN_1756 & _GEN_46370 : ~_GEN_1755 & _GEN_46370;
  wire       _GEN_46755 = _GEN_1383 ? ~_GEN_1770 & _GEN_46371 : ~_GEN_1769 & _GEN_46371;
  wire       _GEN_46756 = _GEN_1383 ? ~_GEN_1784 & _GEN_46372 : ~_GEN_1783 & _GEN_46372;
  wire       _GEN_46757 = _GEN_1383 ? ~_GEN_1798 & _GEN_46373 : ~_GEN_1797 & _GEN_46373;
  wire       _GEN_46758 = _GEN_1383 ? ~_GEN_1812 & _GEN_46374 : ~_GEN_1811 & _GEN_46374;
  wire       _GEN_46759 = _GEN_1383 ? ~_GEN_1826 & _GEN_46375 : ~_GEN_1825 & _GEN_46375;
  wire       _GEN_47112 = _GEN_1382 ? ~_GEN_1394 & _GEN_46728 : ~_GEN_1393 & _GEN_46728;
  wire       _GEN_47113 = _GEN_1382 ? ~_GEN_1408 & _GEN_46729 : ~_GEN_1407 & _GEN_46729;
  wire       _GEN_47114 = _GEN_1382 ? ~_GEN_1422 & _GEN_46730 : ~_GEN_1421 & _GEN_46730;
  wire       _GEN_47115 = _GEN_1382 ? ~_GEN_1436 & _GEN_46731 : ~_GEN_1435 & _GEN_46731;
  wire       _GEN_47116 = _GEN_1382 ? ~_GEN_1450 & _GEN_46732 : ~_GEN_1449 & _GEN_46732;
  wire       _GEN_47117 = _GEN_1382 ? ~_GEN_1464 & _GEN_46733 : ~_GEN_1463 & _GEN_46733;
  wire       _GEN_47118 = _GEN_1382 ? ~_GEN_1478 & _GEN_46734 : ~_GEN_1477 & _GEN_46734;
  wire       _GEN_47119 = _GEN_1382 ? ~_GEN_1492 & _GEN_46735 : ~_GEN_1491 & _GEN_46735;
  wire       _GEN_47120 = _GEN_1382 ? ~_GEN_1506 & _GEN_46736 : ~_GEN_1505 & _GEN_46736;
  wire       _GEN_47121 = _GEN_1382 ? ~_GEN_1520 & _GEN_46737 : ~_GEN_1519 & _GEN_46737;
  wire       _GEN_47122 = _GEN_1382 ? ~_GEN_1534 & _GEN_46738 : ~_GEN_1533 & _GEN_46738;
  wire       _GEN_47123 = _GEN_1382 ? ~_GEN_1548 & _GEN_46739 : ~_GEN_1547 & _GEN_46739;
  wire       _GEN_47124 = _GEN_1382 ? ~_GEN_1562 & _GEN_46740 : ~_GEN_1561 & _GEN_46740;
  wire       _GEN_47125 = _GEN_1382 ? ~_GEN_1576 & _GEN_46741 : ~_GEN_1575 & _GEN_46741;
  wire       _GEN_47126 = _GEN_1382 ? ~_GEN_1590 & _GEN_46742 : ~_GEN_1589 & _GEN_46742;
  wire       _GEN_47127 = _GEN_1382 ? ~_GEN_1604 & _GEN_46743 : ~_GEN_1603 & _GEN_46743;
  wire       _GEN_47128 = _GEN_1382 ? ~_GEN_1618 & _GEN_46744 : ~_GEN_1617 & _GEN_46744;
  wire       _GEN_47129 = _GEN_1382 ? ~_GEN_1632 & _GEN_46745 : ~_GEN_1631 & _GEN_46745;
  wire       _GEN_47130 = _GEN_1382 ? ~_GEN_1646 & _GEN_46746 : ~_GEN_1645 & _GEN_46746;
  wire       _GEN_47131 = _GEN_1382 ? ~_GEN_1660 & _GEN_46747 : ~_GEN_1659 & _GEN_46747;
  wire       _GEN_47132 = _GEN_1382 ? ~_GEN_1674 & _GEN_46748 : ~_GEN_1673 & _GEN_46748;
  wire       _GEN_47133 = _GEN_1382 ? ~_GEN_1688 & _GEN_46749 : ~_GEN_1687 & _GEN_46749;
  wire       _GEN_47134 = _GEN_1382 ? ~_GEN_1702 & _GEN_46750 : ~_GEN_1701 & _GEN_46750;
  wire       _GEN_47135 = _GEN_1382 ? ~_GEN_1716 & _GEN_46751 : ~_GEN_1715 & _GEN_46751;
  wire       _GEN_47136 = _GEN_1382 ? ~_GEN_1730 & _GEN_46752 : ~_GEN_1729 & _GEN_46752;
  wire       _GEN_47137 = _GEN_1382 ? ~_GEN_1744 & _GEN_46753 : ~_GEN_1743 & _GEN_46753;
  wire       _GEN_47138 = _GEN_1382 ? ~_GEN_1758 & _GEN_46754 : ~_GEN_1757 & _GEN_46754;
  wire       _GEN_47139 = _GEN_1382 ? ~_GEN_1772 & _GEN_46755 : ~_GEN_1771 & _GEN_46755;
  wire       _GEN_47140 = _GEN_1382 ? ~_GEN_1786 & _GEN_46756 : ~_GEN_1785 & _GEN_46756;
  wire       _GEN_47141 = _GEN_1382 ? ~_GEN_1800 & _GEN_46757 : ~_GEN_1799 & _GEN_46757;
  wire       _GEN_47142 = _GEN_1382 ? ~_GEN_1814 & _GEN_46758 : ~_GEN_1813 & _GEN_46758;
  wire       _GEN_47143 = _GEN_1382 ? ~_GEN_1828 & _GEN_46759 : ~_GEN_1827 & _GEN_46759;
  wire       _GEN_47496 = _GEN_1381 ? ~_GEN_1396 & _GEN_47112 : ~_GEN_1395 & _GEN_47112;
  wire       _GEN_47497 = _GEN_1381 ? ~_GEN_1410 & _GEN_47113 : ~_GEN_1409 & _GEN_47113;
  wire       _GEN_47498 = _GEN_1381 ? ~_GEN_1424 & _GEN_47114 : ~_GEN_1423 & _GEN_47114;
  wire       _GEN_47499 = _GEN_1381 ? ~_GEN_1438 & _GEN_47115 : ~_GEN_1437 & _GEN_47115;
  wire       _GEN_47500 = _GEN_1381 ? ~_GEN_1452 & _GEN_47116 : ~_GEN_1451 & _GEN_47116;
  wire       _GEN_47501 = _GEN_1381 ? ~_GEN_1466 & _GEN_47117 : ~_GEN_1465 & _GEN_47117;
  wire       _GEN_47502 = _GEN_1381 ? ~_GEN_1480 & _GEN_47118 : ~_GEN_1479 & _GEN_47118;
  wire       _GEN_47503 = _GEN_1381 ? ~_GEN_1494 & _GEN_47119 : ~_GEN_1493 & _GEN_47119;
  wire       _GEN_47504 = _GEN_1381 ? ~_GEN_1508 & _GEN_47120 : ~_GEN_1507 & _GEN_47120;
  wire       _GEN_47505 = _GEN_1381 ? ~_GEN_1522 & _GEN_47121 : ~_GEN_1521 & _GEN_47121;
  wire       _GEN_47506 = _GEN_1381 ? ~_GEN_1536 & _GEN_47122 : ~_GEN_1535 & _GEN_47122;
  wire       _GEN_47507 = _GEN_1381 ? ~_GEN_1550 & _GEN_47123 : ~_GEN_1549 & _GEN_47123;
  wire       _GEN_47508 = _GEN_1381 ? ~_GEN_1564 & _GEN_47124 : ~_GEN_1563 & _GEN_47124;
  wire       _GEN_47509 = _GEN_1381 ? ~_GEN_1578 & _GEN_47125 : ~_GEN_1577 & _GEN_47125;
  wire       _GEN_47510 = _GEN_1381 ? ~_GEN_1592 & _GEN_47126 : ~_GEN_1591 & _GEN_47126;
  wire       _GEN_47511 = _GEN_1381 ? ~_GEN_1606 & _GEN_47127 : ~_GEN_1605 & _GEN_47127;
  wire       _GEN_47512 = _GEN_1381 ? ~_GEN_1620 & _GEN_47128 : ~_GEN_1619 & _GEN_47128;
  wire       _GEN_47513 = _GEN_1381 ? ~_GEN_1634 & _GEN_47129 : ~_GEN_1633 & _GEN_47129;
  wire       _GEN_47514 = _GEN_1381 ? ~_GEN_1648 & _GEN_47130 : ~_GEN_1647 & _GEN_47130;
  wire       _GEN_47515 = _GEN_1381 ? ~_GEN_1662 & _GEN_47131 : ~_GEN_1661 & _GEN_47131;
  wire       _GEN_47516 = _GEN_1381 ? ~_GEN_1676 & _GEN_47132 : ~_GEN_1675 & _GEN_47132;
  wire       _GEN_47517 = _GEN_1381 ? ~_GEN_1690 & _GEN_47133 : ~_GEN_1689 & _GEN_47133;
  wire       _GEN_47518 = _GEN_1381 ? ~_GEN_1704 & _GEN_47134 : ~_GEN_1703 & _GEN_47134;
  wire       _GEN_47519 = _GEN_1381 ? ~_GEN_1718 & _GEN_47135 : ~_GEN_1717 & _GEN_47135;
  wire       _GEN_47520 = _GEN_1381 ? ~_GEN_1732 & _GEN_47136 : ~_GEN_1731 & _GEN_47136;
  wire       _GEN_47521 = _GEN_1381 ? ~_GEN_1746 & _GEN_47137 : ~_GEN_1745 & _GEN_47137;
  wire       _GEN_47522 = _GEN_1381 ? ~_GEN_1760 & _GEN_47138 : ~_GEN_1759 & _GEN_47138;
  wire       _GEN_47523 = _GEN_1381 ? ~_GEN_1774 & _GEN_47139 : ~_GEN_1773 & _GEN_47139;
  wire       _GEN_47524 = _GEN_1381 ? ~_GEN_1788 & _GEN_47140 : ~_GEN_1787 & _GEN_47140;
  wire       _GEN_47525 = _GEN_1381 ? ~_GEN_1802 & _GEN_47141 : ~_GEN_1801 & _GEN_47141;
  wire       _GEN_47526 = _GEN_1381 ? ~_GEN_1816 & _GEN_47142 : ~_GEN_1815 & _GEN_47142;
  wire       _GEN_47527 = _GEN_1381 ? ~_GEN_1830 & _GEN_47143 : ~_GEN_1829 & _GEN_47143;
  always @(posedge clock) begin
    if (_GEN_1993) begin
      assert__assert: assert(~casez_tmp);
      assert__assert_1: assert(_GEN_1852);
    end
    if (_GEN_1994) begin
      assert__assert_2: assert(casez_tmp_0);
      assert__assert_3: assert(casez_tmp_1);
    end
    if (_GEN_1995) begin
      assert__assert_4: assert(casez_tmp_2);
      assert__assert_5: assert(casez_tmp_3);
    end
    if (_GEN_1996) begin
      assert__assert_6: assert(casez_tmp_4);
      assert__assert_7: assert(casez_tmp_5);
    end
    if (_GEN_1997)
      assert__assert_8: assert(casez_tmp_6);
    if (~reset) begin
      assert__assert_9: assert(~_GEN_1854);
      assert__assert_10: assert(~_GEN_1855);
      assert__assert_11: assert(~_GEN_1856);
      assert__assert_12: assert(~_GEN_1857);
      assert__assert_13: assert(~_GEN_1858);
      assert__assert_14: assert(~_GEN_1859);
      assert__assert_15: assert(~_GEN_1860);
      assert__assert_16: assert(~_GEN_1861);
      assert__assert_17: assert(~_GEN_1862);
      assert__assert_18: assert(~_GEN_1863);
      assert__assert_19: assert(~_GEN_1864);
      assert__assert_20: assert(~_GEN_1865);
      assert__assert_21: assert(~_GEN_1866);
      assert__assert_22: assert(~_GEN_1867);
      assert__assert_23: assert(~_GEN_1868);
      assert__assert_24: assert(~_GEN_1869);
      assert__assert_25: assert(~_GEN_1870);
      assert__assert_26: assert(~_GEN_1871);
      assert__assert_27: assert(~_GEN_1872);
      assert__assert_28: assert(~_GEN_1873);
      assert__assert_29: assert(~_GEN_1874);
      assert__assert_30: assert(~_GEN_1875);
      assert__assert_31: assert(~_GEN_1876);
      assert__assert_32: assert(~_GEN_1877);
      assert__assert_33: assert(~_GEN_1878);
      assert__assert_34: assert(~_GEN_1879);
      assert__assert_35: assert(~_GEN_1880);
      assert__assert_36: assert(~_GEN_1881);
      assert__assert_37: assert(~_GEN_1882);
      assert__assert_38: assert(~_GEN_1883);
      assert__assert_39: assert(~_GEN_1884);
    end
    if (_GEN_1998) begin
      assert__assert_40: assert(~casez_tmp_50);
      assert__assert_41: assert(_GEN_1885);
    end
    if (_GEN_1999) begin
      assert__assert_42: assert(casez_tmp_51);
      assert__assert_43: assert(casez_tmp_52);
    end
    if (_GEN_2000) begin
      assert__assert_44: assert(casez_tmp_53);
      assert__assert_45: assert(casez_tmp_54);
    end
    if (_GEN_2001) begin
      assert__assert_46: assert(casez_tmp_55);
      assert__assert_47: assert(casez_tmp_56);
    end
    if (_GEN_2002)
      assert__assert_48: assert(casez_tmp_57);
    if (~reset) begin
      assert__assert_49: assert(~_GEN_1854);
      assert__assert_50: assert(~_GEN_1886);
      assert__assert_51: assert(~_GEN_1887);
      assert__assert_52: assert(~_GEN_1888);
      assert__assert_53: assert(~_GEN_1889);
      assert__assert_54: assert(~_GEN_1890);
      assert__assert_55: assert(~_GEN_1891);
      assert__assert_56: assert(~_GEN_1892);
      assert__assert_57: assert(~_GEN_1893);
      assert__assert_58: assert(~_GEN_1894);
      assert__assert_59: assert(~_GEN_1895);
      assert__assert_60: assert(~_GEN_1896);
      assert__assert_61: assert(~_GEN_1897);
      assert__assert_62: assert(~_GEN_1898);
      assert__assert_63: assert(~_GEN_1899);
      assert__assert_64: assert(~_GEN_1900);
      assert__assert_65: assert(~_GEN_1901);
      assert__assert_66: assert(~_GEN_1902);
      assert__assert_67: assert(~_GEN_1903);
      assert__assert_68: assert(~_GEN_1904);
      assert__assert_69: assert(~_GEN_1905);
      assert__assert_70: assert(~_GEN_1906);
      assert__assert_71: assert(~_GEN_1907);
      assert__assert_72: assert(~_GEN_1908);
      assert__assert_73: assert(~_GEN_1909);
      assert__assert_74: assert(~_GEN_1910);
      assert__assert_75: assert(~_GEN_1911);
      assert__assert_76: assert(~_GEN_1912);
      assert__assert_77: assert(~_GEN_1913);
      assert__assert_78: assert(~_GEN_1914);
      assert__assert_79: assert(~_GEN_1915);
    end
    if (_GEN_2003) begin
      assert__assert_80: assert(~casez_tmp_101);
      assert__assert_81: assert(_GEN_1916);
    end
    if (_GEN_2004) begin
      assert__assert_82: assert(casez_tmp_102);
      assert__assert_83: assert(casez_tmp_103);
    end
    if (_GEN_2005) begin
      assert__assert_84: assert(casez_tmp_104);
      assert__assert_85: assert(casez_tmp_105);
    end
    if (_GEN_2006) begin
      assert__assert_86: assert(casez_tmp_106);
      assert__assert_87: assert(casez_tmp_107);
    end
    if (_GEN_2007)
      assert__assert_88: assert(casez_tmp_108);
    if (~reset) begin
      assert__assert_89: assert(~_GEN_1854);
      assert__assert_90: assert(~_GEN_1917);
      assert__assert_91: assert(~_GEN_1918);
      assert__assert_92: assert(~_GEN_1919);
      assert__assert_93: assert(~_GEN_1920);
      assert__assert_94: assert(~_GEN_1921);
      assert__assert_95: assert(~_GEN_1922);
      assert__assert_96: assert(~_GEN_1923);
      assert__assert_97: assert(~_GEN_1924);
      assert__assert_98: assert(~_GEN_1925);
      assert__assert_99: assert(~_GEN_1926);
      assert__assert_100: assert(~_GEN_1927);
      assert__assert_101: assert(~_GEN_1928);
      assert__assert_102: assert(~_GEN_1929);
      assert__assert_103: assert(~_GEN_1930);
      assert__assert_104: assert(~_GEN_1931);
      assert__assert_105: assert(~_GEN_1932);
      assert__assert_106: assert(~_GEN_1933);
      assert__assert_107: assert(~_GEN_1934);
      assert__assert_108: assert(~_GEN_1935);
      assert__assert_109: assert(~_GEN_1936);
      assert__assert_110: assert(~_GEN_1937);
      assert__assert_111: assert(~_GEN_1938);
      assert__assert_112: assert(~_GEN_1939);
      assert__assert_113: assert(~_GEN_1940);
      assert__assert_114: assert(~_GEN_1941);
      assert__assert_115: assert(~_GEN_1942);
      assert__assert_116: assert(~_GEN_1943);
      assert__assert_117: assert(~_GEN_1944);
      assert__assert_118: assert(~_GEN_1945);
      assert__assert_119: assert(~_GEN_1946);
    end
    if (_GEN_2008) begin
      assert__assert_120: assert(~casez_tmp_152);
      assert__assert_121: assert(_GEN_1947);
    end
    if (_GEN_2009) begin
      assert__assert_122: assert(casez_tmp_153);
      assert__assert_123: assert(casez_tmp_154);
    end
    if (_GEN_2010) begin
      assert__assert_124: assert(casez_tmp_155);
      assert__assert_125: assert(casez_tmp_156);
    end
    if (_GEN_2011) begin
      assert__assert_126: assert(casez_tmp_157);
      assert__assert_127: assert(casez_tmp_158);
    end
    if (_GEN_2012)
      assert__assert_128: assert(casez_tmp_159);
    if (~reset) begin
      assert__assert_129: assert(~_GEN_1854);
      assert__assert_130: assert(~_GEN_1948);
      assert__assert_131: assert(~_GEN_1949);
      assert__assert_132: assert(~_GEN_1950);
      assert__assert_133: assert(~_GEN_1951);
      assert__assert_134: assert(~_GEN_1952);
      assert__assert_135: assert(~_GEN_1953);
      assert__assert_136: assert(~_GEN_1954);
      assert__assert_137: assert(~_GEN_1955);
      assert__assert_138: assert(~_GEN_1956);
      assert__assert_139: assert(~_GEN_1957);
      assert__assert_140: assert(~_GEN_1958);
      assert__assert_141: assert(~_GEN_1959);
      assert__assert_142: assert(~_GEN_1960);
      assert__assert_143: assert(~_GEN_1961);
      assert__assert_144: assert(~_GEN_1962);
      assert__assert_145: assert(~_GEN_1963);
      assert__assert_146: assert(~_GEN_1964);
      assert__assert_147: assert(~_GEN_1965);
      assert__assert_148: assert(~_GEN_1966);
      assert__assert_149: assert(~_GEN_1967);
      assert__assert_150: assert(~_GEN_1968);
      assert__assert_151: assert(~_GEN_1969);
      assert__assert_152: assert(~_GEN_1970);
      assert__assert_153: assert(~_GEN_1971);
      assert__assert_154: assert(~_GEN_1972);
      assert__assert_155: assert(~_GEN_1973);
      assert__assert_156: assert(~_GEN_1974);
      assert__assert_157: assert(~_GEN_1975);
      assert__assert_158: assert(~_GEN_1976);
      assert__assert_159: assert(~_GEN_1977);
      assert__assert_160: assert(~(|(_GEN_1978[2:1])));
      assert__assert_161: assert(~_GEN_1979);
      assert__assert_162: assert(~_GEN_1980);
      assert__assert_163: assert(~_GEN_1981);
      assert__assert_164: assert(~_GEN_1982);
      assert__assert_165: assert(~_GEN_1983);
      assert__assert_166: assert(~_GEN_1984);
      assert__assert_167: assert(~_GEN_1985);
      assert__assert_168: assert(~_GEN_1986);
      assert__assert_169: assert(~_GEN_1987);
      assert__assert_170: assert(~_GEN_1988);
      assert__assert_171: assert(~_GEN_1989);
      assert__assert_172: assert(_GEN_1991);
      assert__assert_173: assert(_GEN_1992);
    end
    if (reset) begin
      rob_pnr <= 5'h0;
      rob_pnr_lsb <= 2'h0;
      pnr_maybe_at_tail <= 1'h0;
    end
    else begin
      if (empty & _GEN_1839) begin
        rob_pnr <= rob_head;
        if (io_enq_valids_0)
          rob_pnr_lsb <= 2'h0;
        else if (io_enq_valids_1)
          rob_pnr_lsb <= 2'h1;
        else
          rob_pnr_lsb <= {1'h1, ~io_enq_valids_2};
      end
      else if (safe_to_inc & do_inc_row) begin
        rob_pnr <= rob_pnr + 5'h1;
        rob_pnr_lsb <= 2'h0;
      end
      else if (safe_to_inc & (_do_inc_row_T_4 | full & ~pnr_maybe_at_tail)) begin
        if (rob_pnr_unsafe_0)
          rob_pnr_lsb <= 2'h0;
        else if (rob_pnr_unsafe_1)
          rob_pnr_lsb <= 2'h1;
        else
          rob_pnr_lsb <= {1'h1, ~rob_pnr_unsafe_2};
      end
      else if (safe_to_inc & _io_ready_T_1 & ~empty) begin
        if (_rob_pnr_lsb_T_16[0])
          rob_pnr_lsb <= 2'h0;
        else if (_rob_pnr_lsb_T_16[1])
          rob_pnr_lsb <= 2'h1;
        else
          rob_pnr_lsb <= {1'h1, ~(_rob_pnr_lsb_T_16[2])};
      end
      else if (full & pnr_maybe_at_tail)
        rob_pnr_lsb <= 2'h0;
      pnr_maybe_at_tail <= _maybe_full_T & (do_inc_row | pnr_maybe_at_tail);
    end
    rob_unsafe__0 <= ~_GEN_22 & (_GEN_3 ? ~_GEN_21 & _GEN_7404 : ~_GEN_20 & _GEN_7404);
    rob_unsafe__1 <= ~_GEN_36 & (_GEN_3 ? ~_GEN_35 & _GEN_7405 : ~_GEN_34 & _GEN_7405);
    rob_unsafe__2 <= ~_GEN_50 & (_GEN_3 ? ~_GEN_49 & _GEN_7406 : ~_GEN_48 & _GEN_7406);
    rob_unsafe__3 <= ~_GEN_64 & (_GEN_3 ? ~_GEN_63 & _GEN_7407 : ~_GEN_62 & _GEN_7407);
    rob_unsafe__4 <= ~_GEN_78 & (_GEN_3 ? ~_GEN_77 & _GEN_7408 : ~_GEN_76 & _GEN_7408);
    rob_unsafe__5 <= ~_GEN_92 & (_GEN_3 ? ~_GEN_91 & _GEN_7409 : ~_GEN_90 & _GEN_7409);
    rob_unsafe__6 <= ~_GEN_106 & (_GEN_3 ? ~_GEN_105 & _GEN_7410 : ~_GEN_104 & _GEN_7410);
    rob_unsafe__7 <= ~_GEN_120 & (_GEN_3 ? ~_GEN_119 & _GEN_7411 : ~_GEN_118 & _GEN_7411);
    rob_unsafe__8 <= ~_GEN_134 & (_GEN_3 ? ~_GEN_133 & _GEN_7412 : ~_GEN_132 & _GEN_7412);
    rob_unsafe__9 <= ~_GEN_148 & (_GEN_3 ? ~_GEN_147 & _GEN_7413 : ~_GEN_146 & _GEN_7413);
    rob_unsafe__10 <= ~_GEN_162 & (_GEN_3 ? ~_GEN_161 & _GEN_7414 : ~_GEN_160 & _GEN_7414);
    rob_unsafe__11 <= ~_GEN_176 & (_GEN_3 ? ~_GEN_175 & _GEN_7415 : ~_GEN_174 & _GEN_7415);
    rob_unsafe__12 <= ~_GEN_190 & (_GEN_3 ? ~_GEN_189 & _GEN_7416 : ~_GEN_188 & _GEN_7416);
    rob_unsafe__13 <= ~_GEN_204 & (_GEN_3 ? ~_GEN_203 & _GEN_7417 : ~_GEN_202 & _GEN_7417);
    rob_unsafe__14 <= ~_GEN_218 & (_GEN_3 ? ~_GEN_217 & _GEN_7418 : ~_GEN_216 & _GEN_7418);
    rob_unsafe__15 <= ~_GEN_232 & (_GEN_3 ? ~_GEN_231 & _GEN_7419 : ~_GEN_230 & _GEN_7419);
    rob_unsafe__16 <= ~_GEN_246 & (_GEN_3 ? ~_GEN_245 & _GEN_7420 : ~_GEN_244 & _GEN_7420);
    rob_unsafe__17 <= ~_GEN_260 & (_GEN_3 ? ~_GEN_259 & _GEN_7421 : ~_GEN_258 & _GEN_7421);
    rob_unsafe__18 <= ~_GEN_274 & (_GEN_3 ? ~_GEN_273 & _GEN_7422 : ~_GEN_272 & _GEN_7422);
    rob_unsafe__19 <= ~_GEN_288 & (_GEN_3 ? ~_GEN_287 & _GEN_7423 : ~_GEN_286 & _GEN_7423);
    rob_unsafe__20 <= ~_GEN_302 & (_GEN_3 ? ~_GEN_301 & _GEN_7424 : ~_GEN_300 & _GEN_7424);
    rob_unsafe__21 <= ~_GEN_316 & (_GEN_3 ? ~_GEN_315 & _GEN_7425 : ~_GEN_314 & _GEN_7425);
    rob_unsafe__22 <= ~_GEN_330 & (_GEN_3 ? ~_GEN_329 & _GEN_7426 : ~_GEN_328 & _GEN_7426);
    rob_unsafe__23 <= ~_GEN_344 & (_GEN_3 ? ~_GEN_343 & _GEN_7427 : ~_GEN_342 & _GEN_7427);
    rob_unsafe__24 <= ~_GEN_358 & (_GEN_3 ? ~_GEN_357 & _GEN_7428 : ~_GEN_356 & _GEN_7428);
    rob_unsafe__25 <= ~_GEN_372 & (_GEN_3 ? ~_GEN_371 & _GEN_7429 : ~_GEN_370 & _GEN_7429);
    rob_unsafe__26 <= ~_GEN_386 & (_GEN_3 ? ~_GEN_385 & _GEN_7430 : ~_GEN_384 & _GEN_7430);
    rob_unsafe__27 <= ~_GEN_400 & (_GEN_3 ? ~_GEN_399 & _GEN_7431 : ~_GEN_398 & _GEN_7431);
    rob_unsafe__28 <= ~_GEN_414 & (_GEN_3 ? ~_GEN_413 & _GEN_7432 : ~_GEN_412 & _GEN_7432);
    rob_unsafe__29 <= ~_GEN_428 & (_GEN_3 ? ~_GEN_427 & _GEN_7433 : ~_GEN_426 & _GEN_7433);
    rob_unsafe__30 <= ~_GEN_442 & (_GEN_3 ? ~_GEN_441 & _GEN_7434 : ~_GEN_440 & _GEN_7434);
    rob_unsafe__31 <= ~_GEN_456 & (_GEN_3 ? ~_GEN_455 & _GEN_7435 : ~_GEN_454 & _GEN_7435);
    rob_unsafe_1_0 <= ~_GEN_481 & (_GEN_462 ? ~_GEN_480 & _GEN_20768 : ~_GEN_479 & _GEN_20768);
    rob_unsafe_1_1 <= ~_GEN_495 & (_GEN_462 ? ~_GEN_494 & _GEN_20769 : ~_GEN_493 & _GEN_20769);
    rob_unsafe_1_2 <= ~_GEN_509 & (_GEN_462 ? ~_GEN_508 & _GEN_20770 : ~_GEN_507 & _GEN_20770);
    rob_unsafe_1_3 <= ~_GEN_523 & (_GEN_462 ? ~_GEN_522 & _GEN_20771 : ~_GEN_521 & _GEN_20771);
    rob_unsafe_1_4 <= ~_GEN_537 & (_GEN_462 ? ~_GEN_536 & _GEN_20772 : ~_GEN_535 & _GEN_20772);
    rob_unsafe_1_5 <= ~_GEN_551 & (_GEN_462 ? ~_GEN_550 & _GEN_20773 : ~_GEN_549 & _GEN_20773);
    rob_unsafe_1_6 <= ~_GEN_565 & (_GEN_462 ? ~_GEN_564 & _GEN_20774 : ~_GEN_563 & _GEN_20774);
    rob_unsafe_1_7 <= ~_GEN_579 & (_GEN_462 ? ~_GEN_578 & _GEN_20775 : ~_GEN_577 & _GEN_20775);
    rob_unsafe_1_8 <= ~_GEN_593 & (_GEN_462 ? ~_GEN_592 & _GEN_20776 : ~_GEN_591 & _GEN_20776);
    rob_unsafe_1_9 <= ~_GEN_607 & (_GEN_462 ? ~_GEN_606 & _GEN_20777 : ~_GEN_605 & _GEN_20777);
    rob_unsafe_1_10 <= ~_GEN_621 & (_GEN_462 ? ~_GEN_620 & _GEN_20778 : ~_GEN_619 & _GEN_20778);
    rob_unsafe_1_11 <= ~_GEN_635 & (_GEN_462 ? ~_GEN_634 & _GEN_20779 : ~_GEN_633 & _GEN_20779);
    rob_unsafe_1_12 <= ~_GEN_649 & (_GEN_462 ? ~_GEN_648 & _GEN_20780 : ~_GEN_647 & _GEN_20780);
    rob_unsafe_1_13 <= ~_GEN_663 & (_GEN_462 ? ~_GEN_662 & _GEN_20781 : ~_GEN_661 & _GEN_20781);
    rob_unsafe_1_14 <= ~_GEN_677 & (_GEN_462 ? ~_GEN_676 & _GEN_20782 : ~_GEN_675 & _GEN_20782);
    rob_unsafe_1_15 <= ~_GEN_691 & (_GEN_462 ? ~_GEN_690 & _GEN_20783 : ~_GEN_689 & _GEN_20783);
    rob_unsafe_1_16 <= ~_GEN_705 & (_GEN_462 ? ~_GEN_704 & _GEN_20784 : ~_GEN_703 & _GEN_20784);
    rob_unsafe_1_17 <= ~_GEN_719 & (_GEN_462 ? ~_GEN_718 & _GEN_20785 : ~_GEN_717 & _GEN_20785);
    rob_unsafe_1_18 <= ~_GEN_733 & (_GEN_462 ? ~_GEN_732 & _GEN_20786 : ~_GEN_731 & _GEN_20786);
    rob_unsafe_1_19 <= ~_GEN_747 & (_GEN_462 ? ~_GEN_746 & _GEN_20787 : ~_GEN_745 & _GEN_20787);
    rob_unsafe_1_20 <= ~_GEN_761 & (_GEN_462 ? ~_GEN_760 & _GEN_20788 : ~_GEN_759 & _GEN_20788);
    rob_unsafe_1_21 <= ~_GEN_775 & (_GEN_462 ? ~_GEN_774 & _GEN_20789 : ~_GEN_773 & _GEN_20789);
    rob_unsafe_1_22 <= ~_GEN_789 & (_GEN_462 ? ~_GEN_788 & _GEN_20790 : ~_GEN_787 & _GEN_20790);
    rob_unsafe_1_23 <= ~_GEN_803 & (_GEN_462 ? ~_GEN_802 & _GEN_20791 : ~_GEN_801 & _GEN_20791);
    rob_unsafe_1_24 <= ~_GEN_817 & (_GEN_462 ? ~_GEN_816 & _GEN_20792 : ~_GEN_815 & _GEN_20792);
    rob_unsafe_1_25 <= ~_GEN_831 & (_GEN_462 ? ~_GEN_830 & _GEN_20793 : ~_GEN_829 & _GEN_20793);
    rob_unsafe_1_26 <= ~_GEN_845 & (_GEN_462 ? ~_GEN_844 & _GEN_20794 : ~_GEN_843 & _GEN_20794);
    rob_unsafe_1_27 <= ~_GEN_859 & (_GEN_462 ? ~_GEN_858 & _GEN_20795 : ~_GEN_857 & _GEN_20795);
    rob_unsafe_1_28 <= ~_GEN_873 & (_GEN_462 ? ~_GEN_872 & _GEN_20796 : ~_GEN_871 & _GEN_20796);
    rob_unsafe_1_29 <= ~_GEN_887 & (_GEN_462 ? ~_GEN_886 & _GEN_20797 : ~_GEN_885 & _GEN_20797);
    rob_unsafe_1_30 <= ~_GEN_901 & (_GEN_462 ? ~_GEN_900 & _GEN_20798 : ~_GEN_899 & _GEN_20798);
    rob_unsafe_1_31 <= ~_GEN_915 & (_GEN_462 ? ~_GEN_914 & _GEN_20799 : ~_GEN_913 & _GEN_20799);
    rob_unsafe_2_0 <= ~_GEN_940 & (_GEN_921 ? ~_GEN_939 & _GEN_34132 : ~_GEN_938 & _GEN_34132);
    rob_unsafe_2_1 <= ~_GEN_954 & (_GEN_921 ? ~_GEN_953 & _GEN_34133 : ~_GEN_952 & _GEN_34133);
    rob_unsafe_2_2 <= ~_GEN_968 & (_GEN_921 ? ~_GEN_967 & _GEN_34134 : ~_GEN_966 & _GEN_34134);
    rob_unsafe_2_3 <= ~_GEN_982 & (_GEN_921 ? ~_GEN_981 & _GEN_34135 : ~_GEN_980 & _GEN_34135);
    rob_unsafe_2_4 <= ~_GEN_996 & (_GEN_921 ? ~_GEN_995 & _GEN_34136 : ~_GEN_994 & _GEN_34136);
    rob_unsafe_2_5 <= ~_GEN_1010 & (_GEN_921 ? ~_GEN_1009 & _GEN_34137 : ~_GEN_1008 & _GEN_34137);
    rob_unsafe_2_6 <= ~_GEN_1024 & (_GEN_921 ? ~_GEN_1023 & _GEN_34138 : ~_GEN_1022 & _GEN_34138);
    rob_unsafe_2_7 <= ~_GEN_1038 & (_GEN_921 ? ~_GEN_1037 & _GEN_34139 : ~_GEN_1036 & _GEN_34139);
    rob_unsafe_2_8 <= ~_GEN_1052 & (_GEN_921 ? ~_GEN_1051 & _GEN_34140 : ~_GEN_1050 & _GEN_34140);
    rob_unsafe_2_9 <= ~_GEN_1066 & (_GEN_921 ? ~_GEN_1065 & _GEN_34141 : ~_GEN_1064 & _GEN_34141);
    rob_unsafe_2_10 <= ~_GEN_1080 & (_GEN_921 ? ~_GEN_1079 & _GEN_34142 : ~_GEN_1078 & _GEN_34142);
    rob_unsafe_2_11 <= ~_GEN_1094 & (_GEN_921 ? ~_GEN_1093 & _GEN_34143 : ~_GEN_1092 & _GEN_34143);
    rob_unsafe_2_12 <= ~_GEN_1108 & (_GEN_921 ? ~_GEN_1107 & _GEN_34144 : ~_GEN_1106 & _GEN_34144);
    rob_unsafe_2_13 <= ~_GEN_1122 & (_GEN_921 ? ~_GEN_1121 & _GEN_34145 : ~_GEN_1120 & _GEN_34145);
    rob_unsafe_2_14 <= ~_GEN_1136 & (_GEN_921 ? ~_GEN_1135 & _GEN_34146 : ~_GEN_1134 & _GEN_34146);
    rob_unsafe_2_15 <= ~_GEN_1150 & (_GEN_921 ? ~_GEN_1149 & _GEN_34147 : ~_GEN_1148 & _GEN_34147);
    rob_unsafe_2_16 <= ~_GEN_1164 & (_GEN_921 ? ~_GEN_1163 & _GEN_34148 : ~_GEN_1162 & _GEN_34148);
    rob_unsafe_2_17 <= ~_GEN_1178 & (_GEN_921 ? ~_GEN_1177 & _GEN_34149 : ~_GEN_1176 & _GEN_34149);
    rob_unsafe_2_18 <= ~_GEN_1192 & (_GEN_921 ? ~_GEN_1191 & _GEN_34150 : ~_GEN_1190 & _GEN_34150);
    rob_unsafe_2_19 <= ~_GEN_1206 & (_GEN_921 ? ~_GEN_1205 & _GEN_34151 : ~_GEN_1204 & _GEN_34151);
    rob_unsafe_2_20 <= ~_GEN_1220 & (_GEN_921 ? ~_GEN_1219 & _GEN_34152 : ~_GEN_1218 & _GEN_34152);
    rob_unsafe_2_21 <= ~_GEN_1234 & (_GEN_921 ? ~_GEN_1233 & _GEN_34153 : ~_GEN_1232 & _GEN_34153);
    rob_unsafe_2_22 <= ~_GEN_1248 & (_GEN_921 ? ~_GEN_1247 & _GEN_34154 : ~_GEN_1246 & _GEN_34154);
    rob_unsafe_2_23 <= ~_GEN_1262 & (_GEN_921 ? ~_GEN_1261 & _GEN_34155 : ~_GEN_1260 & _GEN_34155);
    rob_unsafe_2_24 <= ~_GEN_1276 & (_GEN_921 ? ~_GEN_1275 & _GEN_34156 : ~_GEN_1274 & _GEN_34156);
    rob_unsafe_2_25 <= ~_GEN_1290 & (_GEN_921 ? ~_GEN_1289 & _GEN_34157 : ~_GEN_1288 & _GEN_34157);
    rob_unsafe_2_26 <= ~_GEN_1304 & (_GEN_921 ? ~_GEN_1303 & _GEN_34158 : ~_GEN_1302 & _GEN_34158);
    rob_unsafe_2_27 <= ~_GEN_1318 & (_GEN_921 ? ~_GEN_1317 & _GEN_34159 : ~_GEN_1316 & _GEN_34159);
    rob_unsafe_2_28 <= ~_GEN_1332 & (_GEN_921 ? ~_GEN_1331 & _GEN_34160 : ~_GEN_1330 & _GEN_34160);
    rob_unsafe_2_29 <= ~_GEN_1346 & (_GEN_921 ? ~_GEN_1345 & _GEN_34161 : ~_GEN_1344 & _GEN_34161);
    rob_unsafe_2_30 <= ~_GEN_1360 & (_GEN_921 ? ~_GEN_1359 & _GEN_34162 : ~_GEN_1358 & _GEN_34162);
    rob_unsafe_2_31 <= ~_GEN_1374 & (_GEN_921 ? ~_GEN_1373 & _GEN_34163 : ~_GEN_1372 & _GEN_34163);
    rob_unsafe_3_0 <= ~_GEN_1399 & (_GEN_1380 ? ~_GEN_1398 & _GEN_47496 : ~_GEN_1397 & _GEN_47496);
    rob_unsafe_3_1 <= ~_GEN_1413 & (_GEN_1380 ? ~_GEN_1412 & _GEN_47497 : ~_GEN_1411 & _GEN_47497);
    rob_unsafe_3_2 <= ~_GEN_1427 & (_GEN_1380 ? ~_GEN_1426 & _GEN_47498 : ~_GEN_1425 & _GEN_47498);
    rob_unsafe_3_3 <= ~_GEN_1441 & (_GEN_1380 ? ~_GEN_1440 & _GEN_47499 : ~_GEN_1439 & _GEN_47499);
    rob_unsafe_3_4 <= ~_GEN_1455 & (_GEN_1380 ? ~_GEN_1454 & _GEN_47500 : ~_GEN_1453 & _GEN_47500);
    rob_unsafe_3_5 <= ~_GEN_1469 & (_GEN_1380 ? ~_GEN_1468 & _GEN_47501 : ~_GEN_1467 & _GEN_47501);
    rob_unsafe_3_6 <= ~_GEN_1483 & (_GEN_1380 ? ~_GEN_1482 & _GEN_47502 : ~_GEN_1481 & _GEN_47502);
    rob_unsafe_3_7 <= ~_GEN_1497 & (_GEN_1380 ? ~_GEN_1496 & _GEN_47503 : ~_GEN_1495 & _GEN_47503);
    rob_unsafe_3_8 <= ~_GEN_1511 & (_GEN_1380 ? ~_GEN_1510 & _GEN_47504 : ~_GEN_1509 & _GEN_47504);
    rob_unsafe_3_9 <= ~_GEN_1525 & (_GEN_1380 ? ~_GEN_1524 & _GEN_47505 : ~_GEN_1523 & _GEN_47505);
    rob_unsafe_3_10 <= ~_GEN_1539 & (_GEN_1380 ? ~_GEN_1538 & _GEN_47506 : ~_GEN_1537 & _GEN_47506);
    rob_unsafe_3_11 <= ~_GEN_1553 & (_GEN_1380 ? ~_GEN_1552 & _GEN_47507 : ~_GEN_1551 & _GEN_47507);
    rob_unsafe_3_12 <= ~_GEN_1567 & (_GEN_1380 ? ~_GEN_1566 & _GEN_47508 : ~_GEN_1565 & _GEN_47508);
    rob_unsafe_3_13 <= ~_GEN_1581 & (_GEN_1380 ? ~_GEN_1580 & _GEN_47509 : ~_GEN_1579 & _GEN_47509);
    rob_unsafe_3_14 <= ~_GEN_1595 & (_GEN_1380 ? ~_GEN_1594 & _GEN_47510 : ~_GEN_1593 & _GEN_47510);
    rob_unsafe_3_15 <= ~_GEN_1609 & (_GEN_1380 ? ~_GEN_1608 & _GEN_47511 : ~_GEN_1607 & _GEN_47511);
    rob_unsafe_3_16 <= ~_GEN_1623 & (_GEN_1380 ? ~_GEN_1622 & _GEN_47512 : ~_GEN_1621 & _GEN_47512);
    rob_unsafe_3_17 <= ~_GEN_1637 & (_GEN_1380 ? ~_GEN_1636 & _GEN_47513 : ~_GEN_1635 & _GEN_47513);
    rob_unsafe_3_18 <= ~_GEN_1651 & (_GEN_1380 ? ~_GEN_1650 & _GEN_47514 : ~_GEN_1649 & _GEN_47514);
    rob_unsafe_3_19 <= ~_GEN_1665 & (_GEN_1380 ? ~_GEN_1664 & _GEN_47515 : ~_GEN_1663 & _GEN_47515);
    rob_unsafe_3_20 <= ~_GEN_1679 & (_GEN_1380 ? ~_GEN_1678 & _GEN_47516 : ~_GEN_1677 & _GEN_47516);
    rob_unsafe_3_21 <= ~_GEN_1693 & (_GEN_1380 ? ~_GEN_1692 & _GEN_47517 : ~_GEN_1691 & _GEN_47517);
    rob_unsafe_3_22 <= ~_GEN_1707 & (_GEN_1380 ? ~_GEN_1706 & _GEN_47518 : ~_GEN_1705 & _GEN_47518);
    rob_unsafe_3_23 <= ~_GEN_1721 & (_GEN_1380 ? ~_GEN_1720 & _GEN_47519 : ~_GEN_1719 & _GEN_47519);
    rob_unsafe_3_24 <= ~_GEN_1735 & (_GEN_1380 ? ~_GEN_1734 & _GEN_47520 : ~_GEN_1733 & _GEN_47520);
    rob_unsafe_3_25 <= ~_GEN_1749 & (_GEN_1380 ? ~_GEN_1748 & _GEN_47521 : ~_GEN_1747 & _GEN_47521);
    rob_unsafe_3_26 <= ~_GEN_1763 & (_GEN_1380 ? ~_GEN_1762 & _GEN_47522 : ~_GEN_1761 & _GEN_47522);
    rob_unsafe_3_27 <= ~_GEN_1777 & (_GEN_1380 ? ~_GEN_1776 & _GEN_47523 : ~_GEN_1775 & _GEN_47523);
    rob_unsafe_3_28 <= ~_GEN_1791 & (_GEN_1380 ? ~_GEN_1790 & _GEN_47524 : ~_GEN_1789 & _GEN_47524);
    rob_unsafe_3_29 <= ~_GEN_1805 & (_GEN_1380 ? ~_GEN_1804 & _GEN_47525 : ~_GEN_1803 & _GEN_47525);
    rob_unsafe_3_30 <= ~_GEN_1819 & (_GEN_1380 ? ~_GEN_1818 & _GEN_47526 : ~_GEN_1817 & _GEN_47526);
    rob_unsafe_3_31 <= ~_GEN_1833 & (_GEN_1380 ? ~_GEN_1832 & _GEN_47527 : ~_GEN_1831 & _GEN_47527);
  end // always @(posedge)
endmodule

