// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

module AXI4UserYanker(
  input         clock,
                reset,
                auto_in_aw_valid,
  input  [3:0]  auto_in_aw_bits_id,
  input  [31:0] auto_in_aw_bits_addr,
  input  [7:0]  auto_in_aw_bits_len,
  input  [2:0]  auto_in_aw_bits_size,
  input  [1:0]  auto_in_aw_bits_burst,
  input         auto_in_aw_bits_lock,
  input  [3:0]  auto_in_aw_bits_cache,
  input  [2:0]  auto_in_aw_bits_prot,
  input  [3:0]  auto_in_aw_bits_qos,
                auto_in_aw_bits_echo_tl_state_size,
  input  [4:0]  auto_in_aw_bits_echo_tl_state_source,
  input         auto_in_aw_bits_echo_extra_id,
                auto_in_w_valid,
  input  [63:0] auto_in_w_bits_data,
  input  [7:0]  auto_in_w_bits_strb,
  input         auto_in_w_bits_last,
                auto_in_b_ready,
                auto_in_ar_valid,
  input  [3:0]  auto_in_ar_bits_id,
  input  [31:0] auto_in_ar_bits_addr,
  input  [7:0]  auto_in_ar_bits_len,
  input  [2:0]  auto_in_ar_bits_size,
  input  [1:0]  auto_in_ar_bits_burst,
  input         auto_in_ar_bits_lock,
  input  [3:0]  auto_in_ar_bits_cache,
  input  [2:0]  auto_in_ar_bits_prot,
  input  [3:0]  auto_in_ar_bits_qos,
                auto_in_ar_bits_echo_tl_state_size,
  input  [4:0]  auto_in_ar_bits_echo_tl_state_source,
  input         auto_in_ar_bits_echo_extra_id,
                auto_in_r_ready,
                auto_out_aw_ready,
                auto_out_w_ready,
                auto_out_b_valid,
  input  [3:0]  auto_out_b_bits_id,
  input  [1:0]  auto_out_b_bits_resp,
  input         auto_out_ar_ready,
                auto_out_r_valid,
  input  [3:0]  auto_out_r_bits_id,
  input  [63:0] auto_out_r_bits_data,
  input  [1:0]  auto_out_r_bits_resp,
  input         auto_out_r_bits_last,
  output        auto_in_aw_ready,
                auto_in_w_ready,
                auto_in_b_valid,
  output [3:0]  auto_in_b_bits_id,
  output [1:0]  auto_in_b_bits_resp,
  output [3:0]  auto_in_b_bits_echo_tl_state_size,
  output [4:0]  auto_in_b_bits_echo_tl_state_source,
  output        auto_in_b_bits_echo_extra_id,
                auto_in_ar_ready,
                auto_in_r_valid,
  output [3:0]  auto_in_r_bits_id,
  output [63:0] auto_in_r_bits_data,
  output [1:0]  auto_in_r_bits_resp,
  output [3:0]  auto_in_r_bits_echo_tl_state_size,
  output [4:0]  auto_in_r_bits_echo_tl_state_source,
  output        auto_in_r_bits_echo_extra_id,
                auto_in_r_bits_last,
                auto_out_aw_valid,
  output [3:0]  auto_out_aw_bits_id,
  output [31:0] auto_out_aw_bits_addr,
  output [7:0]  auto_out_aw_bits_len,
  output [2:0]  auto_out_aw_bits_size,
  output [1:0]  auto_out_aw_bits_burst,
  output        auto_out_aw_bits_lock,
  output [3:0]  auto_out_aw_bits_cache,
  output [2:0]  auto_out_aw_bits_prot,
  output [3:0]  auto_out_aw_bits_qos,
  output        auto_out_w_valid,
  output [63:0] auto_out_w_bits_data,
  output [7:0]  auto_out_w_bits_strb,
  output        auto_out_w_bits_last,
                auto_out_b_ready,
                auto_out_ar_valid,
  output [3:0]  auto_out_ar_bits_id,
  output [31:0] auto_out_ar_bits_addr,
  output [7:0]  auto_out_ar_bits_len,
  output [2:0]  auto_out_ar_bits_size,
  output [1:0]  auto_out_ar_bits_burst,
  output        auto_out_ar_bits_lock,
  output [3:0]  auto_out_ar_bits_cache,
  output [2:0]  auto_out_ar_bits_prot,
  output [3:0]  auto_out_ar_bits_qos,
  output        auto_out_r_ready
);

  wire       _Queue_31_io_enq_ready;
  wire       _Queue_31_io_deq_valid;
  wire [3:0] _Queue_31_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_31_io_deq_bits_tl_state_source;
  wire       _Queue_31_io_deq_bits_extra_id;
  wire       _Queue_30_io_enq_ready;
  wire       _Queue_30_io_deq_valid;
  wire [3:0] _Queue_30_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_30_io_deq_bits_tl_state_source;
  wire       _Queue_30_io_deq_bits_extra_id;
  wire       _Queue_29_io_enq_ready;
  wire       _Queue_29_io_deq_valid;
  wire [3:0] _Queue_29_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_29_io_deq_bits_tl_state_source;
  wire       _Queue_29_io_deq_bits_extra_id;
  wire       _Queue_28_io_enq_ready;
  wire       _Queue_28_io_deq_valid;
  wire [3:0] _Queue_28_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_28_io_deq_bits_tl_state_source;
  wire       _Queue_28_io_deq_bits_extra_id;
  wire       _Queue_27_io_enq_ready;
  wire       _Queue_27_io_deq_valid;
  wire [3:0] _Queue_27_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_27_io_deq_bits_tl_state_source;
  wire       _Queue_27_io_deq_bits_extra_id;
  wire       _Queue_26_io_enq_ready;
  wire       _Queue_26_io_deq_valid;
  wire [3:0] _Queue_26_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_26_io_deq_bits_tl_state_source;
  wire       _Queue_26_io_deq_bits_extra_id;
  wire       _Queue_25_io_enq_ready;
  wire       _Queue_25_io_deq_valid;
  wire [3:0] _Queue_25_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_25_io_deq_bits_tl_state_source;
  wire       _Queue_25_io_deq_bits_extra_id;
  wire       _Queue_24_io_enq_ready;
  wire       _Queue_24_io_deq_valid;
  wire [3:0] _Queue_24_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_24_io_deq_bits_tl_state_source;
  wire       _Queue_24_io_deq_bits_extra_id;
  wire       _Queue_23_io_enq_ready;
  wire       _Queue_23_io_deq_valid;
  wire [3:0] _Queue_23_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_23_io_deq_bits_tl_state_source;
  wire       _Queue_23_io_deq_bits_extra_id;
  wire       _Queue_22_io_enq_ready;
  wire       _Queue_22_io_deq_valid;
  wire [3:0] _Queue_22_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_22_io_deq_bits_tl_state_source;
  wire       _Queue_22_io_deq_bits_extra_id;
  wire       _Queue_21_io_enq_ready;
  wire       _Queue_21_io_deq_valid;
  wire [3:0] _Queue_21_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_21_io_deq_bits_tl_state_source;
  wire       _Queue_21_io_deq_bits_extra_id;
  wire       _Queue_20_io_enq_ready;
  wire       _Queue_20_io_deq_valid;
  wire [3:0] _Queue_20_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_20_io_deq_bits_tl_state_source;
  wire       _Queue_20_io_deq_bits_extra_id;
  wire       _Queue_19_io_enq_ready;
  wire       _Queue_19_io_deq_valid;
  wire [3:0] _Queue_19_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_19_io_deq_bits_tl_state_source;
  wire       _Queue_19_io_deq_bits_extra_id;
  wire       _Queue_18_io_enq_ready;
  wire       _Queue_18_io_deq_valid;
  wire [3:0] _Queue_18_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_18_io_deq_bits_tl_state_source;
  wire       _Queue_18_io_deq_bits_extra_id;
  wire       _Queue_17_io_enq_ready;
  wire       _Queue_17_io_deq_valid;
  wire [3:0] _Queue_17_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_17_io_deq_bits_tl_state_source;
  wire       _Queue_17_io_deq_bits_extra_id;
  wire       _Queue_16_io_enq_ready;
  wire       _Queue_16_io_deq_valid;
  wire [3:0] _Queue_16_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_16_io_deq_bits_tl_state_source;
  wire       _Queue_16_io_deq_bits_extra_id;
  wire       _Queue_15_io_enq_ready;
  wire       _Queue_15_io_deq_valid;
  wire [3:0] _Queue_15_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_15_io_deq_bits_tl_state_source;
  wire       _Queue_15_io_deq_bits_extra_id;
  wire       _Queue_14_io_enq_ready;
  wire       _Queue_14_io_deq_valid;
  wire [3:0] _Queue_14_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_14_io_deq_bits_tl_state_source;
  wire       _Queue_14_io_deq_bits_extra_id;
  wire       _Queue_13_io_enq_ready;
  wire       _Queue_13_io_deq_valid;
  wire [3:0] _Queue_13_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_13_io_deq_bits_tl_state_source;
  wire       _Queue_13_io_deq_bits_extra_id;
  wire       _Queue_12_io_enq_ready;
  wire       _Queue_12_io_deq_valid;
  wire [3:0] _Queue_12_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_12_io_deq_bits_tl_state_source;
  wire       _Queue_12_io_deq_bits_extra_id;
  wire       _Queue_11_io_enq_ready;
  wire       _Queue_11_io_deq_valid;
  wire [3:0] _Queue_11_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_11_io_deq_bits_tl_state_source;
  wire       _Queue_11_io_deq_bits_extra_id;
  wire       _Queue_10_io_enq_ready;
  wire       _Queue_10_io_deq_valid;
  wire [3:0] _Queue_10_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_10_io_deq_bits_tl_state_source;
  wire       _Queue_10_io_deq_bits_extra_id;
  wire       _Queue_9_io_enq_ready;
  wire       _Queue_9_io_deq_valid;
  wire [3:0] _Queue_9_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_9_io_deq_bits_tl_state_source;
  wire       _Queue_9_io_deq_bits_extra_id;
  wire       _Queue_8_io_enq_ready;
  wire       _Queue_8_io_deq_valid;
  wire [3:0] _Queue_8_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_8_io_deq_bits_tl_state_source;
  wire       _Queue_8_io_deq_bits_extra_id;
  wire       _Queue_7_io_enq_ready;
  wire       _Queue_7_io_deq_valid;
  wire [3:0] _Queue_7_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_7_io_deq_bits_tl_state_source;
  wire       _Queue_7_io_deq_bits_extra_id;
  wire       _Queue_6_io_enq_ready;
  wire       _Queue_6_io_deq_valid;
  wire [3:0] _Queue_6_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_6_io_deq_bits_tl_state_source;
  wire       _Queue_6_io_deq_bits_extra_id;
  wire       _Queue_5_io_enq_ready;
  wire       _Queue_5_io_deq_valid;
  wire [3:0] _Queue_5_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_5_io_deq_bits_tl_state_source;
  wire       _Queue_5_io_deq_bits_extra_id;
  wire       _Queue_4_io_enq_ready;
  wire       _Queue_4_io_deq_valid;
  wire [3:0] _Queue_4_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_4_io_deq_bits_tl_state_source;
  wire       _Queue_4_io_deq_bits_extra_id;
  wire       _Queue_3_io_enq_ready;
  wire       _Queue_3_io_deq_valid;
  wire [3:0] _Queue_3_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_3_io_deq_bits_tl_state_source;
  wire       _Queue_3_io_deq_bits_extra_id;
  wire       _Queue_2_io_enq_ready;
  wire       _Queue_2_io_deq_valid;
  wire [3:0] _Queue_2_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_2_io_deq_bits_tl_state_source;
  wire       _Queue_2_io_deq_bits_extra_id;
  wire       _Queue_1_io_enq_ready;
  wire       _Queue_1_io_deq_valid;
  wire [3:0] _Queue_1_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_1_io_deq_bits_tl_state_source;
  wire       _Queue_1_io_deq_bits_extra_id;
  wire       _Queue_io_enq_ready;
  wire       _Queue_io_deq_valid;
  wire [3:0] _Queue_io_deq_bits_tl_state_size;
  wire [4:0] _Queue_io_deq_bits_tl_state_source;
  wire       _Queue_io_deq_bits_extra_id;
  reg        casez_tmp;
  reg        casez_tmp_0;
  reg  [4:0] casez_tmp_1;
  reg  [3:0] casez_tmp_2;
  reg        casez_tmp_3;
  reg        casez_tmp_4;
  reg  [4:0] casez_tmp_5;
  reg  [3:0] casez_tmp_6;
  always @(*) begin
    casez (auto_in_ar_bits_id)
      4'b0000:
        casez_tmp = _Queue_io_enq_ready;
      4'b0001:
        casez_tmp = _Queue_1_io_enq_ready;
      4'b0010:
        casez_tmp = _Queue_2_io_enq_ready;
      4'b0011:
        casez_tmp = _Queue_3_io_enq_ready;
      4'b0100:
        casez_tmp = _Queue_4_io_enq_ready;
      4'b0101:
        casez_tmp = _Queue_5_io_enq_ready;
      4'b0110:
        casez_tmp = _Queue_6_io_enq_ready;
      4'b0111:
        casez_tmp = _Queue_7_io_enq_ready;
      4'b1000:
        casez_tmp = _Queue_8_io_enq_ready;
      4'b1001:
        casez_tmp = _Queue_9_io_enq_ready;
      4'b1010:
        casez_tmp = _Queue_10_io_enq_ready;
      4'b1011:
        casez_tmp = _Queue_11_io_enq_ready;
      4'b1100:
        casez_tmp = _Queue_12_io_enq_ready;
      4'b1101:
        casez_tmp = _Queue_13_io_enq_ready;
      4'b1110:
        casez_tmp = _Queue_14_io_enq_ready;
      default:
        casez_tmp = _Queue_15_io_enq_ready;
    endcase
  end // always @(*)
  always @(*) begin
    casez (auto_out_r_bits_id)
      4'b0000:
        casez_tmp_0 = _Queue_io_deq_bits_extra_id;
      4'b0001:
        casez_tmp_0 = _Queue_1_io_deq_bits_extra_id;
      4'b0010:
        casez_tmp_0 = _Queue_2_io_deq_bits_extra_id;
      4'b0011:
        casez_tmp_0 = _Queue_3_io_deq_bits_extra_id;
      4'b0100:
        casez_tmp_0 = _Queue_4_io_deq_bits_extra_id;
      4'b0101:
        casez_tmp_0 = _Queue_5_io_deq_bits_extra_id;
      4'b0110:
        casez_tmp_0 = _Queue_6_io_deq_bits_extra_id;
      4'b0111:
        casez_tmp_0 = _Queue_7_io_deq_bits_extra_id;
      4'b1000:
        casez_tmp_0 = _Queue_8_io_deq_bits_extra_id;
      4'b1001:
        casez_tmp_0 = _Queue_9_io_deq_bits_extra_id;
      4'b1010:
        casez_tmp_0 = _Queue_10_io_deq_bits_extra_id;
      4'b1011:
        casez_tmp_0 = _Queue_11_io_deq_bits_extra_id;
      4'b1100:
        casez_tmp_0 = _Queue_12_io_deq_bits_extra_id;
      4'b1101:
        casez_tmp_0 = _Queue_13_io_deq_bits_extra_id;
      4'b1110:
        casez_tmp_0 = _Queue_14_io_deq_bits_extra_id;
      default:
        casez_tmp_0 = _Queue_15_io_deq_bits_extra_id;
    endcase
  end // always @(*)
  always @(*) begin
    casez (auto_out_r_bits_id)
      4'b0000:
        casez_tmp_1 = _Queue_io_deq_bits_tl_state_source;
      4'b0001:
        casez_tmp_1 = _Queue_1_io_deq_bits_tl_state_source;
      4'b0010:
        casez_tmp_1 = _Queue_2_io_deq_bits_tl_state_source;
      4'b0011:
        casez_tmp_1 = _Queue_3_io_deq_bits_tl_state_source;
      4'b0100:
        casez_tmp_1 = _Queue_4_io_deq_bits_tl_state_source;
      4'b0101:
        casez_tmp_1 = _Queue_5_io_deq_bits_tl_state_source;
      4'b0110:
        casez_tmp_1 = _Queue_6_io_deq_bits_tl_state_source;
      4'b0111:
        casez_tmp_1 = _Queue_7_io_deq_bits_tl_state_source;
      4'b1000:
        casez_tmp_1 = _Queue_8_io_deq_bits_tl_state_source;
      4'b1001:
        casez_tmp_1 = _Queue_9_io_deq_bits_tl_state_source;
      4'b1010:
        casez_tmp_1 = _Queue_10_io_deq_bits_tl_state_source;
      4'b1011:
        casez_tmp_1 = _Queue_11_io_deq_bits_tl_state_source;
      4'b1100:
        casez_tmp_1 = _Queue_12_io_deq_bits_tl_state_source;
      4'b1101:
        casez_tmp_1 = _Queue_13_io_deq_bits_tl_state_source;
      4'b1110:
        casez_tmp_1 = _Queue_14_io_deq_bits_tl_state_source;
      default:
        casez_tmp_1 = _Queue_15_io_deq_bits_tl_state_source;
    endcase
  end // always @(*)
  always @(*) begin
    casez (auto_out_r_bits_id)
      4'b0000:
        casez_tmp_2 = _Queue_io_deq_bits_tl_state_size;
      4'b0001:
        casez_tmp_2 = _Queue_1_io_deq_bits_tl_state_size;
      4'b0010:
        casez_tmp_2 = _Queue_2_io_deq_bits_tl_state_size;
      4'b0011:
        casez_tmp_2 = _Queue_3_io_deq_bits_tl_state_size;
      4'b0100:
        casez_tmp_2 = _Queue_4_io_deq_bits_tl_state_size;
      4'b0101:
        casez_tmp_2 = _Queue_5_io_deq_bits_tl_state_size;
      4'b0110:
        casez_tmp_2 = _Queue_6_io_deq_bits_tl_state_size;
      4'b0111:
        casez_tmp_2 = _Queue_7_io_deq_bits_tl_state_size;
      4'b1000:
        casez_tmp_2 = _Queue_8_io_deq_bits_tl_state_size;
      4'b1001:
        casez_tmp_2 = _Queue_9_io_deq_bits_tl_state_size;
      4'b1010:
        casez_tmp_2 = _Queue_10_io_deq_bits_tl_state_size;
      4'b1011:
        casez_tmp_2 = _Queue_11_io_deq_bits_tl_state_size;
      4'b1100:
        casez_tmp_2 = _Queue_12_io_deq_bits_tl_state_size;
      4'b1101:
        casez_tmp_2 = _Queue_13_io_deq_bits_tl_state_size;
      4'b1110:
        casez_tmp_2 = _Queue_14_io_deq_bits_tl_state_size;
      default:
        casez_tmp_2 = _Queue_15_io_deq_bits_tl_state_size;
    endcase
  end // always @(*)
  wire       _GEN = auto_out_r_valid & auto_in_r_ready;
  wire       _GEN_0 = auto_in_ar_valid & auto_out_ar_ready;
  always @(*) begin
    casez (auto_in_aw_bits_id)
      4'b0000:
        casez_tmp_3 = _Queue_16_io_enq_ready;
      4'b0001:
        casez_tmp_3 = _Queue_17_io_enq_ready;
      4'b0010:
        casez_tmp_3 = _Queue_18_io_enq_ready;
      4'b0011:
        casez_tmp_3 = _Queue_19_io_enq_ready;
      4'b0100:
        casez_tmp_3 = _Queue_20_io_enq_ready;
      4'b0101:
        casez_tmp_3 = _Queue_21_io_enq_ready;
      4'b0110:
        casez_tmp_3 = _Queue_22_io_enq_ready;
      4'b0111:
        casez_tmp_3 = _Queue_23_io_enq_ready;
      4'b1000:
        casez_tmp_3 = _Queue_24_io_enq_ready;
      4'b1001:
        casez_tmp_3 = _Queue_25_io_enq_ready;
      4'b1010:
        casez_tmp_3 = _Queue_26_io_enq_ready;
      4'b1011:
        casez_tmp_3 = _Queue_27_io_enq_ready;
      4'b1100:
        casez_tmp_3 = _Queue_28_io_enq_ready;
      4'b1101:
        casez_tmp_3 = _Queue_29_io_enq_ready;
      4'b1110:
        casez_tmp_3 = _Queue_30_io_enq_ready;
      default:
        casez_tmp_3 = _Queue_31_io_enq_ready;
    endcase
  end // always @(*)
  always @(*) begin
    casez (auto_out_b_bits_id)
      4'b0000:
        casez_tmp_4 = _Queue_16_io_deq_bits_extra_id;
      4'b0001:
        casez_tmp_4 = _Queue_17_io_deq_bits_extra_id;
      4'b0010:
        casez_tmp_4 = _Queue_18_io_deq_bits_extra_id;
      4'b0011:
        casez_tmp_4 = _Queue_19_io_deq_bits_extra_id;
      4'b0100:
        casez_tmp_4 = _Queue_20_io_deq_bits_extra_id;
      4'b0101:
        casez_tmp_4 = _Queue_21_io_deq_bits_extra_id;
      4'b0110:
        casez_tmp_4 = _Queue_22_io_deq_bits_extra_id;
      4'b0111:
        casez_tmp_4 = _Queue_23_io_deq_bits_extra_id;
      4'b1000:
        casez_tmp_4 = _Queue_24_io_deq_bits_extra_id;
      4'b1001:
        casez_tmp_4 = _Queue_25_io_deq_bits_extra_id;
      4'b1010:
        casez_tmp_4 = _Queue_26_io_deq_bits_extra_id;
      4'b1011:
        casez_tmp_4 = _Queue_27_io_deq_bits_extra_id;
      4'b1100:
        casez_tmp_4 = _Queue_28_io_deq_bits_extra_id;
      4'b1101:
        casez_tmp_4 = _Queue_29_io_deq_bits_extra_id;
      4'b1110:
        casez_tmp_4 = _Queue_30_io_deq_bits_extra_id;
      default:
        casez_tmp_4 = _Queue_31_io_deq_bits_extra_id;
    endcase
  end // always @(*)
  always @(*) begin
    casez (auto_out_b_bits_id)
      4'b0000:
        casez_tmp_5 = _Queue_16_io_deq_bits_tl_state_source;
      4'b0001:
        casez_tmp_5 = _Queue_17_io_deq_bits_tl_state_source;
      4'b0010:
        casez_tmp_5 = _Queue_18_io_deq_bits_tl_state_source;
      4'b0011:
        casez_tmp_5 = _Queue_19_io_deq_bits_tl_state_source;
      4'b0100:
        casez_tmp_5 = _Queue_20_io_deq_bits_tl_state_source;
      4'b0101:
        casez_tmp_5 = _Queue_21_io_deq_bits_tl_state_source;
      4'b0110:
        casez_tmp_5 = _Queue_22_io_deq_bits_tl_state_source;
      4'b0111:
        casez_tmp_5 = _Queue_23_io_deq_bits_tl_state_source;
      4'b1000:
        casez_tmp_5 = _Queue_24_io_deq_bits_tl_state_source;
      4'b1001:
        casez_tmp_5 = _Queue_25_io_deq_bits_tl_state_source;
      4'b1010:
        casez_tmp_5 = _Queue_26_io_deq_bits_tl_state_source;
      4'b1011:
        casez_tmp_5 = _Queue_27_io_deq_bits_tl_state_source;
      4'b1100:
        casez_tmp_5 = _Queue_28_io_deq_bits_tl_state_source;
      4'b1101:
        casez_tmp_5 = _Queue_29_io_deq_bits_tl_state_source;
      4'b1110:
        casez_tmp_5 = _Queue_30_io_deq_bits_tl_state_source;
      default:
        casez_tmp_5 = _Queue_31_io_deq_bits_tl_state_source;
    endcase
  end // always @(*)
  always @(*) begin
    casez (auto_out_b_bits_id)
      4'b0000:
        casez_tmp_6 = _Queue_16_io_deq_bits_tl_state_size;
      4'b0001:
        casez_tmp_6 = _Queue_17_io_deq_bits_tl_state_size;
      4'b0010:
        casez_tmp_6 = _Queue_18_io_deq_bits_tl_state_size;
      4'b0011:
        casez_tmp_6 = _Queue_19_io_deq_bits_tl_state_size;
      4'b0100:
        casez_tmp_6 = _Queue_20_io_deq_bits_tl_state_size;
      4'b0101:
        casez_tmp_6 = _Queue_21_io_deq_bits_tl_state_size;
      4'b0110:
        casez_tmp_6 = _Queue_22_io_deq_bits_tl_state_size;
      4'b0111:
        casez_tmp_6 = _Queue_23_io_deq_bits_tl_state_size;
      4'b1000:
        casez_tmp_6 = _Queue_24_io_deq_bits_tl_state_size;
      4'b1001:
        casez_tmp_6 = _Queue_25_io_deq_bits_tl_state_size;
      4'b1010:
        casez_tmp_6 = _Queue_26_io_deq_bits_tl_state_size;
      4'b1011:
        casez_tmp_6 = _Queue_27_io_deq_bits_tl_state_size;
      4'b1100:
        casez_tmp_6 = _Queue_28_io_deq_bits_tl_state_size;
      4'b1101:
        casez_tmp_6 = _Queue_29_io_deq_bits_tl_state_size;
      4'b1110:
        casez_tmp_6 = _Queue_30_io_deq_bits_tl_state_size;
      default:
        casez_tmp_6 = _Queue_31_io_deq_bits_tl_state_size;
    endcase
  end // always @(*)
  wire       _GEN_1 = auto_out_b_valid & auto_in_b_ready;
  wire       _GEN_2 = auto_in_aw_valid & auto_out_aw_ready;
  Queue_17 Queue (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h0),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h0 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_io_enq_ready),
    .io_deq_valid                (_Queue_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_io_deq_bits_extra_id)
  );
  Queue_17 Queue_1 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h1),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h1 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_1_io_enq_ready),
    .io_deq_valid                (_Queue_1_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_1_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_1_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_1_io_deq_bits_extra_id)
  );
  Queue_17 Queue_2 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h2),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h2 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_2_io_enq_ready),
    .io_deq_valid                (_Queue_2_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_2_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_2_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_2_io_deq_bits_extra_id)
  );
  Queue_17 Queue_3 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h3),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h3 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_3_io_enq_ready),
    .io_deq_valid                (_Queue_3_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_3_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_3_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_3_io_deq_bits_extra_id)
  );
  Queue_21 Queue_4 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h4),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h4 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_4_io_enq_ready),
    .io_deq_valid                (_Queue_4_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_4_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_4_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_4_io_deq_bits_extra_id)
  );
  Queue_21 Queue_5 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h5),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h5 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_5_io_enq_ready),
    .io_deq_valid                (_Queue_5_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_5_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_5_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_5_io_deq_bits_extra_id)
  );
  Queue_21 Queue_6 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h6),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h6 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_6_io_enq_ready),
    .io_deq_valid                (_Queue_6_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_6_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_6_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_6_io_deq_bits_extra_id)
  );
  Queue_21 Queue_7 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h7),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h7 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_7_io_enq_ready),
    .io_deq_valid                (_Queue_7_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_7_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_7_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_7_io_deq_bits_extra_id)
  );
  Queue_21 Queue_8 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h8),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h8 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_8_io_enq_ready),
    .io_deq_valid                (_Queue_8_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_8_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_8_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_8_io_deq_bits_extra_id)
  );
  Queue_21 Queue_9 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'h9),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'h9 & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_9_io_enq_ready),
    .io_deq_valid                (_Queue_9_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_9_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_9_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_9_io_deq_bits_extra_id)
  );
  Queue_21 Queue_10 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'hA),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'hA & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_10_io_enq_ready),
    .io_deq_valid                (_Queue_10_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_10_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_10_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_10_io_deq_bits_extra_id)
  );
  Queue_21 Queue_11 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'hB),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'hB & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_11_io_enq_ready),
    .io_deq_valid                (_Queue_11_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_11_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_11_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_11_io_deq_bits_extra_id)
  );
  Queue_21 Queue_12 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'hC),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'hC & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_12_io_enq_ready),
    .io_deq_valid                (_Queue_12_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_12_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_12_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_12_io_deq_bits_extra_id)
  );
  Queue_21 Queue_13 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'hD),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'hD & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_13_io_enq_ready),
    .io_deq_valid                (_Queue_13_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_13_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_13_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_13_io_deq_bits_extra_id)
  );
  Queue_21 Queue_14 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & auto_in_ar_bits_id == 4'hE),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & auto_out_r_bits_id == 4'hE & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_14_io_enq_ready),
    .io_deq_valid                (_Queue_14_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_14_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_14_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_14_io_deq_bits_extra_id)
  );
  Queue_21 Queue_15 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_0 & (&auto_in_ar_bits_id)),
    .io_enq_bits_tl_state_size   (auto_in_ar_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_ar_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_ar_bits_echo_extra_id),
    .io_deq_ready                (_GEN & (&auto_out_r_bits_id) & auto_out_r_bits_last),
    .io_enq_ready                (_Queue_15_io_enq_ready),
    .io_deq_valid                (_Queue_15_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_15_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_15_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_15_io_deq_bits_extra_id)
  );
  Queue_17 Queue_16 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h0),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h0),
    .io_enq_ready                (_Queue_16_io_enq_ready),
    .io_deq_valid                (_Queue_16_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_16_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_16_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_16_io_deq_bits_extra_id)
  );
  Queue_17 Queue_17 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h1),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h1),
    .io_enq_ready                (_Queue_17_io_enq_ready),
    .io_deq_valid                (_Queue_17_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_17_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_17_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_17_io_deq_bits_extra_id)
  );
  Queue_17 Queue_18 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h2),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h2),
    .io_enq_ready                (_Queue_18_io_enq_ready),
    .io_deq_valid                (_Queue_18_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_18_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_18_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_18_io_deq_bits_extra_id)
  );
  Queue_17 Queue_19 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h3),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h3),
    .io_enq_ready                (_Queue_19_io_enq_ready),
    .io_deq_valid                (_Queue_19_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_19_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_19_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_19_io_deq_bits_extra_id)
  );
  Queue_21 Queue_20 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h4),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h4),
    .io_enq_ready                (_Queue_20_io_enq_ready),
    .io_deq_valid                (_Queue_20_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_20_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_20_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_20_io_deq_bits_extra_id)
  );
  Queue_21 Queue_21 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h5),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h5),
    .io_enq_ready                (_Queue_21_io_enq_ready),
    .io_deq_valid                (_Queue_21_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_21_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_21_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_21_io_deq_bits_extra_id)
  );
  Queue_21 Queue_22 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h6),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h6),
    .io_enq_ready                (_Queue_22_io_enq_ready),
    .io_deq_valid                (_Queue_22_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_22_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_22_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_22_io_deq_bits_extra_id)
  );
  Queue_21 Queue_23 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h7),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h7),
    .io_enq_ready                (_Queue_23_io_enq_ready),
    .io_deq_valid                (_Queue_23_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_23_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_23_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_23_io_deq_bits_extra_id)
  );
  Queue_21 Queue_24 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h8),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h8),
    .io_enq_ready                (_Queue_24_io_enq_ready),
    .io_deq_valid                (_Queue_24_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_24_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_24_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_24_io_deq_bits_extra_id)
  );
  Queue_21 Queue_25 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'h9),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'h9),
    .io_enq_ready                (_Queue_25_io_enq_ready),
    .io_deq_valid                (_Queue_25_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_25_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_25_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_25_io_deq_bits_extra_id)
  );
  Queue_21 Queue_26 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'hA),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'hA),
    .io_enq_ready                (_Queue_26_io_enq_ready),
    .io_deq_valid                (_Queue_26_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_26_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_26_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_26_io_deq_bits_extra_id)
  );
  Queue_21 Queue_27 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'hB),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'hB),
    .io_enq_ready                (_Queue_27_io_enq_ready),
    .io_deq_valid                (_Queue_27_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_27_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_27_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_27_io_deq_bits_extra_id)
  );
  Queue_21 Queue_28 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'hC),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'hC),
    .io_enq_ready                (_Queue_28_io_enq_ready),
    .io_deq_valid                (_Queue_28_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_28_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_28_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_28_io_deq_bits_extra_id)
  );
  Queue_21 Queue_29 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'hD),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'hD),
    .io_enq_ready                (_Queue_29_io_enq_ready),
    .io_deq_valid                (_Queue_29_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_29_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_29_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_29_io_deq_bits_extra_id)
  );
  Queue_21 Queue_30 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & auto_in_aw_bits_id == 4'hE),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & auto_out_b_bits_id == 4'hE),
    .io_enq_ready                (_Queue_30_io_enq_ready),
    .io_deq_valid                (_Queue_30_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_30_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_30_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_30_io_deq_bits_extra_id)
  );
  Queue_21 Queue_31 (
    .clock                       (clock),
    .reset                       (reset),
    .io_enq_valid                (_GEN_2 & (&auto_in_aw_bits_id)),
    .io_enq_bits_tl_state_size   (auto_in_aw_bits_echo_tl_state_size),
    .io_enq_bits_tl_state_source (auto_in_aw_bits_echo_tl_state_source),
    .io_enq_bits_extra_id        (auto_in_aw_bits_echo_extra_id),
    .io_deq_ready                (_GEN_1 & (&auto_out_b_bits_id)),
    .io_enq_ready                (_Queue_31_io_enq_ready),
    .io_deq_valid                (_Queue_31_io_deq_valid),
    .io_deq_bits_tl_state_size   (_Queue_31_io_deq_bits_tl_state_size),
    .io_deq_bits_tl_state_source (_Queue_31_io_deq_bits_tl_state_source),
    .io_deq_bits_extra_id        (_Queue_31_io_deq_bits_extra_id)
  );
  assign auto_in_aw_ready = auto_out_aw_ready & casez_tmp_3;
  assign auto_in_w_ready = auto_out_w_ready;
  assign auto_in_b_valid = auto_out_b_valid;
  assign auto_in_b_bits_id = auto_out_b_bits_id;
  assign auto_in_b_bits_resp = auto_out_b_bits_resp;
  assign auto_in_b_bits_echo_tl_state_size = casez_tmp_6;
  assign auto_in_b_bits_echo_tl_state_source = casez_tmp_5;
  assign auto_in_b_bits_echo_extra_id = casez_tmp_4;
  assign auto_in_ar_ready = auto_out_ar_ready & casez_tmp;
  assign auto_in_r_valid = auto_out_r_valid;
  assign auto_in_r_bits_id = auto_out_r_bits_id;
  assign auto_in_r_bits_data = auto_out_r_bits_data;
  assign auto_in_r_bits_resp = auto_out_r_bits_resp;
  assign auto_in_r_bits_echo_tl_state_size = casez_tmp_2;
  assign auto_in_r_bits_echo_tl_state_source = casez_tmp_1;
  assign auto_in_r_bits_echo_extra_id = casez_tmp_0;
  assign auto_in_r_bits_last = auto_out_r_bits_last;
  assign auto_out_aw_valid = auto_in_aw_valid & casez_tmp_3;
  assign auto_out_aw_bits_id = auto_in_aw_bits_id;
  assign auto_out_aw_bits_addr = auto_in_aw_bits_addr;
  assign auto_out_aw_bits_len = auto_in_aw_bits_len;
  assign auto_out_aw_bits_size = auto_in_aw_bits_size;
  assign auto_out_aw_bits_burst = auto_in_aw_bits_burst;
  assign auto_out_aw_bits_lock = auto_in_aw_bits_lock;
  assign auto_out_aw_bits_cache = auto_in_aw_bits_cache;
  assign auto_out_aw_bits_prot = auto_in_aw_bits_prot;
  assign auto_out_aw_bits_qos = auto_in_aw_bits_qos;
  assign auto_out_w_valid = auto_in_w_valid;
  assign auto_out_w_bits_data = auto_in_w_bits_data;
  assign auto_out_w_bits_strb = auto_in_w_bits_strb;
  assign auto_out_w_bits_last = auto_in_w_bits_last;
  assign auto_out_b_ready = auto_in_b_ready;
  assign auto_out_ar_valid = auto_in_ar_valid & casez_tmp;
  assign auto_out_ar_bits_id = auto_in_ar_bits_id;
  assign auto_out_ar_bits_addr = auto_in_ar_bits_addr;
  assign auto_out_ar_bits_len = auto_in_ar_bits_len;
  assign auto_out_ar_bits_size = auto_in_ar_bits_size;
  assign auto_out_ar_bits_burst = auto_in_ar_bits_burst;
  assign auto_out_ar_bits_lock = auto_in_ar_bits_lock;
  assign auto_out_ar_bits_cache = auto_in_ar_bits_cache;
  assign auto_out_ar_bits_prot = auto_in_ar_bits_prot;
  assign auto_out_ar_bits_qos = auto_in_ar_bits_qos;
  assign auto_out_r_ready = auto_in_r_ready;
endmodule

