module weights_replay_and_save_wrapper;
  weights_replay_and_save_ip weights_replay_and_save_ip (
      .clk(clk),
      .rst(rst)
  );
endmodule
