// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

module ALUExeUnit_2(
  input         clock,
                reset,
                io_req_valid,
  input  [6:0]  io_req_bits_uop_uopc,
  input         io_req_bits_uop_is_rvc,
  input  [9:0]  io_req_bits_uop_fu_code,
  input  [3:0]  io_req_bits_uop_ctrl_br_type,
  input  [1:0]  io_req_bits_uop_ctrl_op1_sel,
  input  [2:0]  io_req_bits_uop_ctrl_op2_sel,
                io_req_bits_uop_ctrl_imm_sel,
  input  [3:0]  io_req_bits_uop_ctrl_op_fcn,
  input         io_req_bits_uop_ctrl_fcn_dw,
                io_req_bits_uop_is_br,
                io_req_bits_uop_is_jalr,
                io_req_bits_uop_is_jal,
                io_req_bits_uop_is_sfb,
  input  [19:0] io_req_bits_uop_br_mask,
  input  [4:0]  io_req_bits_uop_br_tag,
  input  [5:0]  io_req_bits_uop_ftq_idx,
  input         io_req_bits_uop_edge_inst,
  input  [5:0]  io_req_bits_uop_pc_lob,
  input         io_req_bits_uop_taken,
  input  [19:0] io_req_bits_uop_imm_packed,
  input  [6:0]  io_req_bits_uop_rob_idx,
  input  [4:0]  io_req_bits_uop_ldq_idx,
                io_req_bits_uop_stq_idx,
  input  [6:0]  io_req_bits_uop_pdst,
                io_req_bits_uop_prs1,
  input         io_req_bits_uop_bypassable,
                io_req_bits_uop_is_amo,
                io_req_bits_uop_uses_stq,
  input  [1:0]  io_req_bits_uop_dst_rtype,
  input         io_req_bits_uop_fp_val,
  input  [64:0] io_req_bits_rs1_data,
                io_req_bits_rs2_data,
  input         io_req_bits_kill,
                io_ll_fresp_ready,
  input  [19:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input         io_get_ftq_pc_entry_cfi_idx_valid,
  input  [2:0]  io_get_ftq_pc_entry_cfi_idx_bits,
  input         io_get_ftq_pc_entry_start_bank,
  input  [39:0] io_get_ftq_pc_pc,
  input         io_get_ftq_pc_next_val,
  input  [39:0] io_get_ftq_pc_next_pc,
  input  [2:0]  io_fcsr_rm,
  output [9:0]  io_fu_types,
  output        io_iresp_valid,
  output [6:0]  io_iresp_bits_uop_rob_idx,
                io_iresp_bits_uop_pdst,
  output        io_iresp_bits_uop_bypassable,
                io_iresp_bits_uop_is_amo,
                io_iresp_bits_uop_uses_stq,
  output [1:0]  io_iresp_bits_uop_dst_rtype,
  output [64:0] io_iresp_bits_data,
  output        io_ll_fresp_valid,
  output [6:0]  io_ll_fresp_bits_uop_uopc,
  output [19:0] io_ll_fresp_bits_uop_br_mask,
  output [6:0]  io_ll_fresp_bits_uop_rob_idx,
  output [4:0]  io_ll_fresp_bits_uop_stq_idx,
  output [6:0]  io_ll_fresp_bits_uop_pdst,
  output        io_ll_fresp_bits_uop_is_amo,
                io_ll_fresp_bits_uop_uses_stq,
  output [1:0]  io_ll_fresp_bits_uop_dst_rtype,
  output        io_ll_fresp_bits_uop_fp_val,
  output [64:0] io_ll_fresp_bits_data,
  output        io_ll_fresp_bits_predicated,
                io_ll_fresp_bits_fflags_valid,
  output [6:0]  io_ll_fresp_bits_fflags_bits_uop_rob_idx,
  output [4:0]  io_ll_fresp_bits_fflags_bits_flags,
  output        io_bypass_0_valid,
  output [6:0]  io_bypass_0_bits_uop_pdst,
  output [1:0]  io_bypass_0_bits_uop_dst_rtype,
  output [64:0] io_bypass_0_bits_data,
  output        io_brinfo_uop_is_rvc,
  output [19:0] io_brinfo_uop_br_mask,
  output [4:0]  io_brinfo_uop_br_tag,
  output [5:0]  io_brinfo_uop_ftq_idx,
  output        io_brinfo_uop_edge_inst,
  output [5:0]  io_brinfo_uop_pc_lob,
  output [6:0]  io_brinfo_uop_rob_idx,
  output [4:0]  io_brinfo_uop_ldq_idx,
                io_brinfo_uop_stq_idx,
  output        io_brinfo_valid,
                io_brinfo_mispredict,
                io_brinfo_taken,
  output [2:0]  io_brinfo_cfi_type,
  output [1:0]  io_brinfo_pc_sel,
  output [39:0] io_brinfo_jalr_target,
  output [20:0] io_brinfo_target_offset
);

  wire        _queue_io_enq_ready;
  wire        _queue_io_empty;
  wire        _IntToFPUnit_io_resp_valid;
  wire [6:0]  _IntToFPUnit_io_resp_bits_uop_uopc;
  wire [19:0] _IntToFPUnit_io_resp_bits_uop_br_mask;
  wire [6:0]  _IntToFPUnit_io_resp_bits_uop_rob_idx;
  wire [4:0]  _IntToFPUnit_io_resp_bits_uop_stq_idx;
  wire [6:0]  _IntToFPUnit_io_resp_bits_uop_pdst;
  wire        _IntToFPUnit_io_resp_bits_uop_is_amo;
  wire        _IntToFPUnit_io_resp_bits_uop_uses_stq;
  wire [1:0]  _IntToFPUnit_io_resp_bits_uop_dst_rtype;
  wire        _IntToFPUnit_io_resp_bits_uop_fp_val;
  wire [64:0] _IntToFPUnit_io_resp_bits_data;
  wire        _IntToFPUnit_io_resp_bits_fflags_valid;
  wire [6:0]  _IntToFPUnit_io_resp_bits_fflags_bits_uop_rob_idx;
  wire [4:0]  _IntToFPUnit_io_resp_bits_fflags_bits_flags;
  wire [63:0] _ALUUnit_io_resp_bits_data;
  wire [63:0] _ALUUnit_io_bypass_0_bits_data;
  ALUUnit ALUUnit (
    .clock                             (clock),
    .reset                             (reset),
    .io_req_valid                      (io_req_valid & (io_req_bits_uop_fu_code == 10'h1 | io_req_bits_uop_fu_code == 10'h2 | io_req_bits_uop_fu_code == 10'h20 & io_req_bits_uop_uopc != 7'h6C)),
    .io_req_bits_uop_uopc              (io_req_bits_uop_uopc),
    .io_req_bits_uop_is_rvc            (io_req_bits_uop_is_rvc),
    .io_req_bits_uop_ctrl_br_type      (io_req_bits_uop_ctrl_br_type),
    .io_req_bits_uop_ctrl_op1_sel      (io_req_bits_uop_ctrl_op1_sel),
    .io_req_bits_uop_ctrl_op2_sel      (io_req_bits_uop_ctrl_op2_sel),
    .io_req_bits_uop_ctrl_imm_sel      (io_req_bits_uop_ctrl_imm_sel),
    .io_req_bits_uop_ctrl_op_fcn       (io_req_bits_uop_ctrl_op_fcn),
    .io_req_bits_uop_ctrl_fcn_dw       (io_req_bits_uop_ctrl_fcn_dw),
    .io_req_bits_uop_is_br             (io_req_bits_uop_is_br),
    .io_req_bits_uop_is_jalr           (io_req_bits_uop_is_jalr),
    .io_req_bits_uop_is_jal            (io_req_bits_uop_is_jal),
    .io_req_bits_uop_is_sfb            (io_req_bits_uop_is_sfb),
    .io_req_bits_uop_br_mask           (io_req_bits_uop_br_mask),
    .io_req_bits_uop_br_tag            (io_req_bits_uop_br_tag),
    .io_req_bits_uop_ftq_idx           (io_req_bits_uop_ftq_idx),
    .io_req_bits_uop_edge_inst         (io_req_bits_uop_edge_inst),
    .io_req_bits_uop_pc_lob            (io_req_bits_uop_pc_lob),
    .io_req_bits_uop_taken             (io_req_bits_uop_taken),
    .io_req_bits_uop_imm_packed        (io_req_bits_uop_imm_packed),
    .io_req_bits_uop_rob_idx           (io_req_bits_uop_rob_idx),
    .io_req_bits_uop_ldq_idx           (io_req_bits_uop_ldq_idx),
    .io_req_bits_uop_stq_idx           (io_req_bits_uop_stq_idx),
    .io_req_bits_uop_pdst              (io_req_bits_uop_pdst),
    .io_req_bits_uop_prs1              (io_req_bits_uop_prs1),
    .io_req_bits_uop_bypassable        (io_req_bits_uop_bypassable),
    .io_req_bits_uop_is_amo            (io_req_bits_uop_is_amo),
    .io_req_bits_uop_uses_stq          (io_req_bits_uop_uses_stq),
    .io_req_bits_uop_dst_rtype         (io_req_bits_uop_dst_rtype),
    .io_req_bits_rs1_data              (io_req_bits_rs1_data[63:0]),
    .io_req_bits_rs2_data              (io_req_bits_rs2_data[63:0]),
    .io_req_bits_kill                  (io_req_bits_kill),
    .io_brupdate_b1_resolve_mask       (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask    (io_brupdate_b1_mispredict_mask),
    .io_get_ftq_pc_entry_cfi_idx_valid (io_get_ftq_pc_entry_cfi_idx_valid),
    .io_get_ftq_pc_entry_cfi_idx_bits  (io_get_ftq_pc_entry_cfi_idx_bits),
    .io_get_ftq_pc_entry_start_bank    (io_get_ftq_pc_entry_start_bank),
    .io_get_ftq_pc_pc                  (io_get_ftq_pc_pc),
    .io_get_ftq_pc_next_val            (io_get_ftq_pc_next_val),
    .io_get_ftq_pc_next_pc             (io_get_ftq_pc_next_pc),
    .io_resp_valid                     (io_iresp_valid),
    .io_resp_bits_uop_rob_idx          (io_iresp_bits_uop_rob_idx),
    .io_resp_bits_uop_pdst             (io_iresp_bits_uop_pdst),
    .io_resp_bits_uop_bypassable       (io_iresp_bits_uop_bypassable),
    .io_resp_bits_uop_is_amo           (io_iresp_bits_uop_is_amo),
    .io_resp_bits_uop_uses_stq         (io_iresp_bits_uop_uses_stq),
    .io_resp_bits_uop_dst_rtype        (io_iresp_bits_uop_dst_rtype),
    .io_resp_bits_data                 (_ALUUnit_io_resp_bits_data),
    .io_bypass_0_valid                 (io_bypass_0_valid),
    .io_bypass_0_bits_uop_pdst         (io_bypass_0_bits_uop_pdst),
    .io_bypass_0_bits_uop_dst_rtype    (io_bypass_0_bits_uop_dst_rtype),
    .io_bypass_0_bits_data             (_ALUUnit_io_bypass_0_bits_data),
    .io_brinfo_uop_is_rvc              (io_brinfo_uop_is_rvc),
    .io_brinfo_uop_br_mask             (io_brinfo_uop_br_mask),
    .io_brinfo_uop_br_tag              (io_brinfo_uop_br_tag),
    .io_brinfo_uop_ftq_idx             (io_brinfo_uop_ftq_idx),
    .io_brinfo_uop_edge_inst           (io_brinfo_uop_edge_inst),
    .io_brinfo_uop_pc_lob              (io_brinfo_uop_pc_lob),
    .io_brinfo_uop_rob_idx             (io_brinfo_uop_rob_idx),
    .io_brinfo_uop_ldq_idx             (io_brinfo_uop_ldq_idx),
    .io_brinfo_uop_stq_idx             (io_brinfo_uop_stq_idx),
    .io_brinfo_valid                   (io_brinfo_valid),
    .io_brinfo_mispredict              (io_brinfo_mispredict),
    .io_brinfo_taken                   (io_brinfo_taken),
    .io_brinfo_cfi_type                (io_brinfo_cfi_type),
    .io_brinfo_pc_sel                  (io_brinfo_pc_sel),
    .io_brinfo_jalr_target             (io_brinfo_jalr_target),
    .io_brinfo_target_offset           (io_brinfo_target_offset)
  );
  IntToFPUnit IntToFPUnit (
    .clock                                (clock),
    .reset                                (reset),
    .io_req_valid                         (io_req_valid & io_req_bits_uop_fu_code[8]),
    .io_req_bits_uop_uopc                 (io_req_bits_uop_uopc),
    .io_req_bits_uop_br_mask              (io_req_bits_uop_br_mask),
    .io_req_bits_uop_imm_packed           (io_req_bits_uop_imm_packed),
    .io_req_bits_uop_rob_idx              (io_req_bits_uop_rob_idx),
    .io_req_bits_uop_stq_idx              (io_req_bits_uop_stq_idx),
    .io_req_bits_uop_pdst                 (io_req_bits_uop_pdst),
    .io_req_bits_uop_is_amo               (io_req_bits_uop_is_amo),
    .io_req_bits_uop_uses_stq             (io_req_bits_uop_uses_stq),
    .io_req_bits_uop_dst_rtype            (io_req_bits_uop_dst_rtype),
    .io_req_bits_uop_fp_val               (io_req_bits_uop_fp_val),
    .io_req_bits_rs1_data                 (io_req_bits_rs1_data),
    .io_req_bits_kill                     (io_req_bits_kill),
    .io_brupdate_b1_resolve_mask          (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask       (io_brupdate_b1_mispredict_mask),
    .io_fcsr_rm                           (io_fcsr_rm),
    .io_resp_valid                        (_IntToFPUnit_io_resp_valid),
    .io_resp_bits_uop_uopc                (_IntToFPUnit_io_resp_bits_uop_uopc),
    .io_resp_bits_uop_br_mask             (_IntToFPUnit_io_resp_bits_uop_br_mask),
    .io_resp_bits_uop_rob_idx             (_IntToFPUnit_io_resp_bits_uop_rob_idx),
    .io_resp_bits_uop_stq_idx             (_IntToFPUnit_io_resp_bits_uop_stq_idx),
    .io_resp_bits_uop_pdst                (_IntToFPUnit_io_resp_bits_uop_pdst),
    .io_resp_bits_uop_is_amo              (_IntToFPUnit_io_resp_bits_uop_is_amo),
    .io_resp_bits_uop_uses_stq            (_IntToFPUnit_io_resp_bits_uop_uses_stq),
    .io_resp_bits_uop_dst_rtype           (_IntToFPUnit_io_resp_bits_uop_dst_rtype),
    .io_resp_bits_uop_fp_val              (_IntToFPUnit_io_resp_bits_uop_fp_val),
    .io_resp_bits_data                    (_IntToFPUnit_io_resp_bits_data),
    .io_resp_bits_fflags_valid            (_IntToFPUnit_io_resp_bits_fflags_valid),
    .io_resp_bits_fflags_bits_uop_rob_idx (_IntToFPUnit_io_resp_bits_fflags_bits_uop_rob_idx),
    .io_resp_bits_fflags_bits_flags       (_IntToFPUnit_io_resp_bits_fflags_bits_flags)
  );
  BranchKillableQueue_9 queue (
    .clock                               (clock),
    .reset                               (reset),
    .io_enq_valid                        (_IntToFPUnit_io_resp_valid),
    .io_enq_bits_uop_uopc                (_IntToFPUnit_io_resp_bits_uop_uopc),
    .io_enq_bits_uop_br_mask             (_IntToFPUnit_io_resp_bits_uop_br_mask),
    .io_enq_bits_uop_rob_idx             (_IntToFPUnit_io_resp_bits_uop_rob_idx),
    .io_enq_bits_uop_stq_idx             (_IntToFPUnit_io_resp_bits_uop_stq_idx),
    .io_enq_bits_uop_pdst                (_IntToFPUnit_io_resp_bits_uop_pdst),
    .io_enq_bits_uop_is_amo              (_IntToFPUnit_io_resp_bits_uop_is_amo),
    .io_enq_bits_uop_uses_stq            (_IntToFPUnit_io_resp_bits_uop_uses_stq),
    .io_enq_bits_uop_dst_rtype           (_IntToFPUnit_io_resp_bits_uop_dst_rtype),
    .io_enq_bits_uop_fp_val              (_IntToFPUnit_io_resp_bits_uop_fp_val),
    .io_enq_bits_data                    (_IntToFPUnit_io_resp_bits_data),
    .io_enq_bits_fflags_valid            (_IntToFPUnit_io_resp_bits_fflags_valid),
    .io_enq_bits_fflags_bits_uop_rob_idx (_IntToFPUnit_io_resp_bits_fflags_bits_uop_rob_idx),
    .io_enq_bits_fflags_bits_flags       (_IntToFPUnit_io_resp_bits_fflags_bits_flags),
    .io_deq_ready                        (io_ll_fresp_ready),
    .io_brupdate_b1_resolve_mask         (io_brupdate_b1_resolve_mask),
    .io_brupdate_b1_mispredict_mask      (io_brupdate_b1_mispredict_mask),
    .io_flush                            (io_req_bits_kill),
    .io_enq_ready                        (_queue_io_enq_ready),
    .io_deq_valid                        (io_ll_fresp_valid),
    .io_deq_bits_uop_uopc                (io_ll_fresp_bits_uop_uopc),
    .io_deq_bits_uop_br_mask             (io_ll_fresp_bits_uop_br_mask),
    .io_deq_bits_uop_rob_idx             (io_ll_fresp_bits_uop_rob_idx),
    .io_deq_bits_uop_stq_idx             (io_ll_fresp_bits_uop_stq_idx),
    .io_deq_bits_uop_pdst                (io_ll_fresp_bits_uop_pdst),
    .io_deq_bits_uop_is_amo              (io_ll_fresp_bits_uop_is_amo),
    .io_deq_bits_uop_uses_stq            (io_ll_fresp_bits_uop_uses_stq),
    .io_deq_bits_uop_dst_rtype           (io_ll_fresp_bits_uop_dst_rtype),
    .io_deq_bits_uop_fp_val              (io_ll_fresp_bits_uop_fp_val),
    .io_deq_bits_data                    (io_ll_fresp_bits_data),
    .io_deq_bits_predicated              (io_ll_fresp_bits_predicated),
    .io_deq_bits_fflags_valid            (io_ll_fresp_bits_fflags_valid),
    .io_deq_bits_fflags_bits_uop_rob_idx (io_ll_fresp_bits_fflags_bits_uop_rob_idx),
    .io_deq_bits_fflags_bits_flags       (io_ll_fresp_bits_fflags_bits_flags),
    .io_empty                            (_queue_io_empty)
  );
  assign io_fu_types = {1'h0, _queue_io_empty, 8'h3};
  assign io_iresp_bits_data = {1'h0, _ALUUnit_io_resp_bits_data};
  assign io_bypass_0_bits_data = {1'h0, _ALUUnit_io_bypass_0_bits_data};
endmodule

