// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

// VCS coverage exclude_file
module LSU_assert(
  input        io_core_brupdate_b2_mispredict,
               _stq_stq_execute_head_valid_1,
  input [4:0]  stq_tail,
               stq_execute_head,
               stq_head,
               ldq_tail,
               io_core_dis_uops_0_bits_ldq_idx,
  input        ldq_31_valid,
               ldq_30_valid,
               ldq_29_valid,
               ldq_28_valid,
               ldq_27_valid,
               ldq_26_valid,
               ldq_25_valid,
               ldq_24_valid,
               ldq_23_valid,
               ldq_22_valid,
               ldq_21_valid,
               ldq_20_valid,
               ldq_19_valid,
               ldq_18_valid,
               ldq_17_valid,
               ldq_16_valid,
               ldq_15_valid,
               ldq_14_valid,
               ldq_13_valid,
               ldq_12_valid,
               ldq_11_valid,
               ldq_10_valid,
               ldq_9_valid,
               ldq_8_valid,
               ldq_7_valid,
               ldq_6_valid,
               ldq_5_valid,
               ldq_4_valid,
               ldq_3_valid,
               ldq_2_valid,
               ldq_1_valid,
               ldq_0_valid,
  input [4:0]  io_core_dis_uops_0_bits_stq_idx,
  input        stq_31_valid,
               stq_30_valid,
               stq_29_valid,
               stq_28_valid,
               stq_27_valid,
               stq_26_valid,
               stq_25_valid,
               stq_24_valid,
               stq_23_valid,
               stq_22_valid,
               stq_21_valid,
               stq_20_valid,
               stq_19_valid,
               stq_18_valid,
               stq_17_valid,
               stq_16_valid,
               stq_15_valid,
               stq_14_valid,
               stq_13_valid,
               stq_12_valid,
               stq_11_valid,
               stq_10_valid,
               stq_9_valid,
               stq_8_valid,
               stq_7_valid,
               stq_6_valid,
               stq_5_valid,
               stq_4_valid,
               stq_3_valid,
               stq_2_valid,
               stq_1_valid,
               stq_0_valid,
               dis_ld_val,
               dis_st_val,
  input [4:0]  _GEN,
               io_core_dis_uops_1_bits_ldq_idx,
               _ldq_T_35_bits_youngest_stq_idx,
               io_core_dis_uops_1_bits_stq_idx,
  input        dis_ld_val_1,
               dis_st_val_1,
  input [4:0]  _GEN_0,
               io_core_dis_uops_2_bits_ldq_idx,
               _ldq_T_75_bits_youngest_stq_idx,
               io_core_dis_uops_2_bits_stq_idx,
  input        dis_ld_val_2,
               dis_st_val_2,
  input [4:0]  _GEN_1,
               io_core_dis_uops_3_bits_ldq_idx,
               _ldq_T_115_bits_youngest_stq_idx,
               io_core_dis_uops_3_bits_stq_idx,
  input        dis_ld_val_3,
               dis_st_val_3,
               exe_req_0_valid,
               will_fire_std_incoming_0,
               will_fire_sfence_0,
               _exe_cmd_T,
               will_fire_sta_incoming_0,
               exe_req_1_valid,
               will_fire_std_incoming_1,
               will_fire_sfence_1,
               _exe_cmd_T_7,
               will_fire_sta_incoming_1,
               _GEN_2,
  input [4:0]  hella_req_cmd,
  input        exe_tlb_valid_0,
               _exe_tlb_uop_T_2,
               io_core_exe_1_req_bits_sfence_valid,
               io_core_exe_1_req_bits_uop_is_fence,
               io_core_exe_0_req_bits_uop_is_fence,
               exe_req_0_bits_mxcpt_valid,
               mem_incoming_uop_out_ctrl_is_sta,
               mem_incoming_uop_out_ctrl_is_load,
               can_fire_load_incoming_0,
               will_fire_stad_incoming_0,
               exe_tlb_valid_1,
               _exe_tlb_uop_T_9,
               will_fire_load_retry_1,
               will_fire_sta_retry_1,
  input [4:0]  stq_retry_idx,
  input        stq_31_bits_uop_is_fence,
               stq_30_bits_uop_is_fence,
               stq_29_bits_uop_is_fence,
               stq_28_bits_uop_is_fence,
               stq_27_bits_uop_is_fence,
               stq_26_bits_uop_is_fence,
               stq_25_bits_uop_is_fence,
               stq_24_bits_uop_is_fence,
               stq_23_bits_uop_is_fence,
               stq_22_bits_uop_is_fence,
               stq_21_bits_uop_is_fence,
               stq_20_bits_uop_is_fence,
               stq_19_bits_uop_is_fence,
               stq_18_bits_uop_is_fence,
               stq_17_bits_uop_is_fence,
               stq_16_bits_uop_is_fence,
               stq_15_bits_uop_is_fence,
               stq_14_bits_uop_is_fence,
               stq_13_bits_uop_is_fence,
               stq_12_bits_uop_is_fence,
               stq_11_bits_uop_is_fence,
               stq_10_bits_uop_is_fence,
               stq_9_bits_uop_is_fence,
               stq_8_bits_uop_is_fence,
               stq_7_bits_uop_is_fence,
               stq_6_bits_uop_is_fence,
               stq_5_bits_uop_is_fence,
               stq_4_bits_uop_is_fence,
               stq_3_bits_uop_is_fence,
               stq_2_bits_uop_is_fence,
               stq_1_bits_uop_is_fence,
               stq_0_bits_uop_is_fence,
  input [4:0]  ldq_retry_idx,
  input        clock,
               _GEN_3,
               io_core_dis_uops_3_bits_is_fence,
               _GEN_4,
               io_core_dis_uops_2_bits_is_fence,
               _GEN_5,
               io_core_dis_uops_1_bits_is_fence,
               _GEN_6,
               io_core_dis_uops_0_bits_is_fence,
               _GEN_7,
               _GEN_8,
               _GEN_9,
               _GEN_10,
               _GEN_11,
               _GEN_12,
               _GEN_13,
               _GEN_14,
               _GEN_15,
               _GEN_16,
               _GEN_17,
               _GEN_18,
               _GEN_19,
               _GEN_20,
               _GEN_21,
               _GEN_22,
               _GEN_23,
               _GEN_24,
               _GEN_25,
               _GEN_26,
               _GEN_27,
               _GEN_28,
               _GEN_29,
               _GEN_30,
               _GEN_31,
               _GEN_32,
               _GEN_33,
               _GEN_34,
               _GEN_35,
               _GEN_36,
               _GEN_37,
               _GEN_38,
               _GEN_39,
               _GEN_40,
               _GEN_41,
               _GEN_42,
               _GEN_43,
               _GEN_44,
               _GEN_45,
               _GEN_46,
               _GEN_47,
               _GEN_48,
               _GEN_49,
               _GEN_50,
               _GEN_51,
               _GEN_52,
               _GEN_53,
               _GEN_54,
               _GEN_55,
               _GEN_56,
               _GEN_57,
               _GEN_58,
               _GEN_59,
               _GEN_60,
               _GEN_61,
               _GEN_62,
               _GEN_63,
               _GEN_64,
               _GEN_65,
               _GEN_66,
               _GEN_67,
               _GEN_68,
               _GEN_69,
               _GEN_70,
               _GEN_71,
               _GEN_72,
               _GEN_73,
               _GEN_74,
               _GEN_75,
               _GEN_76,
               _GEN_77,
               _GEN_78,
               _GEN_79,
               _GEN_80,
               _GEN_81,
               _GEN_82,
               _GEN_83,
               _GEN_84,
               _GEN_85,
               _GEN_86,
               _GEN_87,
               _GEN_88,
               _GEN_89,
               _GEN_90,
               _GEN_91,
               _GEN_92,
               _GEN_93,
               _GEN_94,
               _GEN_95,
               _GEN_96,
               _GEN_97,
               _GEN_98,
               _GEN_99,
               _GEN_100,
               _GEN_101,
               _GEN_102,
               _GEN_103,
               _GEN_104,
               _GEN_105,
               _GEN_106,
               _GEN_107,
               _GEN_108,
               _GEN_109,
               _GEN_110,
               _GEN_111,
               _GEN_112,
               _GEN_113,
               _GEN_114,
               _GEN_115,
               _GEN_116,
               _GEN_117,
               _GEN_118,
               _GEN_119,
               _GEN_120,
               _GEN_121,
               _GEN_122,
               _GEN_123,
               _GEN_124,
               _GEN_125,
               _GEN_126,
               _GEN_127,
               _GEN_128,
               _GEN_129,
               _GEN_130,
               io_core_exe_0_req_bits_sfence_valid,
               exe_req_1_bits_mxcpt_valid,
               exe_req_1_bits_uop_ctrl_is_sta,
               io_core_dis_uops_3_bits_ctrl_is_sta,
               io_core_dis_uops_2_bits_ctrl_is_sta,
               io_core_dis_uops_1_bits_ctrl_is_sta,
               io_core_dis_uops_0_bits_ctrl_is_sta,
               _GEN_131,
               _GEN_132,
               _GEN_133,
               _GEN_134,
               _GEN_135,
               _GEN_136,
               _GEN_137,
               _GEN_138,
               _GEN_139,
               _GEN_140,
               _GEN_141,
               _GEN_142,
               _GEN_143,
               _GEN_144,
               _GEN_145,
               _GEN_146,
               _GEN_147,
               _GEN_148,
               _GEN_149,
               _GEN_150,
               _GEN_151,
               _GEN_152,
               _GEN_153,
               _GEN_154,
               _GEN_155,
               _GEN_156,
               _GEN_157,
               _GEN_158,
               _GEN_159,
               _GEN_160,
               _GEN_161,
               _GEN_162,
               _GEN_163,
               _GEN_164,
               _GEN_165,
               _GEN_166,
               _GEN_167,
               _GEN_168,
               _GEN_169,
               _GEN_170,
               _GEN_171,
               _GEN_172,
               _GEN_173,
               _GEN_174,
               _GEN_175,
               _GEN_176,
               _GEN_177,
               _GEN_178,
               _GEN_179,
               _GEN_180,
               _GEN_181,
               _GEN_182,
               _GEN_183,
               _GEN_184,
               _GEN_185,
               _GEN_186,
               _GEN_187,
               _GEN_188,
               _GEN_189,
               _GEN_190,
               _GEN_191,
               _GEN_192,
               _GEN_193,
               _GEN_194,
               _GEN_195,
               _GEN_196,
               _GEN_197,
               _GEN_198,
               _GEN_199,
               _GEN_200,
               _GEN_201,
               _GEN_202,
               _GEN_203,
               _GEN_204,
               _GEN_205,
               _GEN_206,
               _GEN_207,
               _GEN_208,
               _GEN_209,
               _GEN_210,
               _GEN_211,
               _GEN_212,
               _GEN_213,
               _GEN_214,
               _GEN_215,
               _GEN_216,
               _GEN_217,
               _GEN_218,
               _GEN_219,
               _GEN_220,
               _GEN_221,
               _GEN_222,
               _GEN_223,
               _GEN_224,
               _GEN_225,
               _GEN_226,
               _GEN_227,
               _GEN_228,
               _GEN_229,
               _GEN_230,
               _GEN_231,
               _GEN_232,
               _GEN_233,
               _GEN_234,
               _GEN_235,
               _GEN_236,
               _GEN_237,
               _GEN_238,
               _GEN_239,
               _GEN_240,
               _GEN_241,
               _GEN_242,
               _GEN_243,
               _GEN_244,
               _GEN_245,
               _GEN_246,
               _GEN_247,
               _GEN_248,
               _GEN_249,
               _GEN_250,
               _GEN_251,
               _GEN_252,
               _GEN_253,
               _GEN_254,
               _GEN_255,
               _GEN_256,
               _GEN_257,
               _GEN_258,
               _GEN_259,
               exe_req_1_bits_uop_ctrl_is_load,
               io_core_dis_uops_3_bits_ctrl_is_load,
               io_core_dis_uops_2_bits_ctrl_is_load,
               io_core_dis_uops_1_bits_ctrl_is_load,
               io_core_dis_uops_0_bits_ctrl_is_load,
               can_fire_load_incoming_1,
               will_fire_stad_incoming_1,
               exe_req_0_bits_sfence_valid,
  input [31:0] exe_tlb_paddr_0,
               dtlb_io_resp_0_paddr,
  input        mem_xcpt_uops_0_uses_ldq,
               exe_tlb_uop_0_uses_stq,
               exe_req_1_bits_sfence_valid,
  input [31:0] exe_tlb_paddr_1,
               dtlb_io_resp_1_paddr,
  input        mem_xcpt_uops_1_uses_ldq,
               exe_tlb_uop_1_uses_stq,
  input [4:0]  ldq_incoming_idx_0,
  input        ldq_31_bits_executed,
               ldq_30_bits_executed,
               ldq_29_bits_executed,
               ldq_28_bits_executed,
               ldq_27_bits_executed,
               ldq_26_bits_executed,
               ldq_25_bits_executed,
               ldq_24_bits_executed,
               ldq_23_bits_executed,
               ldq_22_bits_executed,
               ldq_21_bits_executed,
               ldq_20_bits_executed,
               ldq_19_bits_executed,
               ldq_18_bits_executed,
               ldq_17_bits_executed,
               ldq_16_bits_executed,
               ldq_15_bits_executed,
               ldq_14_bits_executed,
               ldq_13_bits_executed,
               ldq_12_bits_executed,
               ldq_11_bits_executed,
               ldq_10_bits_executed,
               ldq_9_bits_executed,
               ldq_8_bits_executed,
               ldq_7_bits_executed,
               ldq_6_bits_executed,
               ldq_5_bits_executed,
               ldq_4_bits_executed,
               ldq_3_bits_executed,
               ldq_2_bits_executed,
               ldq_1_bits_executed,
               ldq_0_bits_executed,
               ldq_31_bits_addr_valid,
               ldq_30_bits_addr_valid,
               ldq_29_bits_addr_valid,
               ldq_28_bits_addr_valid,
               ldq_27_bits_addr_valid,
               ldq_26_bits_addr_valid,
               ldq_25_bits_addr_valid,
               ldq_24_bits_addr_valid,
               ldq_23_bits_addr_valid,
               ldq_22_bits_addr_valid,
               ldq_21_bits_addr_valid,
               ldq_20_bits_addr_valid,
               ldq_19_bits_addr_valid,
               ldq_18_bits_addr_valid,
               ldq_17_bits_addr_valid,
               ldq_16_bits_addr_valid,
               ldq_15_bits_addr_valid,
               ldq_14_bits_addr_valid,
               ldq_13_bits_addr_valid,
               ldq_12_bits_addr_valid,
               ldq_11_bits_addr_valid,
               ldq_10_bits_addr_valid,
               ldq_9_bits_addr_valid,
               ldq_8_bits_addr_valid,
               ldq_7_bits_addr_valid,
               ldq_6_bits_addr_valid,
               ldq_5_bits_addr_valid,
               ldq_4_bits_addr_valid,
               ldq_3_bits_addr_valid,
               ldq_2_bits_addr_valid,
               ldq_1_bits_addr_valid,
               ldq_0_bits_addr_valid,
               stq_incoming_e_0_bits_addr_valid,
  input [4:0]  sidx,
  input        stq_31_bits_data_valid,
               stq_30_bits_data_valid,
               stq_29_bits_data_valid,
               stq_28_bits_data_valid,
               stq_27_bits_data_valid,
               stq_26_bits_data_valid,
               stq_25_bits_data_valid,
               stq_24_bits_data_valid,
               stq_23_bits_data_valid,
               stq_22_bits_data_valid,
               stq_21_bits_data_valid,
               stq_20_bits_data_valid,
               stq_19_bits_data_valid,
               stq_18_bits_data_valid,
               stq_17_bits_data_valid,
               stq_16_bits_data_valid,
               stq_15_bits_data_valid,
               stq_14_bits_data_valid,
               stq_13_bits_data_valid,
               stq_12_bits_data_valid,
               stq_11_bits_data_valid,
               stq_10_bits_data_valid,
               stq_9_bits_data_valid,
               stq_8_bits_data_valid,
               stq_7_bits_data_valid,
               stq_6_bits_data_valid,
               stq_5_bits_data_valid,
               stq_4_bits_data_valid,
               stq_3_bits_data_valid,
               stq_2_bits_data_valid,
               stq_1_bits_data_valid,
               stq_0_bits_data_valid,
  input [4:0]  ldq_incoming_idx_1,
  input        mem_ldq_wakeup_e_out_bits_addr_is_virtual,
               mem_ldq_wakeup_e_out_bits_executed,
               _GEN_140251,
               _GEN_140205,
               stq_incoming_e_1_bits_addr_valid,
  input [4:0]  sidx_1,
  input        _GEN_260,
               _GEN_261,
  input [4:0]  io_dmem_nack_0_bits_uop_ldq_idx,
  input        io_dmem_nack_0_bits_uop_uses_stq,
               io_dmem_resp_0_bits_is_hella,
               send_iresp,
               send_fresp,
  input [4:0]  io_dmem_nack_1_bits_uop_ldq_idx,
  input        io_dmem_nack_1_bits_uop_uses_stq,
               io_dmem_resp_1_bits_is_hella,
               send_iresp_1,
               send_fresp_1,
               stq_0_bits_committed,
  input [19:0] _GEN_262,
  input        stq_1_bits_committed,
  input [19:0] _GEN_263,
  input        stq_2_bits_committed,
  input [19:0] _GEN_264,
  input        stq_3_bits_committed,
  input [19:0] _GEN_265,
  input        stq_4_bits_committed,
  input [19:0] _GEN_266,
  input        stq_5_bits_committed,
  input [19:0] _GEN_267,
  input        stq_6_bits_committed,
  input [19:0] _GEN_268,
  input        stq_7_bits_committed,
  input [19:0] _GEN_269,
  input        stq_8_bits_committed,
  input [19:0] _GEN_270,
  input        stq_9_bits_committed,
  input [19:0] _GEN_271,
  input        stq_10_bits_committed,
  input [19:0] _GEN_272,
  input        stq_11_bits_committed,
  input [19:0] _GEN_273,
  input        stq_12_bits_committed,
  input [19:0] _GEN_274,
  input        stq_13_bits_committed,
  input [19:0] _GEN_275,
  input        stq_14_bits_committed,
  input [19:0] _GEN_276,
  input        stq_15_bits_committed,
  input [19:0] _GEN_277,
  input        stq_16_bits_committed,
  input [19:0] _GEN_278,
  input        stq_17_bits_committed,
  input [19:0] _GEN_279,
  input        stq_18_bits_committed,
  input [19:0] _GEN_280,
  input        stq_19_bits_committed,
  input [19:0] _GEN_281,
  input        stq_20_bits_committed,
  input [19:0] _GEN_282,
  input        stq_21_bits_committed,
  input [19:0] _GEN_283,
  input        stq_22_bits_committed,
  input [19:0] _GEN_284,
  input        stq_23_bits_committed,
  input [19:0] _GEN_285,
  input        stq_24_bits_committed,
  input [19:0] _GEN_286,
  input        stq_25_bits_committed,
  input [19:0] _GEN_287,
  input        stq_26_bits_committed,
  input [19:0] _GEN_288,
  input        stq_27_bits_committed,
  input [19:0] _GEN_289,
  input        stq_28_bits_committed,
  input [19:0] _GEN_290,
  input        stq_29_bits_committed,
  input [19:0] _GEN_291,
  input        stq_30_bits_committed,
  input [19:0] _GEN_292,
  input        stq_31_bits_committed,
  input [19:0] _GEN_293,
  input [4:0]  idx,
  input        ldq_31_bits_succeeded,
               ldq_30_bits_succeeded,
               ldq_29_bits_succeeded,
               ldq_28_bits_succeeded,
               ldq_27_bits_succeeded,
               ldq_26_bits_succeeded,
               ldq_25_bits_succeeded,
               ldq_24_bits_succeeded,
               ldq_23_bits_succeeded,
               ldq_22_bits_succeeded,
               ldq_21_bits_succeeded,
               ldq_20_bits_succeeded,
               ldq_19_bits_succeeded,
               ldq_18_bits_succeeded,
               ldq_17_bits_succeeded,
               ldq_16_bits_succeeded,
               ldq_15_bits_succeeded,
               ldq_14_bits_succeeded,
               ldq_13_bits_succeeded,
               ldq_12_bits_succeeded,
               ldq_11_bits_succeeded,
               ldq_10_bits_succeeded,
               ldq_9_bits_succeeded,
               ldq_8_bits_succeeded,
               ldq_7_bits_succeeded,
               ldq_6_bits_succeeded,
               ldq_5_bits_succeeded,
               ldq_4_bits_succeeded,
               ldq_3_bits_succeeded,
               ldq_2_bits_succeeded,
               ldq_1_bits_succeeded,
               ldq_0_bits_succeeded,
               ldq_31_bits_forward_std_val,
               ldq_30_bits_forward_std_val,
               ldq_29_bits_forward_std_val,
               ldq_28_bits_forward_std_val,
               ldq_27_bits_forward_std_val,
               ldq_26_bits_forward_std_val,
               ldq_25_bits_forward_std_val,
               ldq_24_bits_forward_std_val,
               ldq_23_bits_forward_std_val,
               ldq_22_bits_forward_std_val,
               ldq_21_bits_forward_std_val,
               ldq_20_bits_forward_std_val,
               ldq_19_bits_forward_std_val,
               ldq_18_bits_forward_std_val,
               ldq_17_bits_forward_std_val,
               ldq_16_bits_forward_std_val,
               ldq_15_bits_forward_std_val,
               ldq_14_bits_forward_std_val,
               ldq_13_bits_forward_std_val,
               ldq_12_bits_forward_std_val,
               ldq_11_bits_forward_std_val,
               ldq_10_bits_forward_std_val,
               ldq_9_bits_forward_std_val,
               ldq_8_bits_forward_std_val,
               ldq_7_bits_forward_std_val,
               ldq_6_bits_forward_std_val,
               ldq_5_bits_forward_std_val,
               ldq_4_bits_forward_std_val,
               ldq_3_bits_forward_std_val,
               ldq_2_bits_forward_std_val,
               ldq_1_bits_forward_std_val,
               ldq_0_bits_forward_std_val,
  input [4:0]  idx_1,
               idx_2,
               idx_3,
  input        reset,
               mem_xcpt_valids_0,
               mem_xcpt_valids_1,
               _stq_idx_T,
               _GEN_294,
               will_fire_load_wakeup_1,
               will_fire_hella_incoming_1,
               will_fire_hella_wakeup_1,
               _GEN_295,
               _GEN_296,
               _stq_bits_data_bits_T_2,
               _GEN_297,
               io_dmem_nack_0_bits_uop_uses_ldq,
               io_dmem_nack_0_valid,
               io_dmem_nack_0_bits_is_hella,
               _GEN_298,
               io_dmem_resp_0_valid,
               io_dmem_resp_0_bits_uop_uses_stq,
               io_dmem_resp_0_bits_uop_uses_ldq,
               _GEN_299,
               io_dmem_nack_1_bits_uop_uses_ldq,
               io_dmem_nack_1_valid,
               io_dmem_nack_1_bits_is_hella,
               _GEN_300,
               io_dmem_resp_1_valid,
               io_dmem_resp_1_bits_uop_uses_stq,
               io_dmem_resp_1_bits_uop_uses_ldq,
               commit_load,
               commit_store,
               commit_load_1,
               commit_store_1,
               commit_load_2,
               commit_store_2,
               commit_load_3,
               commit_store_3
);

  reg  casez_tmp;
  reg  casez_tmp_0;
  reg  casez_tmp_1;
  reg  casez_tmp_2;
  reg  casez_tmp_3;
  reg  casez_tmp_4;
  reg  casez_tmp_5;
  reg  casez_tmp_6;
  reg  casez_tmp_7;
  reg  casez_tmp_8;
  reg  casez_tmp_9;
  reg  casez_tmp_10;
  reg  casez_tmp_11;
  reg  casez_tmp_12;
  reg  casez_tmp_13;
  reg  casez_tmp_14;
  reg  casez_tmp_15;
  reg  casez_tmp_16;
  reg  casez_tmp_17;
  reg  casez_tmp_18;
  reg  casez_tmp_19;
  reg  casez_tmp_20;
  reg  casez_tmp_21;
  reg  casez_tmp_22;
  reg  casez_tmp_23;
  reg  casez_tmp_24;
  reg  casez_tmp_25;
  reg  casez_tmp_26;
  reg  casez_tmp_27;
  reg  casez_tmp_28;
  reg  casez_tmp_29;
  reg  casez_tmp_30;
  reg  casez_tmp_31;
  reg  casez_tmp_32;
  reg  casez_tmp_33;
  reg  casez_tmp_34;
  reg  casez_tmp_35;
  reg  casez_tmp_36;
  reg  casez_tmp_37;
  reg  ldq_0_bits_uop_ctrl_is_load;
  reg  ldq_0_bits_uop_ctrl_is_sta;
  reg  ldq_0_bits_uop_is_fence;
  reg  ldq_1_bits_uop_ctrl_is_load;
  reg  ldq_1_bits_uop_ctrl_is_sta;
  reg  ldq_1_bits_uop_is_fence;
  reg  ldq_2_bits_uop_ctrl_is_load;
  reg  ldq_2_bits_uop_ctrl_is_sta;
  reg  ldq_2_bits_uop_is_fence;
  reg  ldq_3_bits_uop_ctrl_is_load;
  reg  ldq_3_bits_uop_ctrl_is_sta;
  reg  ldq_3_bits_uop_is_fence;
  reg  ldq_4_bits_uop_ctrl_is_load;
  reg  ldq_4_bits_uop_ctrl_is_sta;
  reg  ldq_4_bits_uop_is_fence;
  reg  ldq_5_bits_uop_ctrl_is_load;
  reg  ldq_5_bits_uop_ctrl_is_sta;
  reg  ldq_5_bits_uop_is_fence;
  reg  ldq_6_bits_uop_ctrl_is_load;
  reg  ldq_6_bits_uop_ctrl_is_sta;
  reg  ldq_6_bits_uop_is_fence;
  reg  ldq_7_bits_uop_ctrl_is_load;
  reg  ldq_7_bits_uop_ctrl_is_sta;
  reg  ldq_7_bits_uop_is_fence;
  reg  ldq_8_bits_uop_ctrl_is_load;
  reg  ldq_8_bits_uop_ctrl_is_sta;
  reg  ldq_8_bits_uop_is_fence;
  reg  ldq_9_bits_uop_ctrl_is_load;
  reg  ldq_9_bits_uop_ctrl_is_sta;
  reg  ldq_9_bits_uop_is_fence;
  reg  ldq_10_bits_uop_ctrl_is_load;
  reg  ldq_10_bits_uop_ctrl_is_sta;
  reg  ldq_10_bits_uop_is_fence;
  reg  ldq_11_bits_uop_ctrl_is_load;
  reg  ldq_11_bits_uop_ctrl_is_sta;
  reg  ldq_11_bits_uop_is_fence;
  reg  ldq_12_bits_uop_ctrl_is_load;
  reg  ldq_12_bits_uop_ctrl_is_sta;
  reg  ldq_12_bits_uop_is_fence;
  reg  ldq_13_bits_uop_ctrl_is_load;
  reg  ldq_13_bits_uop_ctrl_is_sta;
  reg  ldq_13_bits_uop_is_fence;
  reg  ldq_14_bits_uop_ctrl_is_load;
  reg  ldq_14_bits_uop_ctrl_is_sta;
  reg  ldq_14_bits_uop_is_fence;
  reg  ldq_15_bits_uop_ctrl_is_load;
  reg  ldq_15_bits_uop_ctrl_is_sta;
  reg  ldq_15_bits_uop_is_fence;
  reg  ldq_16_bits_uop_ctrl_is_load;
  reg  ldq_16_bits_uop_ctrl_is_sta;
  reg  ldq_16_bits_uop_is_fence;
  reg  ldq_17_bits_uop_ctrl_is_load;
  reg  ldq_17_bits_uop_ctrl_is_sta;
  reg  ldq_17_bits_uop_is_fence;
  reg  ldq_18_bits_uop_ctrl_is_load;
  reg  ldq_18_bits_uop_ctrl_is_sta;
  reg  ldq_18_bits_uop_is_fence;
  reg  ldq_19_bits_uop_ctrl_is_load;
  reg  ldq_19_bits_uop_ctrl_is_sta;
  reg  ldq_19_bits_uop_is_fence;
  reg  ldq_20_bits_uop_ctrl_is_load;
  reg  ldq_20_bits_uop_ctrl_is_sta;
  reg  ldq_20_bits_uop_is_fence;
  reg  ldq_21_bits_uop_ctrl_is_load;
  reg  ldq_21_bits_uop_ctrl_is_sta;
  reg  ldq_21_bits_uop_is_fence;
  reg  ldq_22_bits_uop_ctrl_is_load;
  reg  ldq_22_bits_uop_ctrl_is_sta;
  reg  ldq_22_bits_uop_is_fence;
  reg  ldq_23_bits_uop_ctrl_is_load;
  reg  ldq_23_bits_uop_ctrl_is_sta;
  reg  ldq_23_bits_uop_is_fence;
  reg  ldq_24_bits_uop_ctrl_is_load;
  reg  ldq_24_bits_uop_ctrl_is_sta;
  reg  ldq_24_bits_uop_is_fence;
  reg  ldq_25_bits_uop_ctrl_is_load;
  reg  ldq_25_bits_uop_ctrl_is_sta;
  reg  ldq_25_bits_uop_is_fence;
  reg  ldq_26_bits_uop_ctrl_is_load;
  reg  ldq_26_bits_uop_ctrl_is_sta;
  reg  ldq_26_bits_uop_is_fence;
  reg  ldq_27_bits_uop_ctrl_is_load;
  reg  ldq_27_bits_uop_ctrl_is_sta;
  reg  ldq_27_bits_uop_is_fence;
  reg  ldq_28_bits_uop_ctrl_is_load;
  reg  ldq_28_bits_uop_ctrl_is_sta;
  reg  ldq_28_bits_uop_is_fence;
  reg  ldq_29_bits_uop_ctrl_is_load;
  reg  ldq_29_bits_uop_ctrl_is_sta;
  reg  ldq_29_bits_uop_is_fence;
  reg  ldq_30_bits_uop_ctrl_is_load;
  reg  ldq_30_bits_uop_ctrl_is_sta;
  reg  ldq_30_bits_uop_is_fence;
  reg  ldq_31_bits_uop_ctrl_is_load;
  reg  ldq_31_bits_uop_ctrl_is_sta;
  reg  ldq_31_bits_uop_is_fence;
  reg  stq_0_bits_uop_ctrl_is_load;
  reg  stq_0_bits_uop_ctrl_is_sta;
  reg  stq_1_bits_uop_ctrl_is_load;
  reg  stq_1_bits_uop_ctrl_is_sta;
  reg  stq_2_bits_uop_ctrl_is_load;
  reg  stq_2_bits_uop_ctrl_is_sta;
  reg  stq_3_bits_uop_ctrl_is_load;
  reg  stq_3_bits_uop_ctrl_is_sta;
  reg  stq_4_bits_uop_ctrl_is_load;
  reg  stq_4_bits_uop_ctrl_is_sta;
  reg  stq_5_bits_uop_ctrl_is_load;
  reg  stq_5_bits_uop_ctrl_is_sta;
  reg  stq_6_bits_uop_ctrl_is_load;
  reg  stq_6_bits_uop_ctrl_is_sta;
  reg  stq_7_bits_uop_ctrl_is_load;
  reg  stq_7_bits_uop_ctrl_is_sta;
  reg  stq_8_bits_uop_ctrl_is_load;
  reg  stq_8_bits_uop_ctrl_is_sta;
  reg  stq_9_bits_uop_ctrl_is_load;
  reg  stq_9_bits_uop_ctrl_is_sta;
  reg  stq_10_bits_uop_ctrl_is_load;
  reg  stq_10_bits_uop_ctrl_is_sta;
  reg  stq_11_bits_uop_ctrl_is_load;
  reg  stq_11_bits_uop_ctrl_is_sta;
  reg  stq_12_bits_uop_ctrl_is_load;
  reg  stq_12_bits_uop_ctrl_is_sta;
  reg  stq_13_bits_uop_ctrl_is_load;
  reg  stq_13_bits_uop_ctrl_is_sta;
  reg  stq_14_bits_uop_ctrl_is_load;
  reg  stq_14_bits_uop_ctrl_is_sta;
  reg  stq_15_bits_uop_ctrl_is_load;
  reg  stq_15_bits_uop_ctrl_is_sta;
  reg  stq_16_bits_uop_ctrl_is_load;
  reg  stq_16_bits_uop_ctrl_is_sta;
  reg  stq_17_bits_uop_ctrl_is_load;
  reg  stq_17_bits_uop_ctrl_is_sta;
  reg  stq_18_bits_uop_ctrl_is_load;
  reg  stq_18_bits_uop_ctrl_is_sta;
  reg  stq_19_bits_uop_ctrl_is_load;
  reg  stq_19_bits_uop_ctrl_is_sta;
  reg  stq_20_bits_uop_ctrl_is_load;
  reg  stq_20_bits_uop_ctrl_is_sta;
  reg  stq_21_bits_uop_ctrl_is_load;
  reg  stq_21_bits_uop_ctrl_is_sta;
  reg  stq_22_bits_uop_ctrl_is_load;
  reg  stq_22_bits_uop_ctrl_is_sta;
  reg  stq_23_bits_uop_ctrl_is_load;
  reg  stq_23_bits_uop_ctrl_is_sta;
  reg  stq_24_bits_uop_ctrl_is_load;
  reg  stq_24_bits_uop_ctrl_is_sta;
  reg  stq_25_bits_uop_ctrl_is_load;
  reg  stq_25_bits_uop_ctrl_is_sta;
  reg  stq_26_bits_uop_ctrl_is_load;
  reg  stq_26_bits_uop_ctrl_is_sta;
  reg  stq_27_bits_uop_ctrl_is_load;
  reg  stq_27_bits_uop_ctrl_is_sta;
  reg  stq_28_bits_uop_ctrl_is_load;
  reg  stq_28_bits_uop_ctrl_is_sta;
  reg  stq_29_bits_uop_ctrl_is_load;
  reg  stq_29_bits_uop_ctrl_is_sta;
  reg  stq_30_bits_uop_ctrl_is_load;
  reg  stq_30_bits_uop_ctrl_is_sta;
  reg  stq_31_bits_uop_ctrl_is_load;
  reg  stq_31_bits_uop_ctrl_is_sta;
  wire _GEN_301 = io_core_brupdate_b2_mispredict | _stq_stq_execute_head_valid_1 | stq_head == stq_execute_head | stq_tail == stq_execute_head;
  wire _GEN_302 = ldq_tail == io_core_dis_uops_0_bits_ldq_idx;
  always @(*) begin
    casez (ldq_tail)
      5'b00000:
        casez_tmp = ldq_0_valid;
      5'b00001:
        casez_tmp = ldq_1_valid;
      5'b00010:
        casez_tmp = ldq_2_valid;
      5'b00011:
        casez_tmp = ldq_3_valid;
      5'b00100:
        casez_tmp = ldq_4_valid;
      5'b00101:
        casez_tmp = ldq_5_valid;
      5'b00110:
        casez_tmp = ldq_6_valid;
      5'b00111:
        casez_tmp = ldq_7_valid;
      5'b01000:
        casez_tmp = ldq_8_valid;
      5'b01001:
        casez_tmp = ldq_9_valid;
      5'b01010:
        casez_tmp = ldq_10_valid;
      5'b01011:
        casez_tmp = ldq_11_valid;
      5'b01100:
        casez_tmp = ldq_12_valid;
      5'b01101:
        casez_tmp = ldq_13_valid;
      5'b01110:
        casez_tmp = ldq_14_valid;
      5'b01111:
        casez_tmp = ldq_15_valid;
      5'b10000:
        casez_tmp = ldq_16_valid;
      5'b10001:
        casez_tmp = ldq_17_valid;
      5'b10010:
        casez_tmp = ldq_18_valid;
      5'b10011:
        casez_tmp = ldq_19_valid;
      5'b10100:
        casez_tmp = ldq_20_valid;
      5'b10101:
        casez_tmp = ldq_21_valid;
      5'b10110:
        casez_tmp = ldq_22_valid;
      5'b10111:
        casez_tmp = ldq_23_valid;
      5'b11000:
        casez_tmp = ldq_24_valid;
      5'b11001:
        casez_tmp = ldq_25_valid;
      5'b11010:
        casez_tmp = ldq_26_valid;
      5'b11011:
        casez_tmp = ldq_27_valid;
      5'b11100:
        casez_tmp = ldq_28_valid;
      5'b11101:
        casez_tmp = ldq_29_valid;
      5'b11110:
        casez_tmp = ldq_30_valid;
      default:
        casez_tmp = ldq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_303 = stq_tail == io_core_dis_uops_0_bits_stq_idx;
  always @(*) begin
    casez (stq_tail)
      5'b00000:
        casez_tmp_0 = stq_0_valid;
      5'b00001:
        casez_tmp_0 = stq_1_valid;
      5'b00010:
        casez_tmp_0 = stq_2_valid;
      5'b00011:
        casez_tmp_0 = stq_3_valid;
      5'b00100:
        casez_tmp_0 = stq_4_valid;
      5'b00101:
        casez_tmp_0 = stq_5_valid;
      5'b00110:
        casez_tmp_0 = stq_6_valid;
      5'b00111:
        casez_tmp_0 = stq_7_valid;
      5'b01000:
        casez_tmp_0 = stq_8_valid;
      5'b01001:
        casez_tmp_0 = stq_9_valid;
      5'b01010:
        casez_tmp_0 = stq_10_valid;
      5'b01011:
        casez_tmp_0 = stq_11_valid;
      5'b01100:
        casez_tmp_0 = stq_12_valid;
      5'b01101:
        casez_tmp_0 = stq_13_valid;
      5'b01110:
        casez_tmp_0 = stq_14_valid;
      5'b01111:
        casez_tmp_0 = stq_15_valid;
      5'b10000:
        casez_tmp_0 = stq_16_valid;
      5'b10001:
        casez_tmp_0 = stq_17_valid;
      5'b10010:
        casez_tmp_0 = stq_18_valid;
      5'b10011:
        casez_tmp_0 = stq_19_valid;
      5'b10100:
        casez_tmp_0 = stq_20_valid;
      5'b10101:
        casez_tmp_0 = stq_21_valid;
      5'b10110:
        casez_tmp_0 = stq_22_valid;
      5'b10111:
        casez_tmp_0 = stq_23_valid;
      5'b11000:
        casez_tmp_0 = stq_24_valid;
      5'b11001:
        casez_tmp_0 = stq_25_valid;
      5'b11010:
        casez_tmp_0 = stq_26_valid;
      5'b11011:
        casez_tmp_0 = stq_27_valid;
      5'b11100:
        casez_tmp_0 = stq_28_valid;
      5'b11101:
        casez_tmp_0 = stq_29_valid;
      5'b11110:
        casez_tmp_0 = stq_30_valid;
      default:
        casez_tmp_0 = stq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_304 = dis_ld_val & dis_st_val;
  wire _GEN_305 = _GEN == io_core_dis_uops_1_bits_ldq_idx;
  always @(*) begin
    casez (_GEN)
      5'b00000:
        casez_tmp_1 = ldq_0_valid;
      5'b00001:
        casez_tmp_1 = ldq_1_valid;
      5'b00010:
        casez_tmp_1 = ldq_2_valid;
      5'b00011:
        casez_tmp_1 = ldq_3_valid;
      5'b00100:
        casez_tmp_1 = ldq_4_valid;
      5'b00101:
        casez_tmp_1 = ldq_5_valid;
      5'b00110:
        casez_tmp_1 = ldq_6_valid;
      5'b00111:
        casez_tmp_1 = ldq_7_valid;
      5'b01000:
        casez_tmp_1 = ldq_8_valid;
      5'b01001:
        casez_tmp_1 = ldq_9_valid;
      5'b01010:
        casez_tmp_1 = ldq_10_valid;
      5'b01011:
        casez_tmp_1 = ldq_11_valid;
      5'b01100:
        casez_tmp_1 = ldq_12_valid;
      5'b01101:
        casez_tmp_1 = ldq_13_valid;
      5'b01110:
        casez_tmp_1 = ldq_14_valid;
      5'b01111:
        casez_tmp_1 = ldq_15_valid;
      5'b10000:
        casez_tmp_1 = ldq_16_valid;
      5'b10001:
        casez_tmp_1 = ldq_17_valid;
      5'b10010:
        casez_tmp_1 = ldq_18_valid;
      5'b10011:
        casez_tmp_1 = ldq_19_valid;
      5'b10100:
        casez_tmp_1 = ldq_20_valid;
      5'b10101:
        casez_tmp_1 = ldq_21_valid;
      5'b10110:
        casez_tmp_1 = ldq_22_valid;
      5'b10111:
        casez_tmp_1 = ldq_23_valid;
      5'b11000:
        casez_tmp_1 = ldq_24_valid;
      5'b11001:
        casez_tmp_1 = ldq_25_valid;
      5'b11010:
        casez_tmp_1 = ldq_26_valid;
      5'b11011:
        casez_tmp_1 = ldq_27_valid;
      5'b11100:
        casez_tmp_1 = ldq_28_valid;
      5'b11101:
        casez_tmp_1 = ldq_29_valid;
      5'b11110:
        casez_tmp_1 = ldq_30_valid;
      default:
        casez_tmp_1 = ldq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_306 = _ldq_T_35_bits_youngest_stq_idx == io_core_dis_uops_1_bits_stq_idx;
  always @(*) begin
    casez (_ldq_T_35_bits_youngest_stq_idx)
      5'b00000:
        casez_tmp_2 = stq_0_valid;
      5'b00001:
        casez_tmp_2 = stq_1_valid;
      5'b00010:
        casez_tmp_2 = stq_2_valid;
      5'b00011:
        casez_tmp_2 = stq_3_valid;
      5'b00100:
        casez_tmp_2 = stq_4_valid;
      5'b00101:
        casez_tmp_2 = stq_5_valid;
      5'b00110:
        casez_tmp_2 = stq_6_valid;
      5'b00111:
        casez_tmp_2 = stq_7_valid;
      5'b01000:
        casez_tmp_2 = stq_8_valid;
      5'b01001:
        casez_tmp_2 = stq_9_valid;
      5'b01010:
        casez_tmp_2 = stq_10_valid;
      5'b01011:
        casez_tmp_2 = stq_11_valid;
      5'b01100:
        casez_tmp_2 = stq_12_valid;
      5'b01101:
        casez_tmp_2 = stq_13_valid;
      5'b01110:
        casez_tmp_2 = stq_14_valid;
      5'b01111:
        casez_tmp_2 = stq_15_valid;
      5'b10000:
        casez_tmp_2 = stq_16_valid;
      5'b10001:
        casez_tmp_2 = stq_17_valid;
      5'b10010:
        casez_tmp_2 = stq_18_valid;
      5'b10011:
        casez_tmp_2 = stq_19_valid;
      5'b10100:
        casez_tmp_2 = stq_20_valid;
      5'b10101:
        casez_tmp_2 = stq_21_valid;
      5'b10110:
        casez_tmp_2 = stq_22_valid;
      5'b10111:
        casez_tmp_2 = stq_23_valid;
      5'b11000:
        casez_tmp_2 = stq_24_valid;
      5'b11001:
        casez_tmp_2 = stq_25_valid;
      5'b11010:
        casez_tmp_2 = stq_26_valid;
      5'b11011:
        casez_tmp_2 = stq_27_valid;
      5'b11100:
        casez_tmp_2 = stq_28_valid;
      5'b11101:
        casez_tmp_2 = stq_29_valid;
      5'b11110:
        casez_tmp_2 = stq_30_valid;
      default:
        casez_tmp_2 = stq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_307 = dis_ld_val_1 & dis_st_val_1;
  wire _GEN_308 = _GEN_0 == io_core_dis_uops_2_bits_ldq_idx;
  always @(*) begin
    casez (_GEN_0)
      5'b00000:
        casez_tmp_3 = ldq_0_valid;
      5'b00001:
        casez_tmp_3 = ldq_1_valid;
      5'b00010:
        casez_tmp_3 = ldq_2_valid;
      5'b00011:
        casez_tmp_3 = ldq_3_valid;
      5'b00100:
        casez_tmp_3 = ldq_4_valid;
      5'b00101:
        casez_tmp_3 = ldq_5_valid;
      5'b00110:
        casez_tmp_3 = ldq_6_valid;
      5'b00111:
        casez_tmp_3 = ldq_7_valid;
      5'b01000:
        casez_tmp_3 = ldq_8_valid;
      5'b01001:
        casez_tmp_3 = ldq_9_valid;
      5'b01010:
        casez_tmp_3 = ldq_10_valid;
      5'b01011:
        casez_tmp_3 = ldq_11_valid;
      5'b01100:
        casez_tmp_3 = ldq_12_valid;
      5'b01101:
        casez_tmp_3 = ldq_13_valid;
      5'b01110:
        casez_tmp_3 = ldq_14_valid;
      5'b01111:
        casez_tmp_3 = ldq_15_valid;
      5'b10000:
        casez_tmp_3 = ldq_16_valid;
      5'b10001:
        casez_tmp_3 = ldq_17_valid;
      5'b10010:
        casez_tmp_3 = ldq_18_valid;
      5'b10011:
        casez_tmp_3 = ldq_19_valid;
      5'b10100:
        casez_tmp_3 = ldq_20_valid;
      5'b10101:
        casez_tmp_3 = ldq_21_valid;
      5'b10110:
        casez_tmp_3 = ldq_22_valid;
      5'b10111:
        casez_tmp_3 = ldq_23_valid;
      5'b11000:
        casez_tmp_3 = ldq_24_valid;
      5'b11001:
        casez_tmp_3 = ldq_25_valid;
      5'b11010:
        casez_tmp_3 = ldq_26_valid;
      5'b11011:
        casez_tmp_3 = ldq_27_valid;
      5'b11100:
        casez_tmp_3 = ldq_28_valid;
      5'b11101:
        casez_tmp_3 = ldq_29_valid;
      5'b11110:
        casez_tmp_3 = ldq_30_valid;
      default:
        casez_tmp_3 = ldq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_309 = _ldq_T_75_bits_youngest_stq_idx == io_core_dis_uops_2_bits_stq_idx;
  always @(*) begin
    casez (_ldq_T_75_bits_youngest_stq_idx)
      5'b00000:
        casez_tmp_4 = stq_0_valid;
      5'b00001:
        casez_tmp_4 = stq_1_valid;
      5'b00010:
        casez_tmp_4 = stq_2_valid;
      5'b00011:
        casez_tmp_4 = stq_3_valid;
      5'b00100:
        casez_tmp_4 = stq_4_valid;
      5'b00101:
        casez_tmp_4 = stq_5_valid;
      5'b00110:
        casez_tmp_4 = stq_6_valid;
      5'b00111:
        casez_tmp_4 = stq_7_valid;
      5'b01000:
        casez_tmp_4 = stq_8_valid;
      5'b01001:
        casez_tmp_4 = stq_9_valid;
      5'b01010:
        casez_tmp_4 = stq_10_valid;
      5'b01011:
        casez_tmp_4 = stq_11_valid;
      5'b01100:
        casez_tmp_4 = stq_12_valid;
      5'b01101:
        casez_tmp_4 = stq_13_valid;
      5'b01110:
        casez_tmp_4 = stq_14_valid;
      5'b01111:
        casez_tmp_4 = stq_15_valid;
      5'b10000:
        casez_tmp_4 = stq_16_valid;
      5'b10001:
        casez_tmp_4 = stq_17_valid;
      5'b10010:
        casez_tmp_4 = stq_18_valid;
      5'b10011:
        casez_tmp_4 = stq_19_valid;
      5'b10100:
        casez_tmp_4 = stq_20_valid;
      5'b10101:
        casez_tmp_4 = stq_21_valid;
      5'b10110:
        casez_tmp_4 = stq_22_valid;
      5'b10111:
        casez_tmp_4 = stq_23_valid;
      5'b11000:
        casez_tmp_4 = stq_24_valid;
      5'b11001:
        casez_tmp_4 = stq_25_valid;
      5'b11010:
        casez_tmp_4 = stq_26_valid;
      5'b11011:
        casez_tmp_4 = stq_27_valid;
      5'b11100:
        casez_tmp_4 = stq_28_valid;
      5'b11101:
        casez_tmp_4 = stq_29_valid;
      5'b11110:
        casez_tmp_4 = stq_30_valid;
      default:
        casez_tmp_4 = stq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_310 = dis_ld_val_2 & dis_st_val_2;
  wire _GEN_311 = _GEN_1 == io_core_dis_uops_3_bits_ldq_idx;
  always @(*) begin
    casez (_GEN_1)
      5'b00000:
        casez_tmp_5 = ldq_0_valid;
      5'b00001:
        casez_tmp_5 = ldq_1_valid;
      5'b00010:
        casez_tmp_5 = ldq_2_valid;
      5'b00011:
        casez_tmp_5 = ldq_3_valid;
      5'b00100:
        casez_tmp_5 = ldq_4_valid;
      5'b00101:
        casez_tmp_5 = ldq_5_valid;
      5'b00110:
        casez_tmp_5 = ldq_6_valid;
      5'b00111:
        casez_tmp_5 = ldq_7_valid;
      5'b01000:
        casez_tmp_5 = ldq_8_valid;
      5'b01001:
        casez_tmp_5 = ldq_9_valid;
      5'b01010:
        casez_tmp_5 = ldq_10_valid;
      5'b01011:
        casez_tmp_5 = ldq_11_valid;
      5'b01100:
        casez_tmp_5 = ldq_12_valid;
      5'b01101:
        casez_tmp_5 = ldq_13_valid;
      5'b01110:
        casez_tmp_5 = ldq_14_valid;
      5'b01111:
        casez_tmp_5 = ldq_15_valid;
      5'b10000:
        casez_tmp_5 = ldq_16_valid;
      5'b10001:
        casez_tmp_5 = ldq_17_valid;
      5'b10010:
        casez_tmp_5 = ldq_18_valid;
      5'b10011:
        casez_tmp_5 = ldq_19_valid;
      5'b10100:
        casez_tmp_5 = ldq_20_valid;
      5'b10101:
        casez_tmp_5 = ldq_21_valid;
      5'b10110:
        casez_tmp_5 = ldq_22_valid;
      5'b10111:
        casez_tmp_5 = ldq_23_valid;
      5'b11000:
        casez_tmp_5 = ldq_24_valid;
      5'b11001:
        casez_tmp_5 = ldq_25_valid;
      5'b11010:
        casez_tmp_5 = ldq_26_valid;
      5'b11011:
        casez_tmp_5 = ldq_27_valid;
      5'b11100:
        casez_tmp_5 = ldq_28_valid;
      5'b11101:
        casez_tmp_5 = ldq_29_valid;
      5'b11110:
        casez_tmp_5 = ldq_30_valid;
      default:
        casez_tmp_5 = ldq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_312 = _ldq_T_115_bits_youngest_stq_idx == io_core_dis_uops_3_bits_stq_idx;
  always @(*) begin
    casez (_ldq_T_115_bits_youngest_stq_idx)
      5'b00000:
        casez_tmp_6 = stq_0_valid;
      5'b00001:
        casez_tmp_6 = stq_1_valid;
      5'b00010:
        casez_tmp_6 = stq_2_valid;
      5'b00011:
        casez_tmp_6 = stq_3_valid;
      5'b00100:
        casez_tmp_6 = stq_4_valid;
      5'b00101:
        casez_tmp_6 = stq_5_valid;
      5'b00110:
        casez_tmp_6 = stq_6_valid;
      5'b00111:
        casez_tmp_6 = stq_7_valid;
      5'b01000:
        casez_tmp_6 = stq_8_valid;
      5'b01001:
        casez_tmp_6 = stq_9_valid;
      5'b01010:
        casez_tmp_6 = stq_10_valid;
      5'b01011:
        casez_tmp_6 = stq_11_valid;
      5'b01100:
        casez_tmp_6 = stq_12_valid;
      5'b01101:
        casez_tmp_6 = stq_13_valid;
      5'b01110:
        casez_tmp_6 = stq_14_valid;
      5'b01111:
        casez_tmp_6 = stq_15_valid;
      5'b10000:
        casez_tmp_6 = stq_16_valid;
      5'b10001:
        casez_tmp_6 = stq_17_valid;
      5'b10010:
        casez_tmp_6 = stq_18_valid;
      5'b10011:
        casez_tmp_6 = stq_19_valid;
      5'b10100:
        casez_tmp_6 = stq_20_valid;
      5'b10101:
        casez_tmp_6 = stq_21_valid;
      5'b10110:
        casez_tmp_6 = stq_22_valid;
      5'b10111:
        casez_tmp_6 = stq_23_valid;
      5'b11000:
        casez_tmp_6 = stq_24_valid;
      5'b11001:
        casez_tmp_6 = stq_25_valid;
      5'b11010:
        casez_tmp_6 = stq_26_valid;
      5'b11011:
        casez_tmp_6 = stq_27_valid;
      5'b11100:
        casez_tmp_6 = stq_28_valid;
      5'b11101:
        casez_tmp_6 = stq_29_valid;
      5'b11110:
        casez_tmp_6 = stq_30_valid;
      default:
        casez_tmp_6 = stq_31_valid;
    endcase
  end // always @(*)
  wire _GEN_313 = dis_ld_val_3 & dis_st_val_3;
  always @(*) begin
    casez (ldq_incoming_idx_0)
      5'b00000:
        casez_tmp_7 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_7 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_7 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_7 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_7 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_7 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_7 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_7 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_7 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_7 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_7 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_7 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_7 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_7 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_7 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_7 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_7 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_7 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_7 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_7 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_7 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_7 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_7 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_7 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_7 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_7 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_7 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_7 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_7 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_7 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_7 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_7 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_0)
      5'b00000:
        casez_tmp_8 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_8 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_8 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_8 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_8 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_8 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_8 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_8 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_8 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_8 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_8 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_8 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_8 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_8 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_8 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_8 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_8 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_8 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_8 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_8 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_8 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_8 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_8 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_8 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_8 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_8 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_8 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_8 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_8 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_8 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_8 = ldq_30_bits_executed;
      default:
        casez_tmp_8 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_1)
      5'b00000:
        casez_tmp_9 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_9 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_9 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_9 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_9 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_9 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_9 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_9 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_9 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_9 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_9 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_9 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_9 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_9 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_9 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_9 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_9 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_9 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_9 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_9 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_9 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_9 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_9 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_9 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_9 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_9 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_9 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_9 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_9 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_9 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_9 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_9 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_1)
      5'b00000:
        casez_tmp_10 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_10 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_10 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_10 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_10 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_10 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_10 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_10 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_10 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_10 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_10 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_10 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_10 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_10 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_10 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_10 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_10 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_10 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_10 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_10 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_10 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_10 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_10 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_10 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_10 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_10 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_10 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_10 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_10 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_10 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_10 = ldq_30_bits_executed;
      default:
        casez_tmp_10 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  wire _GEN_314 = _exe_cmd_T | will_fire_sta_incoming_0;
  wire _GEN_315 = exe_req_0_valid & ~(_GEN_314 | will_fire_std_incoming_0 | will_fire_sfence_0);
  wire _GEN_316 = _exe_cmd_T_7 | will_fire_sta_incoming_1;
  wire _GEN_317 = exe_req_1_valid & ~(_GEN_316 | will_fire_std_incoming_1 | will_fire_sfence_1);
  wire _GEN_318 = (will_fire_sfence_0 | will_fire_sfence_1) & ~(will_fire_sfence_0 & will_fire_sfence_1);
  wire _GEN_319 = _GEN_2 & hella_req_cmd == 5'h14;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_11 = stq_0_bits_uop_ctrl_is_load;
      5'b00001:
        casez_tmp_11 = stq_1_bits_uop_ctrl_is_load;
      5'b00010:
        casez_tmp_11 = stq_2_bits_uop_ctrl_is_load;
      5'b00011:
        casez_tmp_11 = stq_3_bits_uop_ctrl_is_load;
      5'b00100:
        casez_tmp_11 = stq_4_bits_uop_ctrl_is_load;
      5'b00101:
        casez_tmp_11 = stq_5_bits_uop_ctrl_is_load;
      5'b00110:
        casez_tmp_11 = stq_6_bits_uop_ctrl_is_load;
      5'b00111:
        casez_tmp_11 = stq_7_bits_uop_ctrl_is_load;
      5'b01000:
        casez_tmp_11 = stq_8_bits_uop_ctrl_is_load;
      5'b01001:
        casez_tmp_11 = stq_9_bits_uop_ctrl_is_load;
      5'b01010:
        casez_tmp_11 = stq_10_bits_uop_ctrl_is_load;
      5'b01011:
        casez_tmp_11 = stq_11_bits_uop_ctrl_is_load;
      5'b01100:
        casez_tmp_11 = stq_12_bits_uop_ctrl_is_load;
      5'b01101:
        casez_tmp_11 = stq_13_bits_uop_ctrl_is_load;
      5'b01110:
        casez_tmp_11 = stq_14_bits_uop_ctrl_is_load;
      5'b01111:
        casez_tmp_11 = stq_15_bits_uop_ctrl_is_load;
      5'b10000:
        casez_tmp_11 = stq_16_bits_uop_ctrl_is_load;
      5'b10001:
        casez_tmp_11 = stq_17_bits_uop_ctrl_is_load;
      5'b10010:
        casez_tmp_11 = stq_18_bits_uop_ctrl_is_load;
      5'b10011:
        casez_tmp_11 = stq_19_bits_uop_ctrl_is_load;
      5'b10100:
        casez_tmp_11 = stq_20_bits_uop_ctrl_is_load;
      5'b10101:
        casez_tmp_11 = stq_21_bits_uop_ctrl_is_load;
      5'b10110:
        casez_tmp_11 = stq_22_bits_uop_ctrl_is_load;
      5'b10111:
        casez_tmp_11 = stq_23_bits_uop_ctrl_is_load;
      5'b11000:
        casez_tmp_11 = stq_24_bits_uop_ctrl_is_load;
      5'b11001:
        casez_tmp_11 = stq_25_bits_uop_ctrl_is_load;
      5'b11010:
        casez_tmp_11 = stq_26_bits_uop_ctrl_is_load;
      5'b11011:
        casez_tmp_11 = stq_27_bits_uop_ctrl_is_load;
      5'b11100:
        casez_tmp_11 = stq_28_bits_uop_ctrl_is_load;
      5'b11101:
        casez_tmp_11 = stq_29_bits_uop_ctrl_is_load;
      5'b11110:
        casez_tmp_11 = stq_30_bits_uop_ctrl_is_load;
      default:
        casez_tmp_11 = stq_31_bits_uop_ctrl_is_load;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_12 = stq_0_bits_uop_ctrl_is_sta;
      5'b00001:
        casez_tmp_12 = stq_1_bits_uop_ctrl_is_sta;
      5'b00010:
        casez_tmp_12 = stq_2_bits_uop_ctrl_is_sta;
      5'b00011:
        casez_tmp_12 = stq_3_bits_uop_ctrl_is_sta;
      5'b00100:
        casez_tmp_12 = stq_4_bits_uop_ctrl_is_sta;
      5'b00101:
        casez_tmp_12 = stq_5_bits_uop_ctrl_is_sta;
      5'b00110:
        casez_tmp_12 = stq_6_bits_uop_ctrl_is_sta;
      5'b00111:
        casez_tmp_12 = stq_7_bits_uop_ctrl_is_sta;
      5'b01000:
        casez_tmp_12 = stq_8_bits_uop_ctrl_is_sta;
      5'b01001:
        casez_tmp_12 = stq_9_bits_uop_ctrl_is_sta;
      5'b01010:
        casez_tmp_12 = stq_10_bits_uop_ctrl_is_sta;
      5'b01011:
        casez_tmp_12 = stq_11_bits_uop_ctrl_is_sta;
      5'b01100:
        casez_tmp_12 = stq_12_bits_uop_ctrl_is_sta;
      5'b01101:
        casez_tmp_12 = stq_13_bits_uop_ctrl_is_sta;
      5'b01110:
        casez_tmp_12 = stq_14_bits_uop_ctrl_is_sta;
      5'b01111:
        casez_tmp_12 = stq_15_bits_uop_ctrl_is_sta;
      5'b10000:
        casez_tmp_12 = stq_16_bits_uop_ctrl_is_sta;
      5'b10001:
        casez_tmp_12 = stq_17_bits_uop_ctrl_is_sta;
      5'b10010:
        casez_tmp_12 = stq_18_bits_uop_ctrl_is_sta;
      5'b10011:
        casez_tmp_12 = stq_19_bits_uop_ctrl_is_sta;
      5'b10100:
        casez_tmp_12 = stq_20_bits_uop_ctrl_is_sta;
      5'b10101:
        casez_tmp_12 = stq_21_bits_uop_ctrl_is_sta;
      5'b10110:
        casez_tmp_12 = stq_22_bits_uop_ctrl_is_sta;
      5'b10111:
        casez_tmp_12 = stq_23_bits_uop_ctrl_is_sta;
      5'b11000:
        casez_tmp_12 = stq_24_bits_uop_ctrl_is_sta;
      5'b11001:
        casez_tmp_12 = stq_25_bits_uop_ctrl_is_sta;
      5'b11010:
        casez_tmp_12 = stq_26_bits_uop_ctrl_is_sta;
      5'b11011:
        casez_tmp_12 = stq_27_bits_uop_ctrl_is_sta;
      5'b11100:
        casez_tmp_12 = stq_28_bits_uop_ctrl_is_sta;
      5'b11101:
        casez_tmp_12 = stq_29_bits_uop_ctrl_is_sta;
      5'b11110:
        casez_tmp_12 = stq_30_bits_uop_ctrl_is_sta;
      default:
        casez_tmp_12 = stq_31_bits_uop_ctrl_is_sta;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_13 = stq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_13 = stq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_13 = stq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_13 = stq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_13 = stq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_13 = stq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_13 = stq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_13 = stq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_13 = stq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_13 = stq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_13 = stq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_13 = stq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_13 = stq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_13 = stq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_13 = stq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_13 = stq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_13 = stq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_13 = stq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_13 = stq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_13 = stq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_13 = stq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_13 = stq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_13 = stq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_13 = stq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_13 = stq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_13 = stq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_13 = stq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_13 = stq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_13 = stq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_13 = stq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_13 = stq_30_bits_uop_is_fence;
      default:
        casez_tmp_13 = stq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_14 = ldq_0_bits_uop_ctrl_is_load;
      5'b00001:
        casez_tmp_14 = ldq_1_bits_uop_ctrl_is_load;
      5'b00010:
        casez_tmp_14 = ldq_2_bits_uop_ctrl_is_load;
      5'b00011:
        casez_tmp_14 = ldq_3_bits_uop_ctrl_is_load;
      5'b00100:
        casez_tmp_14 = ldq_4_bits_uop_ctrl_is_load;
      5'b00101:
        casez_tmp_14 = ldq_5_bits_uop_ctrl_is_load;
      5'b00110:
        casez_tmp_14 = ldq_6_bits_uop_ctrl_is_load;
      5'b00111:
        casez_tmp_14 = ldq_7_bits_uop_ctrl_is_load;
      5'b01000:
        casez_tmp_14 = ldq_8_bits_uop_ctrl_is_load;
      5'b01001:
        casez_tmp_14 = ldq_9_bits_uop_ctrl_is_load;
      5'b01010:
        casez_tmp_14 = ldq_10_bits_uop_ctrl_is_load;
      5'b01011:
        casez_tmp_14 = ldq_11_bits_uop_ctrl_is_load;
      5'b01100:
        casez_tmp_14 = ldq_12_bits_uop_ctrl_is_load;
      5'b01101:
        casez_tmp_14 = ldq_13_bits_uop_ctrl_is_load;
      5'b01110:
        casez_tmp_14 = ldq_14_bits_uop_ctrl_is_load;
      5'b01111:
        casez_tmp_14 = ldq_15_bits_uop_ctrl_is_load;
      5'b10000:
        casez_tmp_14 = ldq_16_bits_uop_ctrl_is_load;
      5'b10001:
        casez_tmp_14 = ldq_17_bits_uop_ctrl_is_load;
      5'b10010:
        casez_tmp_14 = ldq_18_bits_uop_ctrl_is_load;
      5'b10011:
        casez_tmp_14 = ldq_19_bits_uop_ctrl_is_load;
      5'b10100:
        casez_tmp_14 = ldq_20_bits_uop_ctrl_is_load;
      5'b10101:
        casez_tmp_14 = ldq_21_bits_uop_ctrl_is_load;
      5'b10110:
        casez_tmp_14 = ldq_22_bits_uop_ctrl_is_load;
      5'b10111:
        casez_tmp_14 = ldq_23_bits_uop_ctrl_is_load;
      5'b11000:
        casez_tmp_14 = ldq_24_bits_uop_ctrl_is_load;
      5'b11001:
        casez_tmp_14 = ldq_25_bits_uop_ctrl_is_load;
      5'b11010:
        casez_tmp_14 = ldq_26_bits_uop_ctrl_is_load;
      5'b11011:
        casez_tmp_14 = ldq_27_bits_uop_ctrl_is_load;
      5'b11100:
        casez_tmp_14 = ldq_28_bits_uop_ctrl_is_load;
      5'b11101:
        casez_tmp_14 = ldq_29_bits_uop_ctrl_is_load;
      5'b11110:
        casez_tmp_14 = ldq_30_bits_uop_ctrl_is_load;
      default:
        casez_tmp_14 = ldq_31_bits_uop_ctrl_is_load;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_15 = ldq_0_bits_uop_ctrl_is_sta;
      5'b00001:
        casez_tmp_15 = ldq_1_bits_uop_ctrl_is_sta;
      5'b00010:
        casez_tmp_15 = ldq_2_bits_uop_ctrl_is_sta;
      5'b00011:
        casez_tmp_15 = ldq_3_bits_uop_ctrl_is_sta;
      5'b00100:
        casez_tmp_15 = ldq_4_bits_uop_ctrl_is_sta;
      5'b00101:
        casez_tmp_15 = ldq_5_bits_uop_ctrl_is_sta;
      5'b00110:
        casez_tmp_15 = ldq_6_bits_uop_ctrl_is_sta;
      5'b00111:
        casez_tmp_15 = ldq_7_bits_uop_ctrl_is_sta;
      5'b01000:
        casez_tmp_15 = ldq_8_bits_uop_ctrl_is_sta;
      5'b01001:
        casez_tmp_15 = ldq_9_bits_uop_ctrl_is_sta;
      5'b01010:
        casez_tmp_15 = ldq_10_bits_uop_ctrl_is_sta;
      5'b01011:
        casez_tmp_15 = ldq_11_bits_uop_ctrl_is_sta;
      5'b01100:
        casez_tmp_15 = ldq_12_bits_uop_ctrl_is_sta;
      5'b01101:
        casez_tmp_15 = ldq_13_bits_uop_ctrl_is_sta;
      5'b01110:
        casez_tmp_15 = ldq_14_bits_uop_ctrl_is_sta;
      5'b01111:
        casez_tmp_15 = ldq_15_bits_uop_ctrl_is_sta;
      5'b10000:
        casez_tmp_15 = ldq_16_bits_uop_ctrl_is_sta;
      5'b10001:
        casez_tmp_15 = ldq_17_bits_uop_ctrl_is_sta;
      5'b10010:
        casez_tmp_15 = ldq_18_bits_uop_ctrl_is_sta;
      5'b10011:
        casez_tmp_15 = ldq_19_bits_uop_ctrl_is_sta;
      5'b10100:
        casez_tmp_15 = ldq_20_bits_uop_ctrl_is_sta;
      5'b10101:
        casez_tmp_15 = ldq_21_bits_uop_ctrl_is_sta;
      5'b10110:
        casez_tmp_15 = ldq_22_bits_uop_ctrl_is_sta;
      5'b10111:
        casez_tmp_15 = ldq_23_bits_uop_ctrl_is_sta;
      5'b11000:
        casez_tmp_15 = ldq_24_bits_uop_ctrl_is_sta;
      5'b11001:
        casez_tmp_15 = ldq_25_bits_uop_ctrl_is_sta;
      5'b11010:
        casez_tmp_15 = ldq_26_bits_uop_ctrl_is_sta;
      5'b11011:
        casez_tmp_15 = ldq_27_bits_uop_ctrl_is_sta;
      5'b11100:
        casez_tmp_15 = ldq_28_bits_uop_ctrl_is_sta;
      5'b11101:
        casez_tmp_15 = ldq_29_bits_uop_ctrl_is_sta;
      5'b11110:
        casez_tmp_15 = ldq_30_bits_uop_ctrl_is_sta;
      default:
        casez_tmp_15 = ldq_31_bits_uop_ctrl_is_sta;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_16 = ldq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_16 = ldq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_16 = ldq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_16 = ldq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_16 = ldq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_16 = ldq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_16 = ldq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_16 = ldq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_16 = ldq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_16 = ldq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_16 = ldq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_16 = ldq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_16 = ldq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_16 = ldq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_16 = ldq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_16 = ldq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_16 = ldq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_16 = ldq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_16 = ldq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_16 = ldq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_16 = ldq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_16 = ldq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_16 = ldq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_16 = ldq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_16 = ldq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_16 = ldq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_16 = ldq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_16 = ldq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_16 = ldq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_16 = ldq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_16 = ldq_30_bits_uop_is_fence;
      default:
        casez_tmp_16 = ldq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  reg  mem_xcpt_uops_0_uses_stq;
  reg  mem_xcpt_uops_1_uses_stq;
  wire _GEN_320 = exe_tlb_valid_0 & _exe_tlb_uop_T_2 & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_fence : io_core_exe_0_req_bits_uop_is_fence);
  wire _GEN_321 = (can_fire_load_incoming_0 | will_fire_sta_incoming_0 | will_fire_stad_incoming_0) & exe_req_0_bits_mxcpt_valid & exe_tlb_valid_0 & ~(_exe_tlb_uop_T_2 & mem_incoming_uop_out_ctrl_is_load | _exe_tlb_uop_T_2 & mem_incoming_uop_out_ctrl_is_sta);
  wire _GEN_322 = exe_tlb_valid_1 & (_exe_tlb_uop_T_9 ? (io_core_exe_1_req_bits_sfence_valid | ~io_core_exe_0_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_fence : io_core_exe_0_req_bits_uop_is_fence) : will_fire_load_retry_1 ? casez_tmp_16 : will_fire_sta_retry_1 & casez_tmp_13);
  wire _GEN_323 = (can_fire_load_incoming_1 | will_fire_sta_incoming_1 | will_fire_stad_incoming_1) & exe_req_1_bits_mxcpt_valid & exe_tlb_valid_1 & ~((_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_ctrl_is_load : will_fire_load_retry_1 ? casez_tmp_14 : will_fire_sta_retry_1 & casez_tmp_11) | (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_ctrl_is_sta : will_fire_load_retry_1 ? casez_tmp_15 : will_fire_sta_retry_1 & casez_tmp_12));
  wire _GEN_324 = exe_tlb_paddr_0 == dtlb_io_resp_0_paddr | exe_req_0_bits_sfence_valid;
  reg  REG;
  wire _GEN_325 = mem_xcpt_uops_0_uses_ldq ^ mem_xcpt_uops_0_uses_stq;
  wire _GEN_326 = exe_tlb_paddr_1 == dtlb_io_resp_1_paddr | exe_req_1_bits_sfence_valid;
  reg  REG_1;
  wire _GEN_327 = mem_xcpt_uops_1_uses_ldq ^ mem_xcpt_uops_1_uses_stq;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_17 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_17 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_17 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_17 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_17 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_17 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_17 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_17 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_17 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_17 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_17 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_17 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_17 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_17 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_17 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_17 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_17 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_17 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_17 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_17 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_17 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_17 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_17 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_17 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_17 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_17 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_17 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_17 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_17 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_17 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_17 = ldq_30_bits_executed;
      default:
        casez_tmp_17 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  wire _GEN_328 = can_fire_load_incoming_0 & casez_tmp_7;
  wire _GEN_329 = will_fire_sta_incoming_0 & stq_incoming_e_0_bits_addr_valid;
  always @(*) begin
    casez (sidx)
      5'b00000:
        casez_tmp_18 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_18 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_18 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_18 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_18 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_18 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_18 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_18 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_18 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_18 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_18 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_18 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_18 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_18 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_18 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_18 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_18 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_18 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_18 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_18 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_18 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_18 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_18 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_18 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_18 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_18 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_18 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_18 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_18 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_18 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_18 = stq_30_bits_data_valid;
      default:
        casez_tmp_18 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  wire _GEN_330 = ~mem_ldq_wakeup_e_out_bits_executed & ~mem_ldq_wakeup_e_out_bits_addr_is_virtual;
  wire _GEN_331 = can_fire_load_incoming_1 & casez_tmp_9;
  wire _GEN_332 = will_fire_sta_incoming_1 & stq_incoming_e_1_bits_addr_valid;
  always @(*) begin
    casez (sidx_1)
      5'b00000:
        casez_tmp_19 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_19 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_19 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_19 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_19 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_19 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_19 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_19 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_19 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_19 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_19 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_19 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_19 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_19 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_19 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_19 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_19 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_19 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_19 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_19 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_19 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_19 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_19 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_19 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_19 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_19 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_19 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_19 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_19 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_19 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_19 = stq_30_bits_data_valid;
      default:
        casez_tmp_19 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  wire _GEN_333 = _GEN_260 | _GEN_261;
  always @(*) begin
    casez (io_dmem_nack_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_20 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_20 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_20 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_20 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_20 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_20 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_20 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_20 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_20 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_20 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_20 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_20 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_20 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_20 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_20 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_20 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_20 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_20 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_20 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_20 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_20 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_20 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_20 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_20 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_20 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_20 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_20 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_20 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_20 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_20 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_20 = ldq_30_bits_executed;
      default:
        casez_tmp_20 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  wire _GEN_334 = send_iresp ^ send_fresp;
  always @(*) begin
    casez (io_dmem_nack_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_21 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_21 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_21 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_21 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_21 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_21 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_21 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_21 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_21 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_21 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_21 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_21 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_21 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_21 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_21 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_21 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_21 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_21 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_21 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_21 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_21 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_21 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_21 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_21 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_21 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_21 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_21 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_21 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_21 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_21 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_21 = ldq_30_bits_executed;
      default:
        casez_tmp_21 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  wire _GEN_335 = send_iresp_1 ^ send_fresp_1;
  wire _GEN_336 = (|_GEN_262) & stq_0_valid & stq_0_bits_committed;
  wire _GEN_337 = (|_GEN_263) & stq_1_valid & stq_1_bits_committed;
  wire _GEN_338 = (|_GEN_264) & stq_2_valid & stq_2_bits_committed;
  wire _GEN_339 = (|_GEN_265) & stq_3_valid & stq_3_bits_committed;
  wire _GEN_340 = (|_GEN_266) & stq_4_valid & stq_4_bits_committed;
  wire _GEN_341 = (|_GEN_267) & stq_5_valid & stq_5_bits_committed;
  wire _GEN_342 = (|_GEN_268) & stq_6_valid & stq_6_bits_committed;
  wire _GEN_343 = (|_GEN_269) & stq_7_valid & stq_7_bits_committed;
  wire _GEN_344 = (|_GEN_270) & stq_8_valid & stq_8_bits_committed;
  wire _GEN_345 = (|_GEN_271) & stq_9_valid & stq_9_bits_committed;
  wire _GEN_346 = (|_GEN_272) & stq_10_valid & stq_10_bits_committed;
  wire _GEN_347 = (|_GEN_273) & stq_11_valid & stq_11_bits_committed;
  wire _GEN_348 = (|_GEN_274) & stq_12_valid & stq_12_bits_committed;
  wire _GEN_349 = (|_GEN_275) & stq_13_valid & stq_13_bits_committed;
  wire _GEN_350 = (|_GEN_276) & stq_14_valid & stq_14_bits_committed;
  wire _GEN_351 = (|_GEN_277) & stq_15_valid & stq_15_bits_committed;
  wire _GEN_352 = (|_GEN_278) & stq_16_valid & stq_16_bits_committed;
  wire _GEN_353 = (|_GEN_279) & stq_17_valid & stq_17_bits_committed;
  wire _GEN_354 = (|_GEN_280) & stq_18_valid & stq_18_bits_committed;
  wire _GEN_355 = (|_GEN_281) & stq_19_valid & stq_19_bits_committed;
  wire _GEN_356 = (|_GEN_282) & stq_20_valid & stq_20_bits_committed;
  wire _GEN_357 = (|_GEN_283) & stq_21_valid & stq_21_bits_committed;
  wire _GEN_358 = (|_GEN_284) & stq_22_valid & stq_22_bits_committed;
  wire _GEN_359 = (|_GEN_285) & stq_23_valid & stq_23_bits_committed;
  wire _GEN_360 = (|_GEN_286) & stq_24_valid & stq_24_bits_committed;
  wire _GEN_361 = (|_GEN_287) & stq_25_valid & stq_25_bits_committed;
  wire _GEN_362 = (|_GEN_288) & stq_26_valid & stq_26_bits_committed;
  wire _GEN_363 = (|_GEN_289) & stq_27_valid & stq_27_bits_committed;
  wire _GEN_364 = (|_GEN_290) & stq_28_valid & stq_28_bits_committed;
  wire _GEN_365 = (|_GEN_291) & stq_29_valid & stq_29_bits_committed;
  wire _GEN_366 = (|_GEN_292) & stq_30_valid & stq_30_bits_committed;
  wire _GEN_367 = (|_GEN_293) & stq_31_valid & stq_31_bits_committed;
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_22 = ldq_0_valid;
      5'b00001:
        casez_tmp_22 = ldq_1_valid;
      5'b00010:
        casez_tmp_22 = ldq_2_valid;
      5'b00011:
        casez_tmp_22 = ldq_3_valid;
      5'b00100:
        casez_tmp_22 = ldq_4_valid;
      5'b00101:
        casez_tmp_22 = ldq_5_valid;
      5'b00110:
        casez_tmp_22 = ldq_6_valid;
      5'b00111:
        casez_tmp_22 = ldq_7_valid;
      5'b01000:
        casez_tmp_22 = ldq_8_valid;
      5'b01001:
        casez_tmp_22 = ldq_9_valid;
      5'b01010:
        casez_tmp_22 = ldq_10_valid;
      5'b01011:
        casez_tmp_22 = ldq_11_valid;
      5'b01100:
        casez_tmp_22 = ldq_12_valid;
      5'b01101:
        casez_tmp_22 = ldq_13_valid;
      5'b01110:
        casez_tmp_22 = ldq_14_valid;
      5'b01111:
        casez_tmp_22 = ldq_15_valid;
      5'b10000:
        casez_tmp_22 = ldq_16_valid;
      5'b10001:
        casez_tmp_22 = ldq_17_valid;
      5'b10010:
        casez_tmp_22 = ldq_18_valid;
      5'b10011:
        casez_tmp_22 = ldq_19_valid;
      5'b10100:
        casez_tmp_22 = ldq_20_valid;
      5'b10101:
        casez_tmp_22 = ldq_21_valid;
      5'b10110:
        casez_tmp_22 = ldq_22_valid;
      5'b10111:
        casez_tmp_22 = ldq_23_valid;
      5'b11000:
        casez_tmp_22 = ldq_24_valid;
      5'b11001:
        casez_tmp_22 = ldq_25_valid;
      5'b11010:
        casez_tmp_22 = ldq_26_valid;
      5'b11011:
        casez_tmp_22 = ldq_27_valid;
      5'b11100:
        casez_tmp_22 = ldq_28_valid;
      5'b11101:
        casez_tmp_22 = ldq_29_valid;
      5'b11110:
        casez_tmp_22 = ldq_30_valid;
      default:
        casez_tmp_22 = ldq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_23 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_23 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_23 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_23 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_23 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_23 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_23 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_23 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_23 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_23 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_23 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_23 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_23 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_23 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_23 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_23 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_23 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_23 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_23 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_23 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_23 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_23 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_23 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_23 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_23 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_23 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_23 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_23 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_23 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_23 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_23 = ldq_30_bits_executed;
      default:
        casez_tmp_23 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_24 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_24 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_24 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_24 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_24 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_24 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_24 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_24 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_24 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_24 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_24 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_24 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_24 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_24 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_24 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_24 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_24 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_24 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_24 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_24 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_24 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_24 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_24 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_24 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_24 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_24 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_24 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_24 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_24 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_24 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_24 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_24 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx)
      5'b00000:
        casez_tmp_25 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_25 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_25 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_25 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_25 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_25 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_25 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_25 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_25 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_25 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_25 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_25 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_25 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_25 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_25 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_25 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_25 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_25 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_25 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_25 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_25 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_25 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_25 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_25 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_25 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_25 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_25 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_25 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_25 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_25 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_25 = ldq_30_bits_succeeded;
      default:
        casez_tmp_25 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  wire _GEN_368 = (casez_tmp_23 | casez_tmp_24) & casez_tmp_25;
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_26 = ldq_0_valid;
      5'b00001:
        casez_tmp_26 = ldq_1_valid;
      5'b00010:
        casez_tmp_26 = ldq_2_valid;
      5'b00011:
        casez_tmp_26 = ldq_3_valid;
      5'b00100:
        casez_tmp_26 = ldq_4_valid;
      5'b00101:
        casez_tmp_26 = ldq_5_valid;
      5'b00110:
        casez_tmp_26 = ldq_6_valid;
      5'b00111:
        casez_tmp_26 = ldq_7_valid;
      5'b01000:
        casez_tmp_26 = ldq_8_valid;
      5'b01001:
        casez_tmp_26 = ldq_9_valid;
      5'b01010:
        casez_tmp_26 = ldq_10_valid;
      5'b01011:
        casez_tmp_26 = ldq_11_valid;
      5'b01100:
        casez_tmp_26 = ldq_12_valid;
      5'b01101:
        casez_tmp_26 = ldq_13_valid;
      5'b01110:
        casez_tmp_26 = ldq_14_valid;
      5'b01111:
        casez_tmp_26 = ldq_15_valid;
      5'b10000:
        casez_tmp_26 = ldq_16_valid;
      5'b10001:
        casez_tmp_26 = ldq_17_valid;
      5'b10010:
        casez_tmp_26 = ldq_18_valid;
      5'b10011:
        casez_tmp_26 = ldq_19_valid;
      5'b10100:
        casez_tmp_26 = ldq_20_valid;
      5'b10101:
        casez_tmp_26 = ldq_21_valid;
      5'b10110:
        casez_tmp_26 = ldq_22_valid;
      5'b10111:
        casez_tmp_26 = ldq_23_valid;
      5'b11000:
        casez_tmp_26 = ldq_24_valid;
      5'b11001:
        casez_tmp_26 = ldq_25_valid;
      5'b11010:
        casez_tmp_26 = ldq_26_valid;
      5'b11011:
        casez_tmp_26 = ldq_27_valid;
      5'b11100:
        casez_tmp_26 = ldq_28_valid;
      5'b11101:
        casez_tmp_26 = ldq_29_valid;
      5'b11110:
        casez_tmp_26 = ldq_30_valid;
      default:
        casez_tmp_26 = ldq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_27 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_27 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_27 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_27 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_27 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_27 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_27 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_27 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_27 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_27 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_27 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_27 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_27 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_27 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_27 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_27 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_27 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_27 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_27 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_27 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_27 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_27 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_27 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_27 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_27 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_27 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_27 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_27 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_27 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_27 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_27 = ldq_30_bits_executed;
      default:
        casez_tmp_27 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_28 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_28 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_28 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_28 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_28 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_28 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_28 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_28 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_28 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_28 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_28 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_28 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_28 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_28 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_28 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_28 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_28 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_28 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_28 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_28 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_28 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_28 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_28 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_28 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_28 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_28 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_28 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_28 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_28 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_28 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_28 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_28 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_1)
      5'b00000:
        casez_tmp_29 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_29 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_29 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_29 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_29 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_29 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_29 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_29 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_29 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_29 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_29 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_29 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_29 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_29 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_29 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_29 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_29 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_29 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_29 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_29 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_29 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_29 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_29 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_29 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_29 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_29 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_29 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_29 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_29 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_29 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_29 = ldq_30_bits_succeeded;
      default:
        casez_tmp_29 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  wire _GEN_369 = (casez_tmp_27 | casez_tmp_28) & casez_tmp_29;
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_30 = ldq_0_valid;
      5'b00001:
        casez_tmp_30 = ldq_1_valid;
      5'b00010:
        casez_tmp_30 = ldq_2_valid;
      5'b00011:
        casez_tmp_30 = ldq_3_valid;
      5'b00100:
        casez_tmp_30 = ldq_4_valid;
      5'b00101:
        casez_tmp_30 = ldq_5_valid;
      5'b00110:
        casez_tmp_30 = ldq_6_valid;
      5'b00111:
        casez_tmp_30 = ldq_7_valid;
      5'b01000:
        casez_tmp_30 = ldq_8_valid;
      5'b01001:
        casez_tmp_30 = ldq_9_valid;
      5'b01010:
        casez_tmp_30 = ldq_10_valid;
      5'b01011:
        casez_tmp_30 = ldq_11_valid;
      5'b01100:
        casez_tmp_30 = ldq_12_valid;
      5'b01101:
        casez_tmp_30 = ldq_13_valid;
      5'b01110:
        casez_tmp_30 = ldq_14_valid;
      5'b01111:
        casez_tmp_30 = ldq_15_valid;
      5'b10000:
        casez_tmp_30 = ldq_16_valid;
      5'b10001:
        casez_tmp_30 = ldq_17_valid;
      5'b10010:
        casez_tmp_30 = ldq_18_valid;
      5'b10011:
        casez_tmp_30 = ldq_19_valid;
      5'b10100:
        casez_tmp_30 = ldq_20_valid;
      5'b10101:
        casez_tmp_30 = ldq_21_valid;
      5'b10110:
        casez_tmp_30 = ldq_22_valid;
      5'b10111:
        casez_tmp_30 = ldq_23_valid;
      5'b11000:
        casez_tmp_30 = ldq_24_valid;
      5'b11001:
        casez_tmp_30 = ldq_25_valid;
      5'b11010:
        casez_tmp_30 = ldq_26_valid;
      5'b11011:
        casez_tmp_30 = ldq_27_valid;
      5'b11100:
        casez_tmp_30 = ldq_28_valid;
      5'b11101:
        casez_tmp_30 = ldq_29_valid;
      5'b11110:
        casez_tmp_30 = ldq_30_valid;
      default:
        casez_tmp_30 = ldq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_31 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_31 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_31 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_31 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_31 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_31 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_31 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_31 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_31 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_31 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_31 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_31 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_31 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_31 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_31 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_31 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_31 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_31 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_31 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_31 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_31 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_31 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_31 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_31 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_31 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_31 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_31 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_31 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_31 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_31 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_31 = ldq_30_bits_executed;
      default:
        casez_tmp_31 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_32 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_32 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_32 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_32 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_32 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_32 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_32 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_32 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_32 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_32 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_32 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_32 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_32 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_32 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_32 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_32 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_32 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_32 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_32 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_32 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_32 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_32 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_32 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_32 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_32 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_32 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_32 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_32 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_32 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_32 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_32 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_32 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_2)
      5'b00000:
        casez_tmp_33 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_33 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_33 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_33 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_33 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_33 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_33 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_33 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_33 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_33 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_33 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_33 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_33 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_33 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_33 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_33 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_33 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_33 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_33 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_33 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_33 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_33 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_33 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_33 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_33 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_33 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_33 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_33 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_33 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_33 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_33 = ldq_30_bits_succeeded;
      default:
        casez_tmp_33 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  wire _GEN_370 = (casez_tmp_31 | casez_tmp_32) & casez_tmp_33;
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_34 = ldq_0_valid;
      5'b00001:
        casez_tmp_34 = ldq_1_valid;
      5'b00010:
        casez_tmp_34 = ldq_2_valid;
      5'b00011:
        casez_tmp_34 = ldq_3_valid;
      5'b00100:
        casez_tmp_34 = ldq_4_valid;
      5'b00101:
        casez_tmp_34 = ldq_5_valid;
      5'b00110:
        casez_tmp_34 = ldq_6_valid;
      5'b00111:
        casez_tmp_34 = ldq_7_valid;
      5'b01000:
        casez_tmp_34 = ldq_8_valid;
      5'b01001:
        casez_tmp_34 = ldq_9_valid;
      5'b01010:
        casez_tmp_34 = ldq_10_valid;
      5'b01011:
        casez_tmp_34 = ldq_11_valid;
      5'b01100:
        casez_tmp_34 = ldq_12_valid;
      5'b01101:
        casez_tmp_34 = ldq_13_valid;
      5'b01110:
        casez_tmp_34 = ldq_14_valid;
      5'b01111:
        casez_tmp_34 = ldq_15_valid;
      5'b10000:
        casez_tmp_34 = ldq_16_valid;
      5'b10001:
        casez_tmp_34 = ldq_17_valid;
      5'b10010:
        casez_tmp_34 = ldq_18_valid;
      5'b10011:
        casez_tmp_34 = ldq_19_valid;
      5'b10100:
        casez_tmp_34 = ldq_20_valid;
      5'b10101:
        casez_tmp_34 = ldq_21_valid;
      5'b10110:
        casez_tmp_34 = ldq_22_valid;
      5'b10111:
        casez_tmp_34 = ldq_23_valid;
      5'b11000:
        casez_tmp_34 = ldq_24_valid;
      5'b11001:
        casez_tmp_34 = ldq_25_valid;
      5'b11010:
        casez_tmp_34 = ldq_26_valid;
      5'b11011:
        casez_tmp_34 = ldq_27_valid;
      5'b11100:
        casez_tmp_34 = ldq_28_valid;
      5'b11101:
        casez_tmp_34 = ldq_29_valid;
      5'b11110:
        casez_tmp_34 = ldq_30_valid;
      default:
        casez_tmp_34 = ldq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_35 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_35 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_35 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_35 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_35 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_35 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_35 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_35 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_35 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_35 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_35 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_35 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_35 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_35 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_35 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_35 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_35 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_35 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_35 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_35 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_35 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_35 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_35 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_35 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_35 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_35 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_35 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_35 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_35 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_35 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_35 = ldq_30_bits_executed;
      default:
        casez_tmp_35 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_36 = ldq_0_bits_forward_std_val;
      5'b00001:
        casez_tmp_36 = ldq_1_bits_forward_std_val;
      5'b00010:
        casez_tmp_36 = ldq_2_bits_forward_std_val;
      5'b00011:
        casez_tmp_36 = ldq_3_bits_forward_std_val;
      5'b00100:
        casez_tmp_36 = ldq_4_bits_forward_std_val;
      5'b00101:
        casez_tmp_36 = ldq_5_bits_forward_std_val;
      5'b00110:
        casez_tmp_36 = ldq_6_bits_forward_std_val;
      5'b00111:
        casez_tmp_36 = ldq_7_bits_forward_std_val;
      5'b01000:
        casez_tmp_36 = ldq_8_bits_forward_std_val;
      5'b01001:
        casez_tmp_36 = ldq_9_bits_forward_std_val;
      5'b01010:
        casez_tmp_36 = ldq_10_bits_forward_std_val;
      5'b01011:
        casez_tmp_36 = ldq_11_bits_forward_std_val;
      5'b01100:
        casez_tmp_36 = ldq_12_bits_forward_std_val;
      5'b01101:
        casez_tmp_36 = ldq_13_bits_forward_std_val;
      5'b01110:
        casez_tmp_36 = ldq_14_bits_forward_std_val;
      5'b01111:
        casez_tmp_36 = ldq_15_bits_forward_std_val;
      5'b10000:
        casez_tmp_36 = ldq_16_bits_forward_std_val;
      5'b10001:
        casez_tmp_36 = ldq_17_bits_forward_std_val;
      5'b10010:
        casez_tmp_36 = ldq_18_bits_forward_std_val;
      5'b10011:
        casez_tmp_36 = ldq_19_bits_forward_std_val;
      5'b10100:
        casez_tmp_36 = ldq_20_bits_forward_std_val;
      5'b10101:
        casez_tmp_36 = ldq_21_bits_forward_std_val;
      5'b10110:
        casez_tmp_36 = ldq_22_bits_forward_std_val;
      5'b10111:
        casez_tmp_36 = ldq_23_bits_forward_std_val;
      5'b11000:
        casez_tmp_36 = ldq_24_bits_forward_std_val;
      5'b11001:
        casez_tmp_36 = ldq_25_bits_forward_std_val;
      5'b11010:
        casez_tmp_36 = ldq_26_bits_forward_std_val;
      5'b11011:
        casez_tmp_36 = ldq_27_bits_forward_std_val;
      5'b11100:
        casez_tmp_36 = ldq_28_bits_forward_std_val;
      5'b11101:
        casez_tmp_36 = ldq_29_bits_forward_std_val;
      5'b11110:
        casez_tmp_36 = ldq_30_bits_forward_std_val;
      default:
        casez_tmp_36 = ldq_31_bits_forward_std_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx_3)
      5'b00000:
        casez_tmp_37 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_37 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_37 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_37 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_37 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_37 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_37 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_37 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_37 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_37 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_37 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_37 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_37 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_37 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_37 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_37 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_37 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_37 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_37 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_37 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_37 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_37 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_37 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_37 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_37 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_37 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_37 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_37 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_37 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_37 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_37 = ldq_30_bits_succeeded;
      default:
        casez_tmp_37 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  wire _GEN_371 = (casez_tmp_35 | casez_tmp_36) & casez_tmp_37;
  wire _GEN_372 = dis_ld_val & ~reset;
  wire _GEN_373 = ~dis_ld_val & dis_st_val & ~reset;
  wire _GEN_374 = dis_ld_val_1 & ~reset;
  wire _GEN_375 = ~dis_ld_val_1 & dis_st_val_1 & ~reset;
  wire _GEN_376 = dis_ld_val_2 & ~reset;
  wire _GEN_377 = ~dis_ld_val_2 & dis_st_val_2 & ~reset;
  wire _GEN_378 = dis_ld_val_3 & ~reset;
  wire _GEN_379 = ~dis_ld_val_3 & dis_st_val_3 & ~reset;
  wire _GEN_380 = mem_xcpt_valids_0 & ~reset;
  wire _GEN_381 = mem_xcpt_valids_1 & ~reset;
  wire _GEN_382 = can_fire_load_incoming_0 & ~reset;
  wire _GEN_383 = _stq_idx_T & ~reset;
  wire _GEN_384 = _GEN_294 & ~reset;
  wire _GEN_385 = can_fire_load_incoming_1 & ~reset;
  wire _GEN_386 = ~can_fire_load_incoming_1 & will_fire_load_retry_1 & ~reset;
  wire _GEN_387 = ~can_fire_load_incoming_1 & ~will_fire_load_retry_1;
  wire _GEN_388 = _GEN_387 & will_fire_load_wakeup_1 & ~reset;
  wire _GEN_389 = _GEN_387 & ~will_fire_load_wakeup_1;
  wire _GEN_390 = _GEN_389 & will_fire_hella_incoming_1 & ~reset;
  wire _GEN_391 = _GEN_389 & ~will_fire_hella_incoming_1 & will_fire_hella_wakeup_1 & ~reset;
  wire _GEN_392 = _GEN_295 & ~reset;
  wire _GEN_393 = _GEN_296 & ~reset;
  wire _GEN_394 = _stq_bits_data_bits_T_2 & ~reset;
  wire _GEN_395 = _GEN_297 & ~reset;
  wire _GEN_396 = io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella;
  wire _GEN_397 = _GEN_396 & io_dmem_nack_0_bits_uop_uses_ldq & ~reset;
  wire _GEN_398 = _GEN_396 & ~io_dmem_nack_0_bits_uop_uses_ldq & ~reset;
  wire _GEN_399 = _GEN_298 & ~reset;
  wire _GEN_400 = io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & ~reset;
  wire _GEN_401 = _GEN_299 & ~reset;
  wire _GEN_402 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella;
  wire _GEN_403 = _GEN_402 & io_dmem_nack_1_bits_uop_uses_ldq & ~reset;
  wire _GEN_404 = _GEN_402 & ~io_dmem_nack_1_bits_uop_uses_ldq & ~reset;
  wire _GEN_405 = _GEN_300 & ~reset;
  wire _GEN_406 = io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & ~reset;
  wire _GEN_407 = ~commit_store & commit_load & ~reset;
  wire _GEN_408 = ~commit_store_1 & commit_load_1 & ~reset;
  wire _GEN_409 = ~commit_store_2 & commit_load_2 & ~reset;
  wire _GEN_410 = ~commit_store_3 & commit_load_3 & ~reset;
  `ifndef SYNTHESIS
    always @(posedge clock) begin
      if ((`PRINTF_COND_) & ~reset & ~_GEN_301)
        $fwrite(32'h80000002, "Assertion failed: stq_execute_head got off track.\n    at lsu.scala:222 assert (io.core.brupdate.b2.mispredict ||\n");
      if ((`PRINTF_COND_) & _GEN_372 & ~_GEN_302)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_372 & casez_tmp)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
      if ((`PRINTF_COND_) & _GEN_373 & ~_GEN_303)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_373 & casez_tmp_0)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_304)
        $fwrite(32'h80000002, "Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
      if ((`PRINTF_COND_) & _GEN_374 & ~_GEN_305)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_374 & casez_tmp_1)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
      if ((`PRINTF_COND_) & _GEN_375 & ~_GEN_306)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_375 & casez_tmp_2)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_307)
        $fwrite(32'h80000002, "Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
      if ((`PRINTF_COND_) & _GEN_376 & ~_GEN_308)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_376 & casez_tmp_3)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
      if ((`PRINTF_COND_) & _GEN_377 & ~_GEN_309)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_377 & casez_tmp_4)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_310)
        $fwrite(32'h80000002, "Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
      if ((`PRINTF_COND_) & _GEN_378 & ~_GEN_311)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq load tag.\n    at lsu.scala:316 assert (ld_enq_idx === io.core.dis_uops(w).bits.ldq_idx, \"[lsu] mismatch enq load tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_378 & casez_tmp_5)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting ldq entries\n    at lsu.scala:317 assert (!ldq(ld_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting ldq entries\")\n");
      if ((`PRINTF_COND_) & _GEN_379 & ~_GEN_312)
        $fwrite(32'h80000002, "Assertion failed: [lsu] mismatch enq store tag.\n    at lsu.scala:328 assert (st_enq_idx === io.core.dis_uops(w).bits.stq_idx, \"[lsu] mismatch enq store tag.\")\n");
      if ((`PRINTF_COND_) & _GEN_379 & casez_tmp_6)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Enqueuing uop is overwriting stq entries\n    at lsu.scala:329 assert (!stq(st_enq_idx).valid, \"[lsu] Enqueuing uop is overwriting stq entries\")\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_313)
        $fwrite(32'h80000002, "Assertion failed: A UOP is trying to go into both the LDQ and the STQ\n    at lsu.scala:340 assert(!(dis_ld_val && dis_st_val), \"A UOP is trying to go into both the LDQ and the STQ\")\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_315)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:566 assert(!(exe_req(w).valid && !(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) || will_fire_std_incoming(w) || will_fire_sfence(w))))\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_317)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:566 assert(!(exe_req(w).valid && !(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) || will_fire_std_incoming(w) || will_fire_sfence(w))))\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_318)
        $fwrite(32'h80000002, "Assertion failed: Some operations is proceeding down multiple pipes\n    at lsu.scala:577 assert((memWidth == 1).B ||\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_319)
        $fwrite(32'h80000002, "Assertion failed: SFENCE through hella interface not supported\n    at lsu.scala:592 assert(!(hella_state =/= h_ready && hella_req.cmd === rocket.M_SFENCE),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_320)
        $fwrite(32'h80000002, "Assertion failed: Fence is pretending to talk to the TLB\n    at lsu.scala:683 assert (!(dtlb.io.req(w).valid && exe_tlb_uop(w).is_fence), \"Fence is pretending to talk to the TLB\")\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_321)
        $fwrite(32'h80000002, "Assertion failed: A uop that's not a load or store-address is throwing a memory exception.\n    at lsu.scala:684 assert (!((will_fire_load_incoming(w) || will_fire_sta_incoming(w) || will_fire_stad_incoming(w)) &&\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_322)
        $fwrite(32'h80000002, "Assertion failed: Fence is pretending to talk to the TLB\n    at lsu.scala:683 assert (!(dtlb.io.req(w).valid && exe_tlb_uop(w).is_fence), \"Fence is pretending to talk to the TLB\")\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_323)
        $fwrite(32'h80000002, "Assertion failed: A uop that's not a load or store-address is throwing a memory exception.\n    at lsu.scala:684 assert (!((will_fire_load_incoming(w) || will_fire_sta_incoming(w) || will_fire_stad_incoming(w)) &&\n");
      if ((`PRINTF_COND_) & ~reset & ~_GEN_324)
        $fwrite(32'h80000002, "Assertion failed: [lsu] paddrs should match.\n    at lsu.scala:715 assert (exe_tlb_paddr(w) === dtlb.io.resp(w).paddr || exe_req(w).bits.sfence.valid, \"[lsu] paddrs should match.\")\n");
      if ((`PRINTF_COND_) & _GEN_380 & ~REG)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:719 assert(RegNext(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) ||\n");
      if ((`PRINTF_COND_) & _GEN_380 & ~_GEN_325)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:722 assert(mem_xcpt_uops(w).uses_ldq ^ mem_xcpt_uops(w).uses_stq)\n");
      if ((`PRINTF_COND_) & ~reset & ~_GEN_326)
        $fwrite(32'h80000002, "Assertion failed: [lsu] paddrs should match.\n    at lsu.scala:715 assert (exe_tlb_paddr(w) === dtlb.io.resp(w).paddr || exe_req(w).bits.sfence.valid, \"[lsu] paddrs should match.\")\n");
      if ((`PRINTF_COND_) & _GEN_381 & ~REG_1)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:719 assert(RegNext(will_fire_load_incoming(w) || will_fire_stad_incoming(w) || will_fire_sta_incoming(w) ||\n");
      if ((`PRINTF_COND_) & _GEN_381 & ~_GEN_327)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:722 assert(mem_xcpt_uops(w).uses_ldq ^ mem_xcpt_uops(w).uses_stq)\n");
      if ((`PRINTF_COND_) & _GEN_382 & casez_tmp_8)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:773 assert(!ldq_incoming_e(w).bits.executed)\n");
      if ((`PRINTF_COND_) & _GEN_382 & _GEN_328)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Incoming load is overwriting a valid address\n    at lsu.scala:845 assert(!(will_fire_load_incoming(w) && ldq_incoming_e(w).bits.addr.valid),\n");
      if ((`PRINTF_COND_) & _GEN_383 & _GEN_329)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Incoming store is overwriting a valid address\n    at lsu.scala:859 assert(!(will_fire_sta_incoming(w) && stq_incoming_e(w).bits.addr.valid),\n");
      if ((`PRINTF_COND_) & _GEN_384 & casez_tmp_18)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Incoming store is overwriting a valid data entry\n    at lsu.scala:878 assert(!(stq(sidx).bits.data.valid),\n");
      if ((`PRINTF_COND_) & _GEN_385 & casez_tmp_10)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:773 assert(!ldq_incoming_e(w).bits.executed)\n");
      if ((`PRINTF_COND_) & _GEN_386 & casez_tmp_17)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:780 assert(!ldq_retry_e.bits.executed)\n");
      if ((`PRINTF_COND_) & _GEN_388 & ~_GEN_330)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:802 assert(!ldq_wakeup_e.bits.executed && !ldq_wakeup_e.bits.addr_is_virtual)\n");
      if ((`PRINTF_COND_) & _GEN_390 & ~_GEN_140251)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:804 assert(hella_state === h_s1)\n");
      if ((`PRINTF_COND_) & _GEN_391 & ~_GEN_140205)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:821 assert(hella_state === h_replay)\n");
      if ((`PRINTF_COND_) & _GEN_392 & _GEN_331)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Incoming load is overwriting a valid address\n    at lsu.scala:845 assert(!(will_fire_load_incoming(w) && ldq_incoming_e(w).bits.addr.valid),\n");
      if ((`PRINTF_COND_) & _GEN_393 & _GEN_332)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Incoming store is overwriting a valid address\n    at lsu.scala:859 assert(!(will_fire_sta_incoming(w) && stq_incoming_e(w).bits.addr.valid),\n");
      if ((`PRINTF_COND_) & _GEN_394 & casez_tmp_19)
        $fwrite(32'h80000002, "Assertion failed: [lsu] Incoming store is overwriting a valid data entry\n    at lsu.scala:878 assert(!(stq(sidx).bits.data.valid),\n");
      if ((`PRINTF_COND_) & _GEN_395 & ~_GEN_333)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1291 assert(hella_state === h_wait || hella_state === h_dead)\n");
      if ((`PRINTF_COND_) & _GEN_397 & ~casez_tmp_20)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1295 assert(ldq(io.dmem.nack(w).bits.uop.ldq_idx).bits.executed)\n");
      if ((`PRINTF_COND_) & _GEN_398 & ~io_dmem_nack_0_bits_uop_uses_stq)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1301 assert(io.dmem.nack(w).bits.uop.uses_stq)\n");
      if ((`PRINTF_COND_) & _GEN_399 & io_dmem_resp_0_bits_is_hella)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1312 assert(!io.dmem.resp(w).bits.is_hella)\n");
      if ((`PRINTF_COND_) & _GEN_399 & ~_GEN_334)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1324 assert(send_iresp ^ send_fresp)\n");
      if ((`PRINTF_COND_) & _GEN_400 & io_dmem_resp_0_bits_is_hella)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1332 assert(!io.dmem.resp(w).bits.is_hella)\n");
      if ((`PRINTF_COND_) & _GEN_401 & ~_GEN_333)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1291 assert(hella_state === h_wait || hella_state === h_dead)\n");
      if ((`PRINTF_COND_) & _GEN_403 & ~casez_tmp_21)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1295 assert(ldq(io.dmem.nack(w).bits.uop.ldq_idx).bits.executed)\n");
      if ((`PRINTF_COND_) & _GEN_404 & ~io_dmem_nack_1_bits_uop_uses_stq)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1301 assert(io.dmem.nack(w).bits.uop.uses_stq)\n");
      if ((`PRINTF_COND_) & _GEN_405 & io_dmem_resp_1_bits_is_hella)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1312 assert(!io.dmem.resp(w).bits.is_hella)\n");
      if ((`PRINTF_COND_) & _GEN_405 & ~_GEN_335)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1324 assert(send_iresp ^ send_fresp)\n");
      if ((`PRINTF_COND_) & _GEN_406 & io_dmem_resp_1_bits_is_hella)
        $fwrite(32'h80000002, "Assertion failed\n    at lsu.scala:1332 assert(!io.dmem.resp(w).bits.is_hella)\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_336)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_337)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_338)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_339)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_340)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_341)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_342)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_343)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_344)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_345)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_346)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_347)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_348)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_349)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_350)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_351)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_352)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_353)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_354)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_355)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_356)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_357)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_358)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_359)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_360)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_361)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_362)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_363)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_364)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_365)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_366)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & ~reset & _GEN_367)
        $fwrite(32'h80000002, "Assertion failed: Branch is trying to clear a committed store.\n    at lsu.scala:1419 assert (!(IsKilledByBranch(io.core.brupdate, stq(i).bits.uop) && stq(i).valid && stq(i).bits.committed),\n");
      if ((`PRINTF_COND_) & _GEN_407 & ~casez_tmp_22)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_407 & ~_GEN_368)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
      if ((`PRINTF_COND_) & _GEN_408 & ~casez_tmp_26)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_408 & ~_GEN_369)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
      if ((`PRINTF_COND_) & _GEN_409 & ~casez_tmp_30)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_409 & ~_GEN_370)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
      if ((`PRINTF_COND_) & _GEN_410 & ~casez_tmp_34)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-allocated load entry.\n    at lsu.scala:1461 assert (ldq(idx).valid, \"[lsu] trying to commit an un-allocated load entry.\")\n");
      if ((`PRINTF_COND_) & _GEN_410 & ~_GEN_371)
        $fwrite(32'h80000002, "Assertion failed: [lsu] trying to commit an un-executed load entry.\n    at lsu.scala:1462 assert ((ldq(idx).bits.executed || ldq(idx).bits.forward_std_val) && ldq(idx).bits.succeeded ,\n");
    end // always @(posedge)
  `endif // not def SYNTHESIS
  wire _GEN_411 = dis_ld_val | ~_GEN_131;
  wire _GEN_412 = dis_ld_val | ~_GEN_136;
  wire _GEN_413 = dis_ld_val | ~_GEN_140;
  wire _GEN_414 = dis_ld_val | ~_GEN_144;
  wire _GEN_415 = dis_ld_val | ~_GEN_148;
  wire _GEN_416 = dis_ld_val | ~_GEN_152;
  wire _GEN_417 = dis_ld_val | ~_GEN_156;
  wire _GEN_418 = dis_ld_val | ~_GEN_160;
  wire _GEN_419 = dis_ld_val | ~_GEN_164;
  wire _GEN_420 = dis_ld_val | ~_GEN_168;
  wire _GEN_421 = dis_ld_val | ~_GEN_172;
  wire _GEN_422 = dis_ld_val | ~_GEN_176;
  wire _GEN_423 = dis_ld_val | ~_GEN_180;
  wire _GEN_424 = dis_ld_val | ~_GEN_184;
  wire _GEN_425 = dis_ld_val | ~_GEN_188;
  wire _GEN_426 = dis_ld_val | ~_GEN_192;
  wire _GEN_427 = dis_ld_val | ~_GEN_196;
  wire _GEN_428 = dis_ld_val | ~_GEN_200;
  wire _GEN_429 = dis_ld_val | ~_GEN_204;
  wire _GEN_430 = dis_ld_val | ~_GEN_208;
  wire _GEN_431 = dis_ld_val | ~_GEN_212;
  wire _GEN_432 = dis_ld_val | ~_GEN_216;
  wire _GEN_433 = dis_ld_val | ~_GEN_220;
  wire _GEN_434 = dis_ld_val | ~_GEN_224;
  wire _GEN_435 = dis_ld_val | ~_GEN_228;
  wire _GEN_436 = dis_ld_val | ~_GEN_232;
  wire _GEN_437 = dis_ld_val | ~_GEN_236;
  wire _GEN_438 = dis_ld_val | ~_GEN_240;
  wire _GEN_439 = dis_ld_val | ~_GEN_244;
  wire _GEN_440 = dis_ld_val | ~_GEN_248;
  wire _GEN_441 = dis_ld_val | ~_GEN_252;
  wire _GEN_442 = dis_ld_val | ~_GEN_256;
  wire _GEN_443 = dis_ld_val_1 | ~_GEN_132;
  wire _GEN_444 = dis_ld_val_1 | ~_GEN_137;
  wire _GEN_445 = dis_ld_val_1 | ~_GEN_141;
  wire _GEN_446 = dis_ld_val_1 | ~_GEN_145;
  wire _GEN_447 = dis_ld_val_1 | ~_GEN_149;
  wire _GEN_448 = dis_ld_val_1 | ~_GEN_153;
  wire _GEN_449 = dis_ld_val_1 | ~_GEN_157;
  wire _GEN_450 = dis_ld_val_1 | ~_GEN_161;
  wire _GEN_451 = dis_ld_val_1 | ~_GEN_165;
  wire _GEN_452 = dis_ld_val_1 | ~_GEN_169;
  wire _GEN_453 = dis_ld_val_1 | ~_GEN_173;
  wire _GEN_454 = dis_ld_val_1 | ~_GEN_177;
  wire _GEN_455 = dis_ld_val_1 | ~_GEN_181;
  wire _GEN_456 = dis_ld_val_1 | ~_GEN_185;
  wire _GEN_457 = dis_ld_val_1 | ~_GEN_189;
  wire _GEN_458 = dis_ld_val_1 | ~_GEN_193;
  wire _GEN_459 = dis_ld_val_1 | ~_GEN_197;
  wire _GEN_460 = dis_ld_val_1 | ~_GEN_201;
  wire _GEN_461 = dis_ld_val_1 | ~_GEN_205;
  wire _GEN_462 = dis_ld_val_1 | ~_GEN_209;
  wire _GEN_463 = dis_ld_val_1 | ~_GEN_213;
  wire _GEN_464 = dis_ld_val_1 | ~_GEN_217;
  wire _GEN_465 = dis_ld_val_1 | ~_GEN_221;
  wire _GEN_466 = dis_ld_val_1 | ~_GEN_225;
  wire _GEN_467 = dis_ld_val_1 | ~_GEN_229;
  wire _GEN_468 = dis_ld_val_1 | ~_GEN_233;
  wire _GEN_469 = dis_ld_val_1 | ~_GEN_237;
  wire _GEN_470 = dis_ld_val_1 | ~_GEN_241;
  wire _GEN_471 = dis_ld_val_1 | ~_GEN_245;
  wire _GEN_472 = dis_ld_val_1 | ~_GEN_249;
  wire _GEN_473 = dis_ld_val_1 | ~_GEN_253;
  wire _GEN_474 = dis_ld_val_1 | ~_GEN_257;
  wire _GEN_475 = dis_ld_val_2 | ~_GEN_133;
  wire _GEN_476 = dis_ld_val_2 | ~_GEN_138;
  wire _GEN_477 = dis_ld_val_2 | ~_GEN_142;
  wire _GEN_478 = dis_ld_val_2 | ~_GEN_146;
  wire _GEN_479 = dis_ld_val_2 | ~_GEN_150;
  wire _GEN_480 = dis_ld_val_2 | ~_GEN_154;
  wire _GEN_481 = dis_ld_val_2 | ~_GEN_158;
  wire _GEN_482 = dis_ld_val_2 | ~_GEN_162;
  wire _GEN_483 = dis_ld_val_2 | ~_GEN_166;
  wire _GEN_484 = dis_ld_val_2 | ~_GEN_170;
  wire _GEN_485 = dis_ld_val_2 | ~_GEN_174;
  wire _GEN_486 = dis_ld_val_2 | ~_GEN_178;
  wire _GEN_487 = dis_ld_val_2 | ~_GEN_182;
  wire _GEN_488 = dis_ld_val_2 | ~_GEN_186;
  wire _GEN_489 = dis_ld_val_2 | ~_GEN_190;
  wire _GEN_490 = dis_ld_val_2 | ~_GEN_194;
  wire _GEN_491 = dis_ld_val_2 | ~_GEN_198;
  wire _GEN_492 = dis_ld_val_2 | ~_GEN_202;
  wire _GEN_493 = dis_ld_val_2 | ~_GEN_206;
  wire _GEN_494 = dis_ld_val_2 | ~_GEN_210;
  wire _GEN_495 = dis_ld_val_2 | ~_GEN_214;
  wire _GEN_496 = dis_ld_val_2 | ~_GEN_218;
  wire _GEN_497 = dis_ld_val_2 | ~_GEN_222;
  wire _GEN_498 = dis_ld_val_2 | ~_GEN_226;
  wire _GEN_499 = dis_ld_val_2 | ~_GEN_230;
  wire _GEN_500 = dis_ld_val_2 | ~_GEN_234;
  wire _GEN_501 = dis_ld_val_2 | ~_GEN_238;
  wire _GEN_502 = dis_ld_val_2 | ~_GEN_242;
  wire _GEN_503 = dis_ld_val_2 | ~_GEN_246;
  wire _GEN_504 = dis_ld_val_2 | ~_GEN_250;
  wire _GEN_505 = dis_ld_val_2 | ~_GEN_254;
  wire _GEN_506 = dis_ld_val_2 | ~_GEN_258;
  wire _GEN_507 = dis_ld_val_3 | ~_GEN_134;
  wire _GEN_508 = dis_ld_val_3 | ~_GEN_139;
  wire _GEN_509 = dis_ld_val_3 | ~_GEN_143;
  wire _GEN_510 = dis_ld_val_3 | ~_GEN_147;
  wire _GEN_511 = dis_ld_val_3 | ~_GEN_151;
  wire _GEN_512 = dis_ld_val_3 | ~_GEN_155;
  wire _GEN_513 = dis_ld_val_3 | ~_GEN_159;
  wire _GEN_514 = dis_ld_val_3 | ~_GEN_163;
  wire _GEN_515 = dis_ld_val_3 | ~_GEN_167;
  wire _GEN_516 = dis_ld_val_3 | ~_GEN_171;
  wire _GEN_517 = dis_ld_val_3 | ~_GEN_175;
  wire _GEN_518 = dis_ld_val_3 | ~_GEN_179;
  wire _GEN_519 = dis_ld_val_3 | ~_GEN_183;
  wire _GEN_520 = dis_ld_val_3 | ~_GEN_187;
  wire _GEN_521 = dis_ld_val_3 | ~_GEN_191;
  wire _GEN_522 = dis_ld_val_3 | ~_GEN_195;
  wire _GEN_523 = dis_ld_val_3 | ~_GEN_199;
  wire _GEN_524 = dis_ld_val_3 | ~_GEN_203;
  wire _GEN_525 = dis_ld_val_3 | ~_GEN_207;
  wire _GEN_526 = dis_ld_val_3 | ~_GEN_211;
  wire _GEN_527 = dis_ld_val_3 | ~_GEN_215;
  wire _GEN_528 = dis_ld_val_3 | ~_GEN_219;
  wire _GEN_529 = dis_ld_val_3 | ~_GEN_223;
  wire _GEN_530 = dis_ld_val_3 | ~_GEN_227;
  wire _GEN_531 = dis_ld_val_3 | ~_GEN_231;
  wire _GEN_532 = dis_ld_val_3 | ~_GEN_235;
  wire _GEN_533 = dis_ld_val_3 | ~_GEN_239;
  wire _GEN_534 = dis_ld_val_3 | ~_GEN_243;
  wire _GEN_535 = dis_ld_val_3 | ~_GEN_247;
  wire _GEN_536 = dis_ld_val_3 | ~_GEN_251;
  wire _GEN_537 = dis_ld_val_3 | ~_GEN_255;
  wire _GEN_538 = dis_ld_val_3 | ~_GEN_259;
  always @(posedge clock) begin
    if (~reset)
      assert__assert: assert(_GEN_301);
    if (_GEN_372) begin
      assert__assert_1: assert(_GEN_302);
      assert__assert_2: assert(~casez_tmp);
    end
    if (_GEN_373) begin
      assert__assert_3: assert(_GEN_303);
      assert__assert_4: assert(~casez_tmp_0);
    end
    if (~reset)
      assert__assert_5: assert(~_GEN_304);
    if (_GEN_374) begin
      assert__assert_6: assert(_GEN_305);
      assert__assert_7: assert(~casez_tmp_1);
    end
    if (_GEN_375) begin
      assert__assert_8: assert(_GEN_306);
      assert__assert_9: assert(~casez_tmp_2);
    end
    if (~reset)
      assert__assert_10: assert(~_GEN_307);
    if (_GEN_376) begin
      assert__assert_11: assert(_GEN_308);
      assert__assert_12: assert(~casez_tmp_3);
    end
    if (_GEN_377) begin
      assert__assert_13: assert(_GEN_309);
      assert__assert_14: assert(~casez_tmp_4);
    end
    if (~reset)
      assert__assert_15: assert(~_GEN_310);
    if (_GEN_378) begin
      assert__assert_16: assert(_GEN_311);
      assert__assert_17: assert(~casez_tmp_5);
    end
    if (_GEN_379) begin
      assert__assert_18: assert(_GEN_312);
      assert__assert_19: assert(~casez_tmp_6);
    end
    if (~reset) begin
      assert__assert_20: assert(~_GEN_313);
      assert__assert_21: assert(~_GEN_315);
      assert__assert_22: assert(~_GEN_317);
      assert__assert_23: assert(~_GEN_318);
      assert__assert_24: assert(~_GEN_319);
      assert__assert_25: assert(~_GEN_320);
      assert__assert_26: assert(~_GEN_321);
      assert__assert_27: assert(~_GEN_322);
      assert__assert_28: assert(~_GEN_323);
      assert__assert_29: assert(_GEN_324);
    end
    if (_GEN_380) begin
      assert__assert_30: assert(REG);
      assert__assert_31: assert(_GEN_325);
    end
    if (~reset)
      assert__assert_32: assert(_GEN_326);
    if (_GEN_381) begin
      assert__assert_33: assert(REG_1);
      assert__assert_34: assert(_GEN_327);
    end
    if (_GEN_382) begin
      assert__assert_35: assert(~casez_tmp_8);
      assert__assert_40: assert(~_GEN_328);
    end
    if (_GEN_383)
      assert__assert_41: assert(~_GEN_329);
    if (_GEN_384)
      assert__assert_42: assert(~casez_tmp_18);
    if (_GEN_385)
      assert__assert_43: assert(~casez_tmp_10);
    if (_GEN_386)
      assert__assert_44: assert(~casez_tmp_17);
    if (_GEN_388)
      assert__assert_45: assert(_GEN_330);
    if (_GEN_390)
      assert__assert_46: assert(_GEN_140251);
    if (_GEN_391)
      assert__assert_47: assert(_GEN_140205);
    if (_GEN_392)
      assert__assert_48: assert(~_GEN_331);
    if (_GEN_393)
      assert__assert_49: assert(~_GEN_332);
    if (_GEN_394)
      assert__assert_50: assert(~casez_tmp_19);
    if (_GEN_395)
      assert__assert_51: assert(_GEN_333);
    if (_GEN_397)
      assert__assert_52: assert(casez_tmp_20);
    if (_GEN_398)
      assert__assert_53: assert(io_dmem_nack_0_bits_uop_uses_stq);
    if (_GEN_399) begin
      assert__assert_54: assert(~io_dmem_resp_0_bits_is_hella);
      assert__assert_55: assert(_GEN_334);
    end
    if (_GEN_400)
      assert__assert_56: assert(~io_dmem_resp_0_bits_is_hella);
    if (_GEN_401)
      assert__assert_57: assert(_GEN_333);
    if (_GEN_403)
      assert__assert_58: assert(casez_tmp_21);
    if (_GEN_404)
      assert__assert_59: assert(io_dmem_nack_1_bits_uop_uses_stq);
    if (_GEN_405) begin
      assert__assert_60: assert(~io_dmem_resp_1_bits_is_hella);
      assert__assert_61: assert(_GEN_335);
    end
    if (_GEN_406)
      assert__assert_62: assert(~io_dmem_resp_1_bits_is_hella);
    if (~reset) begin
      assert__assert_63: assert(~_GEN_336);
      assert__assert_64: assert(~_GEN_337);
      assert__assert_65: assert(~_GEN_338);
      assert__assert_66: assert(~_GEN_339);
      assert__assert_67: assert(~_GEN_340);
      assert__assert_68: assert(~_GEN_341);
      assert__assert_69: assert(~_GEN_342);
      assert__assert_70: assert(~_GEN_343);
      assert__assert_71: assert(~_GEN_344);
      assert__assert_72: assert(~_GEN_345);
      assert__assert_73: assert(~_GEN_346);
      assert__assert_74: assert(~_GEN_347);
      assert__assert_75: assert(~_GEN_348);
      assert__assert_76: assert(~_GEN_349);
      assert__assert_77: assert(~_GEN_350);
      assert__assert_78: assert(~_GEN_351);
      assert__assert_79: assert(~_GEN_352);
      assert__assert_80: assert(~_GEN_353);
      assert__assert_81: assert(~_GEN_354);
      assert__assert_82: assert(~_GEN_355);
      assert__assert_83: assert(~_GEN_356);
      assert__assert_84: assert(~_GEN_357);
      assert__assert_85: assert(~_GEN_358);
      assert__assert_86: assert(~_GEN_359);
      assert__assert_87: assert(~_GEN_360);
      assert__assert_88: assert(~_GEN_361);
      assert__assert_89: assert(~_GEN_362);
      assert__assert_90: assert(~_GEN_363);
      assert__assert_91: assert(~_GEN_364);
      assert__assert_92: assert(~_GEN_365);
      assert__assert_93: assert(~_GEN_366);
      assert__assert_94: assert(~_GEN_367);
    end
    if (_GEN_407) begin
      assert__assert_95: assert(casez_tmp_22);
      assert__assert_96: assert(_GEN_368);
    end
    if (_GEN_408) begin
      assert__assert_97: assert(casez_tmp_26);
      assert__assert_98: assert(_GEN_369);
    end
    if (_GEN_409) begin
      assert__assert_99: assert(casez_tmp_30);
      assert__assert_100: assert(_GEN_370);
    end
    if (_GEN_410) begin
      assert__assert_101: assert(casez_tmp_34);
      assert__assert_102: assert(_GEN_371);
    end
    if (_GEN_3) begin
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_4) begin
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_5) begin
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_6) begin
      ldq_0_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_0_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_0_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_7) begin
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_8) begin
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_9) begin
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_10) begin
      ldq_1_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_1_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_1_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_11) begin
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_12) begin
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_13) begin
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_14) begin
      ldq_2_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_2_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_2_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_15) begin
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_16) begin
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_17) begin
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_18) begin
      ldq_3_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_3_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_3_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_19) begin
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_20) begin
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_21) begin
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_22) begin
      ldq_4_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_4_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_4_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_23) begin
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_24) begin
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_25) begin
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_26) begin
      ldq_5_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_5_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_5_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_27) begin
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_28) begin
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_29) begin
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_30) begin
      ldq_6_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_6_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_6_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_31) begin
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_32) begin
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_33) begin
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_34) begin
      ldq_7_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_7_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_7_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_35) begin
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_36) begin
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_37) begin
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_38) begin
      ldq_8_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_8_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_8_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_39) begin
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_40) begin
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_41) begin
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_42) begin
      ldq_9_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_9_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_9_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_43) begin
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_44) begin
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_45) begin
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_46) begin
      ldq_10_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_10_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_10_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_47) begin
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_48) begin
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_49) begin
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_50) begin
      ldq_11_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_11_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_11_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_51) begin
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_52) begin
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_53) begin
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_54) begin
      ldq_12_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_12_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_12_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_55) begin
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_56) begin
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_57) begin
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_58) begin
      ldq_13_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_13_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_13_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_59) begin
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_60) begin
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_61) begin
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_62) begin
      ldq_14_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_14_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_14_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_63) begin
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_64) begin
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_65) begin
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_66) begin
      ldq_15_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_15_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_15_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_67) begin
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_68) begin
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_69) begin
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_70) begin
      ldq_16_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_16_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_16_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_71) begin
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_72) begin
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_73) begin
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_74) begin
      ldq_17_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_17_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_17_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_75) begin
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_76) begin
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_77) begin
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_78) begin
      ldq_18_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_18_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_18_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_79) begin
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_80) begin
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_81) begin
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_82) begin
      ldq_19_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_19_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_19_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_83) begin
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_84) begin
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_85) begin
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_86) begin
      ldq_20_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_20_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_20_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_87) begin
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_88) begin
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_89) begin
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_90) begin
      ldq_21_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_21_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_21_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_91) begin
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_92) begin
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_93) begin
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_94) begin
      ldq_22_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_22_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_22_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_95) begin
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_96) begin
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_97) begin
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_98) begin
      ldq_23_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_23_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_23_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_99) begin
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_100) begin
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_101) begin
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_102) begin
      ldq_24_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_24_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_24_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_103) begin
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_104) begin
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_105) begin
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_106) begin
      ldq_25_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_25_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_25_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_107) begin
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_108) begin
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_109) begin
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_110) begin
      ldq_26_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_26_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_26_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_111) begin
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_112) begin
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_113) begin
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_114) begin
      ldq_27_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_27_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_27_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_115) begin
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_116) begin
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_117) begin
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_118) begin
      ldq_28_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_28_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_28_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_119) begin
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_120) begin
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_121) begin
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_122) begin
      ldq_29_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_29_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_29_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_123) begin
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_124) begin
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_125) begin
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_126) begin
      ldq_30_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_30_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_30_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    if (_GEN_127) begin
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_3_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_3_bits_ctrl_is_sta;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_3_bits_is_fence;
    end
    else if (_GEN_128) begin
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_2_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_2_bits_ctrl_is_sta;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_2_bits_is_fence;
    end
    else if (_GEN_129) begin
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_1_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_1_bits_ctrl_is_sta;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_1_bits_is_fence;
    end
    else if (_GEN_130) begin
      ldq_31_bits_uop_ctrl_is_load <= io_core_dis_uops_0_bits_ctrl_is_load;
      ldq_31_bits_uop_ctrl_is_sta <= io_core_dis_uops_0_bits_ctrl_is_sta;
      ldq_31_bits_uop_is_fence <= io_core_dis_uops_0_bits_is_fence;
    end
    stq_0_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_507 ? (_GEN_475 ? (_GEN_443 ? (_GEN_411 ? stq_0_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_0_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_507 ? (_GEN_475 ? (_GEN_443 ? (_GEN_411 ? stq_0_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_1_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_508 ? (_GEN_476 ? (_GEN_444 ? (_GEN_412 ? stq_1_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_1_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_508 ? (_GEN_476 ? (_GEN_444 ? (_GEN_412 ? stq_1_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_2_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_509 ? (_GEN_477 ? (_GEN_445 ? (_GEN_413 ? stq_2_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_2_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_509 ? (_GEN_477 ? (_GEN_445 ? (_GEN_413 ? stq_2_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_3_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_510 ? (_GEN_478 ? (_GEN_446 ? (_GEN_414 ? stq_3_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_3_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_510 ? (_GEN_478 ? (_GEN_446 ? (_GEN_414 ? stq_3_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_4_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_511 ? (_GEN_479 ? (_GEN_447 ? (_GEN_415 ? stq_4_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_4_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_511 ? (_GEN_479 ? (_GEN_447 ? (_GEN_415 ? stq_4_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_5_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_512 ? (_GEN_480 ? (_GEN_448 ? (_GEN_416 ? stq_5_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_5_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_512 ? (_GEN_480 ? (_GEN_448 ? (_GEN_416 ? stq_5_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_6_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_513 ? (_GEN_481 ? (_GEN_449 ? (_GEN_417 ? stq_6_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_6_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_513 ? (_GEN_481 ? (_GEN_449 ? (_GEN_417 ? stq_6_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_7_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_514 ? (_GEN_482 ? (_GEN_450 ? (_GEN_418 ? stq_7_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_7_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_514 ? (_GEN_482 ? (_GEN_450 ? (_GEN_418 ? stq_7_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_8_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_515 ? (_GEN_483 ? (_GEN_451 ? (_GEN_419 ? stq_8_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_8_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_515 ? (_GEN_483 ? (_GEN_451 ? (_GEN_419 ? stq_8_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_9_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_516 ? (_GEN_484 ? (_GEN_452 ? (_GEN_420 ? stq_9_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_9_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_516 ? (_GEN_484 ? (_GEN_452 ? (_GEN_420 ? stq_9_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_10_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_517 ? (_GEN_485 ? (_GEN_453 ? (_GEN_421 ? stq_10_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_10_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_517 ? (_GEN_485 ? (_GEN_453 ? (_GEN_421 ? stq_10_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_11_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_518 ? (_GEN_486 ? (_GEN_454 ? (_GEN_422 ? stq_11_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_11_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_518 ? (_GEN_486 ? (_GEN_454 ? (_GEN_422 ? stq_11_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_12_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_519 ? (_GEN_487 ? (_GEN_455 ? (_GEN_423 ? stq_12_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_12_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_519 ? (_GEN_487 ? (_GEN_455 ? (_GEN_423 ? stq_12_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_13_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_520 ? (_GEN_488 ? (_GEN_456 ? (_GEN_424 ? stq_13_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_13_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_520 ? (_GEN_488 ? (_GEN_456 ? (_GEN_424 ? stq_13_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_14_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_521 ? (_GEN_489 ? (_GEN_457 ? (_GEN_425 ? stq_14_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_14_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_521 ? (_GEN_489 ? (_GEN_457 ? (_GEN_425 ? stq_14_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_15_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_522 ? (_GEN_490 ? (_GEN_458 ? (_GEN_426 ? stq_15_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_15_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_522 ? (_GEN_490 ? (_GEN_458 ? (_GEN_426 ? stq_15_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_16_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_523 ? (_GEN_491 ? (_GEN_459 ? (_GEN_427 ? stq_16_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_16_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_523 ? (_GEN_491 ? (_GEN_459 ? (_GEN_427 ? stq_16_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_17_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_524 ? (_GEN_492 ? (_GEN_460 ? (_GEN_428 ? stq_17_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_17_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_524 ? (_GEN_492 ? (_GEN_460 ? (_GEN_428 ? stq_17_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_18_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_525 ? (_GEN_493 ? (_GEN_461 ? (_GEN_429 ? stq_18_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_18_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_525 ? (_GEN_493 ? (_GEN_461 ? (_GEN_429 ? stq_18_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_19_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_526 ? (_GEN_494 ? (_GEN_462 ? (_GEN_430 ? stq_19_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_19_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_526 ? (_GEN_494 ? (_GEN_462 ? (_GEN_430 ? stq_19_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_20_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_527 ? (_GEN_495 ? (_GEN_463 ? (_GEN_431 ? stq_20_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_20_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_527 ? (_GEN_495 ? (_GEN_463 ? (_GEN_431 ? stq_20_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_21_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_528 ? (_GEN_496 ? (_GEN_464 ? (_GEN_432 ? stq_21_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_21_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_528 ? (_GEN_496 ? (_GEN_464 ? (_GEN_432 ? stq_21_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_22_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_529 ? (_GEN_497 ? (_GEN_465 ? (_GEN_433 ? stq_22_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_22_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_529 ? (_GEN_497 ? (_GEN_465 ? (_GEN_433 ? stq_22_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_23_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_530 ? (_GEN_498 ? (_GEN_466 ? (_GEN_434 ? stq_23_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_23_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_530 ? (_GEN_498 ? (_GEN_466 ? (_GEN_434 ? stq_23_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_24_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_531 ? (_GEN_499 ? (_GEN_467 ? (_GEN_435 ? stq_24_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_24_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_531 ? (_GEN_499 ? (_GEN_467 ? (_GEN_435 ? stq_24_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_25_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_532 ? (_GEN_500 ? (_GEN_468 ? (_GEN_436 ? stq_25_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_25_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_532 ? (_GEN_500 ? (_GEN_468 ? (_GEN_436 ? stq_25_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_26_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_533 ? (_GEN_501 ? (_GEN_469 ? (_GEN_437 ? stq_26_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_26_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_533 ? (_GEN_501 ? (_GEN_469 ? (_GEN_437 ? stq_26_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_27_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_534 ? (_GEN_502 ? (_GEN_470 ? (_GEN_438 ? stq_27_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_27_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_534 ? (_GEN_502 ? (_GEN_470 ? (_GEN_438 ? stq_27_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_28_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_535 ? (_GEN_503 ? (_GEN_471 ? (_GEN_439 ? stq_28_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_28_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_535 ? (_GEN_503 ? (_GEN_471 ? (_GEN_439 ? stq_28_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_29_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_536 ? (_GEN_504 ? (_GEN_472 ? (_GEN_440 ? stq_29_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_29_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_536 ? (_GEN_504 ? (_GEN_472 ? (_GEN_440 ? stq_29_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_30_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_537 ? (_GEN_505 ? (_GEN_473 ? (_GEN_441 ? stq_30_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_30_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_537 ? (_GEN_505 ? (_GEN_473 ? (_GEN_441 ? stq_30_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    stq_31_bits_uop_ctrl_is_load <= ~_GEN_135 & (_GEN_538 ? (_GEN_506 ? (_GEN_474 ? (_GEN_442 ? stq_31_bits_uop_ctrl_is_load : io_core_dis_uops_0_bits_ctrl_is_load) : io_core_dis_uops_1_bits_ctrl_is_load) : io_core_dis_uops_2_bits_ctrl_is_load) : io_core_dis_uops_3_bits_ctrl_is_load);
    stq_31_bits_uop_ctrl_is_sta <= ~_GEN_135 & (_GEN_538 ? (_GEN_506 ? (_GEN_474 ? (_GEN_442 ? stq_31_bits_uop_ctrl_is_sta : io_core_dis_uops_0_bits_ctrl_is_sta) : io_core_dis_uops_1_bits_ctrl_is_sta) : io_core_dis_uops_2_bits_ctrl_is_sta) : io_core_dis_uops_3_bits_ctrl_is_sta);
    mem_xcpt_uops_0_uses_stq <= exe_tlb_uop_0_uses_stq;
    mem_xcpt_uops_1_uses_stq <= exe_tlb_uop_1_uses_stq;
    REG <= _GEN_314;
    REG_1 <= _GEN_316 | will_fire_load_retry_1 | will_fire_sta_retry_1;
  end // always @(posedge)
endmodule

