// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

module TLROM(
  input         clock,
                reset,
                auto_in_a_valid,
  input  [2:0]  auto_in_a_bits_opcode,
                auto_in_a_bits_param,
  input  [1:0]  auto_in_a_bits_size,
  input  [10:0] auto_in_a_bits_source,
  input  [16:0] auto_in_a_bits_address,
  input  [7:0]  auto_in_a_bits_mask,
  input         auto_in_a_bits_corrupt,
                auto_in_d_ready,
  output        auto_in_a_ready,
                auto_in_d_valid,
  output [1:0]  auto_in_d_bits_size,
  output [10:0] auto_in_d_bits_source,
  output [63:0] auto_in_d_bits_data
);

  wire [63:0] _GEN_86 =
    auto_in_a_bits_address[11:3] == 9'h56
      ? 64'h300000000000000
      : auto_in_a_bits_address[11:3] == 9'h55
          ? 64'hB200000004000000
          : auto_in_a_bits_address[11:3] == 9'h54
              ? 64'h300000000757063
              : auto_in_a_bits_address[11:3] == 9'h53
                  ? 64'hA600000004000000
                  : auto_in_a_bits_address[11:3] == 9'h52
                      ? 64'h300000020000000
                      : auto_in_a_bits_address[11:3] == 9'h51
                          ? 64'h9B00000004000000
                          : auto_in_a_bits_address[11:3] == 9'h50
                              ? 64'h300000001000000
                              : auto_in_a_bits_address[11:3] == 9'h4F
                                  ? 64'h9000000004000000
                                  : auto_in_a_bits_address[11:3] == 9'h4E
                                      ? 64'h300000000800000
                                      : auto_in_a_bits_address[11:3] == 9'h4D
                                          ? 64'h8300000004000000
                                          : auto_in_a_bits_address[11:3] == 9'h4C
                                              ? 64'h300000040000000
                                              : auto_in_a_bits_address[11:3] == 9'h4B
                                                  ? 64'h7600000004000000
                                                  : auto_in_a_bits_address[11:3] == 9'h4A
                                                      ? 64'h300000040000000
                                                      : auto_in_a_bits_address[11:3] == 9'h49
                                                          ? 64'h6300000004000000
                                                          : auto_in_a_bits_address[11:3] == 9'h48
                                                              ? 64'h300000000766373
                                                              : auto_in_a_bits_address[11:3] == 9'h47
                                                                  ? 64'h697200306D6F6F62
                                                                  : auto_in_a_bits_address[11:3] == 9'h46
                                                                      ? 64'h2C7261622D626375
                                                                      : auto_in_a_bits_address[11:3] == 9'h45
                                                                          ? 64'h1B00000014000000
                                                                          : auto_in_a_bits_address[11:3] == 9'h44
                                                                              ? 64'h300000000000000
                                                                              : auto_in_a_bits_address[11:3] == 9'h43
                                                                                  ? 64'h5300000004000000
                                                                                  : auto_in_a_bits_address[11:3] == 9'h42
                                                                                      ? 64'h300000000000030
                                                                                      : auto_in_a_bits_address[11:3] == 9'h41
                                                                                          ? 64'h4075706301000000
                                                                                          : auto_in_a_bits_address[11:3] == 9'h40
                                                                                              ? 64'h40420F0040000000
                                                                                              : auto_in_a_bits_address[11:3] == 9'h3F
                                                                                                  ? 64'h400000003000000
                                                                                                  : auto_in_a_bits_address[11:3] == 9'h3E
                                                                                                      ? 64'hF000000
                                                                                                      : auto_in_a_bits_address[11:3] == 9'h3D
                                                                                                          ? 64'h400000003000000
                                                                                                          : auto_in_a_bits_address[11:3] == 9'h3C
                                                                                                              ? 64'h100000000000000
                                                                                                              : auto_in_a_bits_address[11:3] == 9'h3B
                                                                                                                  ? 64'h400000003000000
                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h3A
                                                                                                                      ? 64'h73757063
                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h39
                                                                                                                          ? 64'h100000002000000
                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h38
                                                                                                                              ? 64'h30303030
                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h37
                                                                                                                                  ? 64'h32303031406C6169
                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h36
                                                                                                                                      ? 64'h7265732F636F732F
                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h35
                                                                                                                                          ? 64'h3400000015000000
                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h34
                                                                                                                                              ? 64'h300000000006E65
                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h33
                                                                                                                                                  ? 64'h736F686301000000
                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h32
                                                                                                                                                      ? 64'h200000000000000
                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h31
                                                                                                                                                          ? 64'h3030303032303031
                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h30
                                                                                                                                                              ? 64'h406C61697265732F
                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h2F
                                                                                                                                                                  ? 64'h636F732F2C000000
                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h2E
                                                                                                                                                                      ? 64'h1500000003000000
                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h2D
                                                                                                                                                                          ? 64'h73657361696C61
                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h2C
                                                                                                                                                                              ? 64'h100000000000000
                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h2B
                                                                                                                                                                                  ? 64'h6472617970696863
                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h2A
                                                                                                                                                                                      ? 64'h2C7261622D626375
                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h29
                                                                                                                                                                                          ? 64'h2600000011000000
                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h28
                                                                                                                                                                                              ? 64'h300000000000000
                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h27
                                                                                                                                                                                                  ? 64'h7665642D64726179
                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h26
                                                                                                                                                                                                      ? 64'h706968632C726162
                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h25
                                                                                                                                                                                                          ? 64'h2D6263751B000000
                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h24
                                                                                                                                                                                                              ? 64'h1500000003000000
                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h23
                                                                                                                                                                                                                  ? 64'h10000000F000000
                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h22
                                                                                                                                                                                                                      ? 64'h400000003000000
                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h21
                                                                                                                                                                                                                          ? 64'h100000000000000
                                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h20
                                                                                                                                                                                                                              ? 64'h400000003000000
                                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h1F ? 64'h1000000 : auto_in_a_bits_address[11:3] == 9'h1E | auto_in_a_bits_address[11:3] == 9'h1D ? 64'h0 : auto_in_a_bits_address[11:3] == 9'h1C ? 64'hF409000060020000 : auto_in_a_bits_address[11:3] == 9'h1B ? 64'h10000000 : auto_in_a_bits_address[11:3] == 9'h1A ? 64'h1100000028000000 : auto_in_a_bits_address[11:3] == 9'h19 ? 64'h2C0A000038000000 : auto_in_a_bits_address[11:3] == 9'h18 ? 64'h8C0C0000EDFE0DD0 : auto_in_a_bits_address[11:3] == 9'h17 ? 64'h1330200073 : auto_in_a_bits_address[11:3] == 9'h16 ? 64'h3006307308000613 : auto_in_a_bits_address[11:3] == 9'h15 ? 64'h185859300000597 : auto_in_a_bits_address[11:3] == 9'h14 ? 64'hF140257334151073 : auto_in_a_bits_address[11:3] == 9'h13 ? 64'h5350300004537 : auto_in_a_bits_address[11:3] == 9'h12 ? 64'h5A02300B505B3 : auto_in_a_bits_address[11:3] == 9'h11 ? 64'h251513FE029EE3 : auto_in_a_bits_address[11:3] == 9'h10 ? 64'h5A283FC1FF06F : auto_in_a_bits_address[11:3] == 9'hF ? 64'h0 : auto_in_a_bits_address[11:3] == 9'hE ? 64'hFFDFF06F : auto_in_a_bits_address[11:3] == 9'hD ? 64'h1050007330052073 : auto_in_a_bits_address[11:3] == 9'hC ? 64'h3045107300800513 : auto_in_a_bits_address[11:3] == 9'hB ? 64'h3030107300028463 : auto_in_a_bits_address[11:3] == 9'hA ? 64'h12F2934122D293 : auto_in_a_bits_address[11:3] == 9'h9 ? 64'h301022F330551073 : auto_in_a_bits_address[11:3] == 9'h8 ? 64'hFC05051300000517 : auto_in_a_bits_address[11:3] == 9'h7 | auto_in_a_bits_address[11:3] == 9'h6 ? 64'h0 : auto_in_a_bits_address[11:3] == 9'h5 ? 64'h6C0006F : auto_in_a_bits_address[11:3] == 9'h4 ? 64'hFE069AE3FFC62683 : auto_in_a_bits_address[11:3] == 9'h3 ? 64'h46061300D62023 : auto_in_a_bits_address[11:3] == 9'h2 ? 64'h10069300458613 : auto_in_a_bits_address[11:3] == 9'h1 ? 64'h780006F00050463 : 64'hF1402573020005B7;
  wire [63:0] _GEN_172 =
    auto_in_a_bits_address[11:3] == 9'hAC
      ? 64'h30303030
      : auto_in_a_bits_address[11:3] == 9'hAB
          ? 64'h3130324072656C6C
          : auto_in_a_bits_address[11:3] == 9'hAA
              ? 64'h6F72746E6F632D65
              : auto_in_a_bits_address[11:3] == 9'hA9
                  ? 64'h6863616301000000
                  : auto_in_a_bits_address[11:3] == 9'hA8
                      ? 64'h2000000006C6F72
                      : auto_in_a_bits_address[11:3] == 9'hA7
                          ? 64'h746E6F63A8010000
                          : auto_in_a_bits_address[11:3] == 9'hA6
                              ? 64'h800000003000000
                              : auto_in_a_bits_address[11:3] == 9'hA5
                                  ? 64'h10000000400000
                                  : auto_in_a_bits_address[11:3] == 9'hA4
                                      ? 64'h2E01000008000000
                                      : auto_in_a_bits_address[11:3] == 9'hA3
                                          ? 64'h300000000000030
                                          : auto_in_a_bits_address[11:3] == 9'hA2
                                              ? 64'h303034406765722D
                                              : auto_in_a_bits_address[11:3] == 9'hA1
                                                  ? 64'h737365726464612D
                                                  : auto_in_a_bits_address[11:3] == 9'hA0
                                                      ? 64'h746F6F6201000000
                                                      : auto_in_a_bits_address[11:3] == 9'h9F
                                                          ? 64'hA101000000000000
                                                          : auto_in_a_bits_address[11:3] == 9'h9E
                                                              ? 64'h300000000737562
                                                              : auto_in_a_bits_address[11:3] == 9'h9D
                                                                  ? 64'h2D656C706D697300
                                                                  : auto_in_a_bits_address[11:3] == 9'h9C
                                                                      ? 64'h636F732D64726179
                                                                      : auto_in_a_bits_address[11:3] == 9'h9B
                                                                          ? 64'h706968632C726162
                                                                          : auto_in_a_bits_address[11:3] == 9'h9A
                                                                              ? 64'h2D6263751B000000
                                                                              : auto_in_a_bits_address[11:3] == 9'h99
                                                                                  ? 64'h2000000003000000
                                                                                  : auto_in_a_bits_address[11:3] == 9'h98
                                                                                      ? 64'h10000000F000000
                                                                                      : auto_in_a_bits_address[11:3] == 9'h97
                                                                                          ? 64'h400000003000000
                                                                                          : auto_in_a_bits_address[11:3] == 9'h96
                                                                                              ? 64'h100000000000000
                                                                                              : auto_in_a_bits_address[11:3] == 9'h95
                                                                                                  ? 64'h400000003000000
                                                                                                  : auto_in_a_bits_address[11:3] == 9'h94
                                                                                                      ? 64'h636F7301000000
                                                                                                      : auto_in_a_bits_address[11:3] == 9'h93
                                                                                                          ? 64'h200000002000000
                                                                                                          : auto_in_a_bits_address[11:3] == 9'h92
                                                                                                              ? 64'h9901000004000000
                                                                                                              : auto_in_a_bits_address[11:3] == 9'h91
                                                                                                                  ? 64'h300000000000010
                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h90
                                                                                                                      ? 64'h802E010000
                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h8F
                                                                                                                          ? 64'h800000003000000
                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h8E
                                                                                                                              ? 64'h79726F6D656D
                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h8D
                                                                                                                                  ? 64'hA600000007000000
                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h8C
                                                                                                                                      ? 64'h300000000303030
                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h8B
                                                                                                                                          ? 64'h3030303038407972
                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h8A
                                                                                                                                              ? 64'h6F6D656D01000000
                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h89
                                                                                                                                                  ? 64'h200000000000030
                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h88
                                                                                                                                                      ? 64'h666974682C626375
                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h87
                                                                                                                                                          ? 64'h1B0000000A000000
                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h86
                                                                                                                                                              ? 64'h300000000000000
                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h85
                                                                                                                                                                  ? 64'h6669746801000000
                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h84
                                                                                                                                                                      ? 64'h200000002000000
                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h83
                                                                                                                                                                          ? 64'h200000003000000
                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h82
                                                                                                                                                                              ? 64'h9901000004000000
                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h81
                                                                                                                                                                                  ? 64'h300000084010000
                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h80
                                                                                                                                                                                      ? 64'h3000000
                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h7F
                                                                                                                                                                                          ? 64'h63746E692D75
                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h7E
                                                                                                                                                                                              ? 64'h70632C7663736972
                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h7D
                                                                                                                                                                                                  ? 64'h1B0000000F000000
                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h7C
                                                                                                                                                                                                      ? 64'h300000001000000
                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h7B
                                                                                                                                                                                                          ? 64'h7301000004000000
                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h7A
                                                                                                                                                                                                              ? 64'h300000000000000
                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h79
                                                                                                                                                                                                                  ? 64'h72656C6C6F72746E
                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h78
                                                                                                                                                                                                                      ? 64'h6F632D7470757272
                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h77
                                                                                                                                                                                                                          ? 64'h65746E6901000000
                                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h76
                                                                                                                                                                                                                              ? 64'h6901000000000000
                                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h75
                                                                                                                                                                                                                                  ? 64'h300000040420F00
                                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h74
                                                                                                                                                                                                                                      ? 64'h4000000004000000
                                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h73 ? 64'h300000000000000 : auto_in_a_bits_address[11:3] == 9'h72 ? 64'h79616B6F62010000 : auto_in_a_bits_address[11:3] == 9'h71 ? 64'h500000003000000 : auto_in_a_bits_address[11:3] == 9'h70 ? 64'h800000051010000 : auto_in_a_bits_address[11:3] == 9'h6F ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'h6E ? 64'h40000003C010000 : auto_in_a_bits_address[11:3] == 9'h6D ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'h6C ? 64'h6D7068697A5F : auto_in_a_bits_address[11:3] == 9'h6B ? 64'h6965636E6566697A : auto_in_a_bits_address[11:3] == 9'h6A ? 64'h5F727363697A6364 : auto_in_a_bits_address[11:3] == 9'h69 ? 64'h66616D6934367672 : auto_in_a_bits_address[11:3] == 9'h68 ? 64'h320100001F000000 : auto_in_a_bits_address[11:3] == 9'h67 ? 64'h300000000000000 : auto_in_a_bits_address[11:3] == 9'h66 ? 64'h2E01000004000000 : auto_in_a_bits_address[11:3] == 9'h65 ? 64'h300000001000000 : auto_in_a_bits_address[11:3] == 9'h64 ? 64'h1D01000004000000 : auto_in_a_bits_address[11:3] == 9'h63 ? 64'h300000000003933 : auto_in_a_bits_address[11:3] == 9'h62 ? 64'h76732C7663736972 : auto_in_a_bits_address[11:3] == 9'h61 ? 64'h140100000B000000 : auto_in_a_bits_address[11:3] == 9'h60 ? 64'h300000020000000 : auto_in_a_bits_address[11:3] == 9'h5F ? 64'h901000004000000 : auto_in_a_bits_address[11:3] == 9'h5E ? 64'h300000001000000 : auto_in_a_bits_address[11:3] == 9'h5D ? 64'hFE00000004000000 : auto_in_a_bits_address[11:3] == 9'h5C ? 64'h300000000800000 : auto_in_a_bits_address[11:3] == 9'h5B ? 64'hF100000004000000 : auto_in_a_bits_address[11:3] == 9'h5A ? 64'h300000040000000 : auto_in_a_bits_address[11:3] == 9'h59 ? 64'hE400000004000000 : auto_in_a_bits_address[11:3] == 9'h58 ? 64'h300000040000000 : auto_in_a_bits_address[11:3] == 9'h57 ? 64'hD100000004000000 : _GEN_86;
  wire [63:0] _GEN_258 =
    auto_in_a_bits_address[11:3] == 9'h102
      ? 64'h300000001000000
      : auto_in_a_bits_address[11:3] == 9'h101
          ? 64'h7301000004000000
          : auto_in_a_bits_address[11:3] == 9'h100
              ? 64'h300000000000000
              : auto_in_a_bits_address[11:3] == 9'hFF
                  ? 64'h3030303030306340
                  : auto_in_a_bits_address[11:3] == 9'hFE
                      ? 64'h72656C6C6F72746E
                      : auto_in_a_bits_address[11:3] == 9'hFD
                          ? 64'h6F632D7470757272
                          : auto_in_a_bits_address[11:3] == 9'hFC
                              ? 64'h65746E6901000000
                              : auto_in_a_bits_address[11:3] == 9'hFB
                                  ? 64'h200000000100000
                                  : auto_in_a_bits_address[11:3] == 9'hFA
                                      ? 64'h3000002E010000
                                      : auto_in_a_bits_address[11:3] == 9'hF9
                                          ? 64'h800000003000000
                                          : auto_in_a_bits_address[11:3] == 9'hF8
                                              ? 64'h30726F7272
                                              : auto_in_a_bits_address[11:3] == 9'hF7
                                                  ? 64'h652C657669666973
                                                  : auto_in_a_bits_address[11:3] == 9'hF6
                                                      ? 64'h1B0000000E000000
                                                      : auto_in_a_bits_address[11:3] == 9'hF5
                                                          ? 64'h300000000000030
                                                          : auto_in_a_bits_address[11:3] == 9'hF4
                                                              ? 64'h3030334065636976
                                                              : auto_in_a_bits_address[11:3] == 9'hF3
                                                                  ? 64'h65642D726F727265
                                                                  : auto_in_a_bits_address[11:3] == 9'hF2
                                                                      ? 64'h100000002000000
                                                                      : auto_in_a_bits_address[11:3] == 9'hF1
                                                                          ? 64'h6C6F72746E6F63
                                                                          : auto_in_a_bits_address[11:3] == 9'hF0
                                                                              ? 64'hA801000008000000
                                                                              : auto_in_a_bits_address[11:3] == 9'hEF
                                                                                  ? 64'h300000000100000
                                                                                  : auto_in_a_bits_address[11:3] == 9'hEE
                                                                                      ? 64'h2E010000
                                                                                      : auto_in_a_bits_address[11:3] == 9'hED
                                                                                          ? 64'h800000003000000
                                                                                          : auto_in_a_bits_address[11:3] == 9'hEC
                                                                                              ? 64'hFFFF000003000000
                                                                                              : auto_in_a_bits_address[11:3] == 9'hEB
                                                                                                  ? 64'hDE01000008000000
                                                                                                  : auto_in_a_bits_address[11:3] == 9'hEA
                                                                                                      ? 64'h300000000000000
                                                                                                      : auto_in_a_bits_address[11:3] == 9'hE9
                                                                                                          ? 64'h6761746AF2010000
                                                                                                          : auto_in_a_bits_address[11:3] == 9'hE8
                                                                                                              ? 64'h500000003000000
                                                                                                              : auto_in_a_bits_address[11:3] == 9'hE7
                                                                                                                  ? 64'h3331302D
                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hE6
                                                                                                                      ? 64'h67756265642C7663
                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hE5
                                                                                                                          ? 64'h736972003331302D
                                                                                                                          : auto_in_a_bits_address[11:3] == 9'hE4
                                                                                                                              ? 64'h67756265642C6576
                                                                                                                              : auto_in_a_bits_address[11:3] == 9'hE3
                                                                                                                                  ? 64'h696669731B000000
                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hE2
                                                                                                                                      ? 64'h2100000003000000
                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hE1
                                                                                                                                          ? 64'h304072656C6C
                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'hE0
                                                                                                                                              ? 64'h6F72746E6F632D67
                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'hDF
                                                                                                                                                  ? 64'h7562656401000000
                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hDE
                                                                                                                                                      ? 64'h2000000006C6F72
                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hDD
                                                                                                                                                          ? 64'h746E6F63A8010000
                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'hDC
                                                                                                                                                              ? 64'h800000003000000
                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'hDB
                                                                                                                                                                  ? 64'h10000000001000
                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hDA
                                                                                                                                                                      ? 64'h2E01000008000000
                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hD9
                                                                                                                                                                          ? 64'h300000000003030
                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'hD8
                                                                                                                                                                              ? 64'h3030303140726574
                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'hD7
                                                                                                                                                                                  ? 64'h61672D6B636F6C63
                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hD6
                                                                                                                                                                                      ? 64'h100000002000000
                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hD5
                                                                                                                                                                                          ? 64'h6C6F72746E6F63
                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'hD4
                                                                                                                                                                                              ? 64'hA801000008000000
                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'hD3
                                                                                                                                                                                                  ? 64'h300000000000100
                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hD2
                                                                                                                                                                                                      ? 64'h22E010000
                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hD1
                                                                                                                                                                                                          ? 64'h800000003000000
                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'hD0
                                                                                                                                                                                                              ? 64'h700000003000000
                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'hCF
                                                                                                                                                                                                                  ? 64'h300000003000000
                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hCE
                                                                                                                                                                                                                      ? 64'hDE01000010000000
                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hCD
                                                                                                                                                                                                                          ? 64'h300000000000000
                                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'hCC
                                                                                                                                                                                                                              ? 64'h30746E696C632C76
                                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'hCB
                                                                                                                                                                                                                                  ? 64'h637369721B000000
                                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'hCA
                                                                                                                                                                                                                                      ? 64'hD00000003000000
                                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'hC9 ? 64'h3030303030 : auto_in_a_bits_address[11:3] == 9'hC8 ? 64'h303240746E696C63 : auto_in_a_bits_address[11:3] == 9'hC7 ? 64'h100000002000000 : auto_in_a_bits_address[11:3] == 9'hC6 ? 64'h100000099010000 : auto_in_a_bits_address[11:3] == 9'hC5 ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'hC4 ? 64'hC000000CC010000 : auto_in_a_bits_address[11:3] == 9'hC3 ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'hC2 ? 64'h6C6F72746E6F63 : auto_in_a_bits_address[11:3] == 9'hC1 ? 64'hA801000008000000 : auto_in_a_bits_address[11:3] == 9'hC0 ? 64'h300000000100000 : auto_in_a_bits_address[11:3] == 9'hBF ? 64'h1022E010000 : auto_in_a_bits_address[11:3] == 9'hBE ? 64'h800000003000000 : auto_in_a_bits_address[11:3] == 9'hBD ? 64'h20000001D010000 : auto_in_a_bits_address[11:3] == 9'hBC ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'hBB ? 64'h65686361 : auto_in_a_bits_address[11:3] == 9'hBA ? 64'h6300306568636163 : auto_in_a_bits_address[11:3] == 9'hB9 ? 64'h65766973756C636E : auto_in_a_bits_address[11:3] == 9'hB8 ? 64'h692C657669666973 : auto_in_a_bits_address[11:3] == 9'hB7 ? 64'h1B0000001D000000 : auto_in_a_bits_address[11:3] == 9'hB6 ? 64'h3000000BE010000 : auto_in_a_bits_address[11:3] == 9'hB5 ? 64'h3000000 : auto_in_a_bits_address[11:3] == 9'hB4 ? 64'h80085000000 : auto_in_a_bits_address[11:3] == 9'hB3 ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'hB2 ? 64'h4000078000000 : auto_in_a_bits_address[11:3] == 9'hB1 ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'hB0 ? 64'h2000000B2010000 : auto_in_a_bits_address[11:3] == 9'hAF ? 64'h400000003000000 : auto_in_a_bits_address[11:3] == 9'hAE ? 64'h4000000065000000 : auto_in_a_bits_address[11:3] == 9'hAD ? 64'h400000003000000 : _GEN_172;
  wire [63:0] _GEN_344 =
    auto_in_a_bits_address[11:3] == 9'h158
      ? 64'h10000000001100
      : auto_in_a_bits_address[11:3] == 9'h157
          ? 64'h2E01000008000000
          : auto_in_a_bits_address[11:3] == 9'h156
              ? 64'h300000000000000
              : auto_in_a_bits_address[11:3] == 9'h155
                  ? 64'h3030303031314072
                  : auto_in_a_bits_address[11:3] == 9'h154
                      ? 64'h65747465732D7465
                      : auto_in_a_bits_address[11:3] == 9'h153
                          ? 64'h7365722D656C6974
                          : auto_in_a_bits_address[11:3] == 9'h152
                              ? 64'h100000002000000
                              : auto_in_a_bits_address[11:3] == 9'h151
                                  ? 64'h400000099010000
                                  : auto_in_a_bits_address[11:3] == 9'h150
                                      ? 64'h400000003000000
                                      : auto_in_a_bits_address[11:3] == 9'h14F
                                          ? 64'h6B636F6C632D64
                                          : auto_in_a_bits_address[11:3] == 9'h14E
                                              ? 64'h657869661B000000
                                              : auto_in_a_bits_address[11:3] == 9'h14D
                                                  ? 64'hC00000003000000
                                                  : auto_in_a_bits_address[11:3] == 9'h14C
                                                      ? 64'h6B636F6C
                                                      : auto_in_a_bits_address[11:3] == 9'h14B
                                                          ? 64'h635F737562705F6D
                                                          : auto_in_a_bits_address[11:3] == 9'h14A
                                                              ? 64'h6574737973627573
                                                              : auto_in_a_bits_address[11:3] == 9'h149
                                                                  ? 64'h4D02000015000000
                                                                  : auto_in_a_bits_address[11:3] == 9'h148
                                                                      ? 64'h30000000065CD1D
                                                                      : auto_in_a_bits_address[11:3] == 9'h147
                                                                          ? 64'h5300000004000000
                                                                          : auto_in_a_bits_address[11:3] == 9'h146
                                                                              ? 64'h300000000000000
                                                                              : auto_in_a_bits_address[11:3] == 9'h145
                                                                                  ? 64'h4002000004000000
                                                                                  : auto_in_a_bits_address[11:3] == 9'h144
                                                                                      ? 64'h300000000000000
                                                                                      : auto_in_a_bits_address[11:3] == 9'h143
                                                                                          ? 64'h6B636F6C635F7375
                                                                                          : auto_in_a_bits_address[11:3] == 9'h142
                                                                                              ? 64'h62705F6D65747379
                                                                                              : auto_in_a_bits_address[11:3] == 9'h141
                                                                                                  ? 64'h7362757301000000
                                                                                                  : auto_in_a_bits_address[11:3] == 9'h140
                                                                                                      ? 64'h2000000006B636F
                                                                                                      : auto_in_a_bits_address[11:3] == 9'h13F
                                                                                                          ? 64'h6C632D6465786966
                                                                                                          : auto_in_a_bits_address[11:3] == 9'h13E
                                                                                                              ? 64'h1B0000000C000000
                                                                                                              : auto_in_a_bits_address[11:3] == 9'h13D
                                                                                                                  ? 64'h300000000000000
                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h13C
                                                                                                                      ? 64'h6B636F6C635F7375
                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h13B
                                                                                                                          ? 64'h626D5F6D65747379
                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h13A
                                                                                                                              ? 64'h736275734D020000
                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h139
                                                                                                                                  ? 64'h1500000003000000
                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h138
                                                                                                                                      ? 64'h65CD1D53000000
                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h137
                                                                                                                                          ? 64'h400000003000000
                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h136
                                                                                                                                              ? 64'h40020000
                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h135
                                                                                                                                                  ? 64'h400000003000000
                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h134
                                                                                                                                                      ? 64'h6B636F6C
                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h133
                                                                                                                                                          ? 64'h635F7375626D5F6D
                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h132
                                                                                                                                                              ? 64'h6574737973627573
                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h131
                                                                                                                                                                  ? 64'h100000002000000
                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h130
                                                                                                                                                                      ? 64'h6C6F72746E6F63
                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h12F
                                                                                                                                                                          ? 64'hA801000008000000
                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h12E
                                                                                                                                                                              ? 64'h300000000100000
                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h12D
                                                                                                                                                                                  ? 64'h2102E010000
                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h12C
                                                                                                                                                                                      ? 64'h800000003000000
                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h12B
                                                                                                                                                                                          ? 64'h100000035020000
                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h12A
                                                                                                                                                                                              ? 64'h400000003000000
                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h129
                                                                                                                                                                                                  ? 64'h500000024020000
                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h128
                                                                                                                                                                                                      ? 64'h400000003000000
                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h127
                                                                                                                                                                                                          ? 64'h30747261
                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h126
                                                                                                                                                                                                              ? 64'h752C657669666973
                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h125
                                                                                                                                                                                                                  ? 64'h1B0000000D000000
                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h124
                                                                                                                                                                                                                      ? 64'h300000004000000
                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h123
                                                                                                                                                                                                                          ? 64'h1D02000004000000
                                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h122
                                                                                                                                                                                                                              ? 64'h300000000303030
                                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h121
                                                                                                                                                                                                                                  ? 64'h3032303031406C61
                                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h120
                                                                                                                                                                                                                                      ? 64'h6972657301000000
                                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h11F
                                                                                                                                                                                                                                          ? 64'h2000000006D656D
                                                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h11E ? 64'hA801000004000000 : auto_in_a_bits_address[11:3] == 9'h11D ? 64'h300000000000100 : auto_in_a_bits_address[11:3] == 9'h11C ? 64'h1002E010000 : auto_in_a_bits_address[11:3] == 9'h11B ? 64'h800000003000000 : auto_in_a_bits_address[11:3] == 9'h11A ? 64'h306D6F722C6576 : auto_in_a_bits_address[11:3] == 9'h119 ? 64'h696669731B000000 : auto_in_a_bits_address[11:3] == 9'h118 ? 64'hC00000003000000 : auto_in_a_bits_address[11:3] == 9'h117 ? 64'h3030303031 : auto_in_a_bits_address[11:3] == 9'h116 ? 64'h406D6F7201000000 : auto_in_a_bits_address[11:3] == 9'h115 ? 64'h200000005000000 : auto_in_a_bits_address[11:3] == 9'h114 ? 64'h9901000004000000 : auto_in_a_bits_address[11:3] == 9'h113 ? 64'h300000001000000 : auto_in_a_bits_address[11:3] == 9'h112 ? 64'h1202000004000000 : auto_in_a_bits_address[11:3] == 9'h111 ? 64'h300000001000000 : auto_in_a_bits_address[11:3] == 9'h110 ? 64'hFF01000004000000 : auto_in_a_bits_address[11:3] == 9'h10F ? 64'h3000000006C6F72 : auto_in_a_bits_address[11:3] == 9'h10E ? 64'h746E6F63A8010000 : auto_in_a_bits_address[11:3] == 9'h10D ? 64'h800000003000000 : auto_in_a_bits_address[11:3] == 9'h10C ? 64'h40000000C : auto_in_a_bits_address[11:3] == 9'h10B ? 64'h2E01000008000000 : auto_in_a_bits_address[11:3] == 9'h10A ? 64'h300000009000000 : auto_in_a_bits_address[11:3] == 9'h109 ? 64'h30000000B000000 : auto_in_a_bits_address[11:3] == 9'h108 ? 64'h3000000DE010000 : auto_in_a_bits_address[11:3] == 9'h107 ? 64'h1000000003000000 : auto_in_a_bits_address[11:3] == 9'h106 ? 64'h8401000000000000 : auto_in_a_bits_address[11:3] == 9'h105 ? 64'h300000000306369 : auto_in_a_bits_address[11:3] == 9'h104 ? 64'h6C702C7663736972 : auto_in_a_bits_address[11:3] == 9'h103 ? 64'h1B0000000C000000 : _GEN_258;
  plusarg_reader #(
    .DEFAULT(0),
    .FORMAT("tilelink_timeout=%d"),
    .WIDTH(32)
  ) plusarg_reader_1 (
    .out (/* unused */)
  );
  assign auto_in_a_ready = auto_in_d_ready;
  assign auto_in_d_valid = auto_in_a_valid;
  assign auto_in_d_bits_size = auto_in_a_bits_size;
  assign auto_in_d_bits_source = auto_in_a_bits_source;
  assign auto_in_d_bits_data =
    (|(auto_in_a_bits_address[15:12])) | (&(auto_in_a_bits_address[11:3])) | auto_in_a_bits_address[11:3] == 9'h1FE | auto_in_a_bits_address[11:3] == 9'h1FD | auto_in_a_bits_address[11:3] == 9'h1FC | auto_in_a_bits_address[11:3] == 9'h1FB | auto_in_a_bits_address[11:3] == 9'h1FA | auto_in_a_bits_address[11:3] == 9'h1F9 | auto_in_a_bits_address[11:3] == 9'h1F8 | auto_in_a_bits_address[11:3] == 9'h1F7 | auto_in_a_bits_address[11:3] == 9'h1F6 | auto_in_a_bits_address[11:3] == 9'h1F5 | auto_in_a_bits_address[11:3] == 9'h1F4 | auto_in_a_bits_address[11:3] == 9'h1F3 | auto_in_a_bits_address[11:3] == 9'h1F2 | auto_in_a_bits_address[11:3] == 9'h1F1 | auto_in_a_bits_address[11:3] == 9'h1F0 | auto_in_a_bits_address[11:3] == 9'h1EF | auto_in_a_bits_address[11:3] == 9'h1EE | auto_in_a_bits_address[11:3] == 9'h1ED | auto_in_a_bits_address[11:3] == 9'h1EC | auto_in_a_bits_address[11:3] == 9'h1EB | auto_in_a_bits_address[11:3] == 9'h1EA | auto_in_a_bits_address[11:3] == 9'h1E9 | auto_in_a_bits_address[11:3] == 9'h1E8 | auto_in_a_bits_address[11:3] == 9'h1E7 | auto_in_a_bits_address[11:3] == 9'h1E6 | auto_in_a_bits_address[11:3] == 9'h1E5 | auto_in_a_bits_address[11:3] == 9'h1E4 | auto_in_a_bits_address[11:3] == 9'h1E3 | auto_in_a_bits_address[11:3] == 9'h1E2 | auto_in_a_bits_address[11:3] == 9'h1E1 | auto_in_a_bits_address[11:3] == 9'h1E0 | auto_in_a_bits_address[11:3] == 9'h1DF | auto_in_a_bits_address[11:3] == 9'h1DE | auto_in_a_bits_address[11:3] == 9'h1DD | auto_in_a_bits_address[11:3] == 9'h1DC | auto_in_a_bits_address[11:3] == 9'h1DB | auto_in_a_bits_address[11:3] == 9'h1DA | auto_in_a_bits_address[11:3] == 9'h1D9 | auto_in_a_bits_address[11:3] == 9'h1D8 | auto_in_a_bits_address[11:3] == 9'h1D7 | auto_in_a_bits_address[11:3] == 9'h1D6 | auto_in_a_bits_address[11:3] == 9'h1D5 | auto_in_a_bits_address[11:3] == 9'h1D4 | auto_in_a_bits_address[11:3] == 9'h1D3 | auto_in_a_bits_address[11:3] == 9'h1D2 | auto_in_a_bits_address[11:3] == 9'h1D1 | auto_in_a_bits_address[11:3] == 9'h1D0 | auto_in_a_bits_address[11:3] == 9'h1CF
    | auto_in_a_bits_address[11:3] == 9'h1CE | auto_in_a_bits_address[11:3] == 9'h1CD | auto_in_a_bits_address[11:3] == 9'h1CC | auto_in_a_bits_address[11:3] == 9'h1CB | auto_in_a_bits_address[11:3] == 9'h1CA | auto_in_a_bits_address[11:3] == 9'h1C9 | auto_in_a_bits_address[11:3] == 9'h1C8 | auto_in_a_bits_address[11:3] == 9'h1C7 | auto_in_a_bits_address[11:3] == 9'h1C6 | auto_in_a_bits_address[11:3] == 9'h1C5 | auto_in_a_bits_address[11:3] == 9'h1C4 | auto_in_a_bits_address[11:3] == 9'h1C3 | auto_in_a_bits_address[11:3] == 9'h1C2 | auto_in_a_bits_address[11:3] == 9'h1C1 | auto_in_a_bits_address[11:3] == 9'h1C0 | auto_in_a_bits_address[11:3] == 9'h1BF | auto_in_a_bits_address[11:3] == 9'h1BE | auto_in_a_bits_address[11:3] == 9'h1BD | auto_in_a_bits_address[11:3] == 9'h1BC | auto_in_a_bits_address[11:3] == 9'h1BB | auto_in_a_bits_address[11:3] == 9'h1BA | auto_in_a_bits_address[11:3] == 9'h1B9 | auto_in_a_bits_address[11:3] == 9'h1B8 | auto_in_a_bits_address[11:3] == 9'h1B7 | auto_in_a_bits_address[11:3] == 9'h1B6 | auto_in_a_bits_address[11:3] == 9'h1B5 | auto_in_a_bits_address[11:3] == 9'h1B4 | auto_in_a_bits_address[11:3] == 9'h1B3 | auto_in_a_bits_address[11:3] == 9'h1B2 | auto_in_a_bits_address[11:3] == 9'h1B1 | auto_in_a_bits_address[11:3] == 9'h1B0 | auto_in_a_bits_address[11:3] == 9'h1AF | auto_in_a_bits_address[11:3] == 9'h1AE | auto_in_a_bits_address[11:3] == 9'h1AD | auto_in_a_bits_address[11:3] == 9'h1AC | auto_in_a_bits_address[11:3] == 9'h1AB | auto_in_a_bits_address[11:3] == 9'h1AA
      ? 64'h0
      : auto_in_a_bits_address[11:3] == 9'h1A9
          ? 64'h73656D
          : auto_in_a_bits_address[11:3] == 9'h1A8
              ? 64'h616E2D7475707475
              : auto_in_a_bits_address[11:3] == 9'h1A7
                  ? 64'h6F2D6B636F6C6300
                  : auto_in_a_bits_address[11:3] == 9'h1A6
                      ? 64'h736C6C65632D6B63
                      : auto_in_a_bits_address[11:3] == 9'h1A5
                          ? 64'h6F6C632300737470
                          : auto_in_a_bits_address[11:3] == 9'h1A4
                              ? 64'h75727265746E6900
                              : auto_in_a_bits_address[11:3] == 9'h1A3
                                  ? 64'h746E657261702D74
                                  : auto_in_a_bits_address[11:3] == 9'h1A2
                                      ? 64'h7075727265746E69
                                      : auto_in_a_bits_address[11:3] == 9'h1A1
                                          ? 64'h736B636F6C6300
                                          : auto_in_a_bits_address[11:3] == 9'h1A0
                                              ? 64'h7665646E2C766373
                                              : auto_in_a_bits_address[11:3] == 9'h19F
                                                  ? 64'h697200797469726F
                                                  : auto_in_a_bits_address[11:3] == 9'h19E
                                                      ? 64'h6972702D78616D2C
                                                      : auto_in_a_bits_address[11:3] == 9'h19D
                                                          ? 64'h7663736972006863
                                                          : auto_in_a_bits_address[11:3] == 9'h19C
                                                              ? 64'h617474612D677562
                                                              : auto_in_a_bits_address[11:3] == 9'h19B
                                                                  ? 64'h6564006465646E65
                                                                  : auto_in_a_bits_address[11:3] == 9'h19A
                                                                      ? 64'h7478652D73747075
                                                                      : auto_in_a_bits_address[11:3] == 9'h199
                                                                          ? 64'h727265746E690074
                                                                          : auto_in_a_bits_address[11:3] == 9'h198
                                                                              ? 64'h6E756F632D726873
                                                                              : auto_in_a_bits_address[11:3] == 9'h197
                                                                                  ? 64'h6D2C657669666973
                                                                                  : auto_in_a_bits_address[11:3] == 9'h196
                                                                                      ? 64'h64656966696E75
                                                                                      : auto_in_a_bits_address[11:3] == 9'h195
                                                                                          ? 64'h2D6568636163006C
                                                                                          : auto_in_a_bits_address[11:3] == 9'h194
                                                                                              ? 64'h6576656C2D656863
                                                                                              : auto_in_a_bits_address[11:3] == 9'h193
                                                                                                  ? 64'h61630073656D616E
                                                                                                  : auto_in_a_bits_address[11:3] == 9'h192
                                                                                                      ? 64'h2D67657200736567
                                                                                                      : auto_in_a_bits_address[11:3] == 9'h191
                                                                                                          ? 64'h6E617200656C646E
                                                                                                          : auto_in_a_bits_address[11:3] == 9'h190
                                                                                                              ? 64'h6168700072656C6C
                                                                                                              : auto_in_a_bits_address[11:3] == 9'h18F
                                                                                                                  ? 64'h6F72746E6F632D74
                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h18E
                                                                                                                      ? 64'h7075727265746E69
                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h18D
                                                                                                                          ? 64'h736C6C65632D74
                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h18C
                                                                                                                              ? 64'h7075727265746E69
                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h18B
                                                                                                                                  ? 64'h230074696C70732D
                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h18A
                                                                                                                                      ? 64'h626C740073757461
                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h189
                                                                                                                                          ? 64'h747300736E6F6967
                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h188
                                                                                                                                              ? 64'h6572706D702C7663
                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h187
                                                                                                                                                  ? 64'h7369720079746972
                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h186
                                                                                                                                                      ? 64'h616C756E61726770
                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h185
                                                                                                                                                          ? 64'h6D702C7663736972
                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h184
                                                                                                                                                              ? 64'h6173692C766373
                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h183
                                                                                                                                                                  ? 64'h6972006765720065
                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h182
                                                                                                                                                                      ? 64'h686361632D6C6576
                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h181
                                                                                                                                                                          ? 64'h656C2D7478656E00
                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h180
                                                                                                                                                                              ? 64'h657079742D756D6D
                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h17F
                                                                                                                                                                                  ? 64'h657A69732D626C
                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h17E
                                                                                                                                                                                      ? 64'h742D690073746573
                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h17D
                                                                                                                                                                                          ? 64'h2D626C742D690065
                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h17C
                                                                                                                                                                                              ? 64'h7A69732D65686361
                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h17B
                                                                                                                                                                                                  ? 64'h632D690073746573
                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h17A
                                                                                                                                                                                                      ? 64'h2D65686361632D69
                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h179
                                                                                                                                                                                                          ? 64'h657A69732D6B63
                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h178
                                                                                                                                                                                                              ? 64'h6F6C622D65686361
                                                                                                                                                                                                              : auto_in_a_bits_address[11:3] == 9'h177
                                                                                                                                                                                                                  ? 64'h632D6900746E756F
                                                                                                                                                                                                                  : auto_in_a_bits_address[11:3] == 9'h176
                                                                                                                                                                                                                      ? 64'h632D746E696F706B
                                                                                                                                                                                                                      : auto_in_a_bits_address[11:3] == 9'h175
                                                                                                                                                                                                                          ? 64'h616572622D636578
                                                                                                                                                                                                                          : auto_in_a_bits_address[11:3] == 9'h174 ? 64'h652D657261776472 : auto_in_a_bits_address[11:3] == 9'h173 ? 64'h616800657079745F : auto_in_a_bits_address[11:3] == 9'h172 ? 64'h6563697665640065 : auto_in_a_bits_address[11:3] == 9'h171 ? 64'h7A69732D626C742D : auto_in_a_bits_address[11:3] == 9'h170 ? 64'h6400737465732D62 : auto_in_a_bits_address[11:3] == 9'h16F ? 64'h6C742D6400657A69 : auto_in_a_bits_address[11:3] == 9'h16E ? 64'h732D65686361632D : auto_in_a_bits_address[11:3] == 9'h16D ? 64'h6400737465732D65 : auto_in_a_bits_address[11:3] == 9'h16C ? 64'h686361632D640065 : auto_in_a_bits_address[11:3] == 9'h16B ? 64'h7A69732D6B636F6C : auto_in_a_bits_address[11:3] == 9'h16A ? 64'h622D65686361632D : auto_in_a_bits_address[11:3] == 9'h169 ? 64'h640079636E657571 : auto_in_a_bits_address[11:3] == 9'h168 ? 64'h6572662D6B636F6C : auto_in_a_bits_address[11:3] == 9'h167 ? 64'h630079636E657571 : auto_in_a_bits_address[11:3] == 9'h166 ? 64'h6572662D65736162 : auto_in_a_bits_address[11:3] == 9'h165 ? 64'h656D697400687461 : auto_in_a_bits_address[11:3] == 9'h164 ? 64'h702D74756F647473 : auto_in_a_bits_address[11:3] == 9'h163 ? 64'h306C6169726573 : auto_in_a_bits_address[11:3] == 9'h162 ? 64'h6C65646F6D0065 : auto_in_a_bits_address[11:3] == 9'h161 ? 64'h6C62697461706D6F : auto_in_a_bits_address[11:3] == 9'h160 ? 64'h6300736C6C65632D : auto_in_a_bits_address[11:3] == 9'h15F ? 64'h657A69732300736C : auto_in_a_bits_address[11:3] == 9'h15E ? 64'h6C65632D73736572 : auto_in_a_bits_address[11:3] == 9'h15D ? 64'h6464612309000000 : auto_in_a_bits_address[11:3] == 9'h15C ? 64'h200000002000000 : auto_in_a_bits_address[11:3] == 9'h15B ? 64'h2000000006C6F72 : auto_in_a_bits_address[11:3] == 9'h15A ? 64'h746E6F63A8010000 : auto_in_a_bits_address[11:3] == 9'h159 ? 64'h800000003000000 : _GEN_344;
endmodule

