// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

bind TLXbar TLMonitor_assert TLMonitor_assert (
  .io_in_a_bits_address (auto_in_0_a_bits_address),
  .io_in_a_bits_size    (auto_in_0_a_bits_size),
  .io_in_a_bits_param   (auto_in_0_a_bits_param),
  .io_in_a_bits_mask    (auto_in_0_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_0_a_bits_corrupt),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_d_bits_param   (nodeIn_d_bits_param),
  .io_in_d_bits_corrupt (nodeIn_d_bits_corrupt),
  .io_in_d_bits_denied  (nodeIn_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_0_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_0_a_valid),
  .io_in_a_bits_source  (auto_in_0_a_bits_source),
  .io_in_d_ready        (auto_in_0_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_source  (in_0_d_bits_source),
  .io_in_d_bits_sink    (nodeIn_d_bits_sink)
);
bind TLXbar TLMonitor_1_assert TLMonitor_1_assert (
  .io_in_a_bits_address (auto_in_1_a_bits_address),
  .io_in_a_bits_size    (auto_in_1_a_bits_size),
  .io_in_a_bits_source  (auto_in_1_a_bits_source),
  .io_in_a_bits_param   (auto_in_1_a_bits_param),
  .io_in_a_bits_mask    (auto_in_1_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_1_a_bits_corrupt),
  .io_in_d_bits_opcode  (in_1_d_bits_opcode),
  .io_in_d_bits_source  (in_1_d_bits_source),
  .io_in_d_bits_size    (in_1_d_bits_size),
  .io_in_d_bits_param   (in_1_d_bits_param),
  .io_in_d_bits_corrupt (in_1_d_bits_corrupt),
  .io_in_d_bits_denied  (in_1_d_bits_denied),
  .io_in_b_bits_address (auto_out_1_b_bits_address),
  .io_in_b_bits_param   (auto_out_1_b_bits_param),
  .io_in_c_bits_address (auto_in_1_c_bits_address),
  .io_in_c_bits_source  (auto_in_1_c_bits_source),
  .io_in_c_bits_size    (auto_in_1_c_bits_size),
  .io_in_c_bits_param   (auto_in_1_c_bits_param),
  .io_in_c_bits_corrupt (auto_in_1_c_bits_corrupt),
  .io_in_a_bits_opcode  (auto_in_1_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (in_1_a_ready),
  .io_in_a_valid        (auto_in_1_a_valid),
  .io_in_d_ready        (auto_in_1_d_ready),
  .io_in_d_valid        (in_1_d_valid),
  .io_in_d_bits_sink    (in_1_d_bits_sink),
  .io_in_b_ready        (auto_in_1_b_ready),
  .io_in_b_valid        (auto_out_1_b_valid),
  .io_in_c_bits_opcode  (auto_in_1_c_bits_opcode),
  .io_in_c_ready        (auto_out_1_c_ready),
  .io_in_c_valid        (auto_in_1_c_valid),
  .io_in_e_valid        (auto_in_1_e_valid),
  .io_in_e_bits_sink    (auto_in_1_e_bits_sink)
);
bind TLXbar TLXbar_assert TLXbar_assert (
  .winner__1        (winner__1),
  .prefixOR_1       (prefixOR_1),
  ._out_0_a_valid_T (_out_0_a_valid_T),
  .winner_1_1       (winner_1_1),
  .winner_1_0       (winner_1_0),
  ._out_1_a_valid_T (_out_1_a_valid_T),
  .winner_2_1       (winner_2_1),
  .winner_2_0       (winner_2_0),
  ._in_0_d_valid_T  (_in_0_d_valid_T),
  .winner_3_1       (winner_3_1),
  .winner_3_0       (winner_3_0),
  ._in_1_d_valid_T  (_in_1_d_valid_T),
  .reset            (reset),
  .clock            (clock)
);
bind TLFIFOFixer TLMonitor_2_assert TLMonitor_2_assert (
  .io_in_a_bits_address (auto_in_0_a_bits_address),
  .io_in_a_bits_size    (auto_in_0_a_bits_size),
  .io_in_a_bits_param   (auto_in_0_a_bits_param),
  .io_in_a_bits_mask    (auto_in_0_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_0_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_0_d_bits_opcode),
  .io_in_d_bits_size    (auto_out_0_d_bits_size),
  .io_in_d_bits_param   (auto_out_0_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_0_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_0_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_0_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_0_a_ready),
  .io_in_a_valid        (auto_in_0_a_valid),
  .io_in_a_bits_source  (auto_in_0_a_bits_source),
  .io_in_d_ready        (auto_in_0_d_ready),
  .io_in_d_valid        (auto_out_0_d_valid),
  .io_in_d_bits_source  (auto_out_0_d_bits_source),
  .io_in_d_bits_sink    (auto_out_0_d_bits_sink)
);
bind TLFIFOFixer TLMonitor_3_assert TLMonitor_3_assert (
  .io_in_a_bits_address (auto_in_1_a_bits_address),
  .io_in_a_bits_size    (auto_in_1_a_bits_size),
  .io_in_a_bits_source  (auto_in_1_a_bits_source),
  .io_in_a_bits_param   (auto_in_1_a_bits_param),
  .io_in_a_bits_mask    (auto_in_1_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_1_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_1_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_1_d_bits_source),
  .io_in_d_bits_size    (auto_out_1_d_bits_size),
  .io_in_d_bits_param   (auto_out_1_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_1_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_1_d_bits_denied),
  .io_in_b_bits_address (auto_out_1_b_bits_address),
  .io_in_b_bits_param   (auto_out_1_b_bits_param),
  .io_in_c_bits_address (auto_in_1_c_bits_address),
  .io_in_c_bits_source  (auto_in_1_c_bits_source),
  .io_in_c_bits_size    (auto_in_1_c_bits_size),
  .io_in_c_bits_param   (auto_in_1_c_bits_param),
  .io_in_c_bits_corrupt (auto_in_1_c_bits_corrupt),
  .io_in_a_bits_opcode  (auto_in_1_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_1_a_ready),
  .io_in_a_valid        (auto_in_1_a_valid),
  .io_in_d_ready        (auto_in_1_d_ready),
  .io_in_d_valid        (auto_out_1_d_valid),
  .io_in_d_bits_sink    (auto_out_1_d_bits_sink),
  .io_in_b_ready        (auto_in_1_b_ready),
  .io_in_b_valid        (auto_out_1_b_valid),
  .io_in_c_bits_opcode  (auto_in_1_c_bits_opcode),
  .io_in_c_ready        (auto_out_1_c_ready),
  .io_in_c_valid        (auto_in_1_c_valid),
  .io_in_e_valid        (auto_in_1_e_valid),
  .io_in_e_bits_sink    (auto_in_1_e_bits_sink)
);
bind TLWidthWidget TLMonitor_4_assert TLMonitor_4_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (corrupt_out),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeated_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLWidthWidget_1 TLMonitor_5_assert TLMonitor_5_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_repeated_repeater_io_deq_bits_opcode),
  .io_in_d_bits_size    (_repeated_repeater_io_deq_bits_size),
  .io_in_d_bits_param   (_repeated_repeater_io_deq_bits_param),
  .io_in_d_bits_corrupt (_repeated_repeater_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_repeated_repeater_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_repeated_repeater_io_deq_valid),
  .io_in_d_bits_source  (_repeated_repeater_io_deq_bits_source),
  .io_in_d_bits_sink    (_repeated_repeater_io_deq_bits_sink)
);
bind TLFIFOFixer_1 TLMonitor_6_assert TLMonitor_6_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_out_d_valid)
);
bind TLXbar_2 TLMonitor_7_assert TLMonitor_7_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_source  (nodeIn_d_bits_source),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLXbar_2 TLXbar_2_assert TLXbar_2_assert (
  .winner_1        (winner_1),
  .winner_0        (winner_0),
  ._in_0_d_valid_T (_in_0_d_valid_T),
  .reset           (reset),
  .clock           (clock)
);
bind TLBuffer TLMonitor_8_assert TLMonitor_8_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLAtomicAutomata TLMonitor_9_assert TLMonitor_9_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (nodeIn_d_bits_corrupt),
  .io_in_d_bits_denied  (nodeIn_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLAtomicAutomata TLAtomicAutomata_assert TLAtomicAutomata_assert (
  .winner_1           (winner_1),
  .cam_amo_0          (cam_amo_0),
  ._nodeOut_a_valid_T (_nodeOut_a_valid_T),
  .reset              (reset),
  .clock              (clock)
);
bind TLBuffer_1 TLMonitor_10_assert TLMonitor_10_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLFragmenter TLMonitor_11_assert TLMonitor_11_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLFragmenter TLFragmenter_assert TLFragmenter_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind TLFragmenter_1 TLMonitor_12_assert TLMonitor_12_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLFragmenter_1 TLFragmenter_1_assert TLFragmenter_1_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind PeripheryBus TLMonitor_13_assert TLMonitor_13_assert (
  .io_in_a_bits_source  (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_source),
  .io_in_a_bits_size    (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_size),
  .io_in_a_bits_address (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_address),
  .io_in_a_bits_param   (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_param),
  .io_in_a_bits_mask    (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_mask),
  .io_in_a_bits_corrupt (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN),
  .io_in_d_bits_source  (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_source),
  .io_in_d_bits_size    (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_size),
  .io_in_a_bits_opcode  (_coupler_to_bootaddressreg_auto_fragmenter_out_a_bits_opcode),
  .clock                (_fixedClockNode_auto_out_0_clock),
  .reset                (_fixedClockNode_auto_out_0_reset),
  .io_in_a_ready        (_coupler_to_bootaddressreg_auto_fragmenter_out_d_ready),
  .io_in_a_valid        (_coupler_to_bootaddressreg_auto_fragmenter_out_a_valid),
  .io_in_d_ready        (_coupler_to_bootaddressreg_auto_fragmenter_out_d_ready),
  .io_in_d_valid        (_coupler_to_bootaddressreg_auto_fragmenter_out_a_valid)
);
bind TLBuffer_2 TLMonitor_14_assert TLMonitor_14_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLBuffer_3 TLMonitor_15_assert TLMonitor_15_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLFIFOFixer_2 TLMonitor_16_assert TLMonitor_16_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_out_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLXbar_4 TLMonitor_17_assert TLMonitor_17_assert (
  .io_in_a_bits_address (auto_in_0_a_bits_address),
  .io_in_a_bits_size    (auto_in_0_a_bits_size),
  .io_in_a_bits_source  (auto_in_0_a_bits_source),
  .io_in_a_bits_param   (auto_in_0_a_bits_param),
  .io_in_a_bits_mask    (auto_in_0_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_0_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[5:0]),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_0_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_0_a_valid),
  .io_in_d_ready        (auto_in_0_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLXbar_4 TLMonitor_18_assert TLMonitor_18_assert (
  .io_in_a_bits_address (auto_in_1_a_bits_address),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (in_1_a_ready),
  .io_in_a_valid        (auto_in_1_a_valid),
  .io_in_d_valid        (in_1_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLXbar_4 TLXbar_4_assert TLXbar_4_assert (
  .winner_1         (winner_1),
  .winner_0         (winner_0),
  ._out_0_a_valid_T (_out_0_a_valid_T),
  .reset            (reset),
  .clock            (clock)
);
bind TLXbar_5 TLMonitor_19_assert TLMonitor_19_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_source  (nodeIn_d_bits_source),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_d_bits_param   (nodeIn_d_bits_param),
  .io_in_d_bits_corrupt (nodeIn_d_bits_corrupt),
  .io_in_d_bits_denied  (nodeIn_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (nodeIn_d_bits_sink)
);
bind TLXbar_5 TLXbar_5_assert TLXbar_5_assert (
  .winner_7           (winner_7),
  .winner_6           (winner_6),
  .winner_5           (winner_5),
  .winner_4           (winner_4),
  .winner_3           (winner_3),
  .winner_2           (winner_2),
  .winner_0           (winner_0),
  .winner_1           (winner_1),
  ._in_0_d_valid_T    (_in_0_d_valid_T),
  .auto_out_2_d_valid (auto_out_2_d_valid),
  .auto_out_3_d_valid (auto_out_3_d_valid),
  .auto_out_4_d_valid (auto_out_4_d_valid),
  .auto_out_5_d_valid (auto_out_5_d_valid),
  .auto_out_6_d_valid (auto_out_6_d_valid),
  .auto_out_7_d_valid (auto_out_7_d_valid),
  .reset              (reset),
  .clock              (clock)
);
bind TLBuffer_4 TLMonitor_20_assert TLMonitor_20_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLAtomicAutomata_1 TLMonitor_21_assert TLMonitor_21_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (nodeIn_d_bits_corrupt),
  .io_in_d_bits_denied  (nodeIn_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLAtomicAutomata_1 TLAtomicAutomata_1_assert TLAtomicAutomata_1_assert (
  .winner_1           (winner_1),
  .cam_amo_0          (cam_amo_0),
  ._nodeOut_a_valid_T (_nodeOut_a_valid_T),
  .reset              (reset),
  .clock              (clock)
);
bind TLError TLMonitor_22_assert TLMonitor_22_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (da_bits_opcode),
  .io_in_d_bits_source  (_a_q_io_deq_bits_source),
  .io_in_d_bits_size    (_a_q_io_deq_bits_size),
  .io_in_d_bits_corrupt (da_bits_opcode[0]),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (da_valid)
);
bind TLBuffer_5 TLMonitor_23_assert TLMonitor_23_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLBuffer_6 TLMonitor_24_assert TLMonitor_24_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLFragmenter_2 TLMonitor_25_assert TLMonitor_25_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLFragmenter_2 TLFragmenter_2_assert TLFragmenter_2_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind TLFragmenter_3 TLMonitor_26_assert TLMonitor_26_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLFragmenter_3 TLFragmenter_3_assert TLFragmenter_3_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind TLFragmenter_4 TLMonitor_27_assert TLMonitor_27_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLFragmenter_4 TLFragmenter_4_assert TLFragmenter_4_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind TLFragmenter_5 TLMonitor_28_assert TLMonitor_28_assert (
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLFragmenter_5 TLFragmenter_5_assert TLFragmenter_5_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind TLFragmenter_6 TLMonitor_29_assert TLMonitor_29_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_out_d_valid)
);
bind TLFragmenter_6 TLFragmenter_6_assert TLFragmenter_6_assert (
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .repeater_io_full          (_repeater_io_full),
  .reset                     (reset),
  .clock                     (clock)
);
bind TLFIFOFixer_3 TLMonitor_30_assert TLMonitor_30_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_out_d_valid)
);
bind TLBuffer_8 TLMonitor_31_assert TLMonitor_31_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind TLFIFOFixer_4 TLMonitor_32_assert TLMonitor_32_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_out_d_valid)
);
bind ProbePicker TLMonitor_33_assert TLMonitor_33_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_out_d_valid)
);
bind AXI4UserYanker AXI4UserYanker_assert AXI4UserYanker_assert (
  .auto_out_r_bits_id    (auto_out_r_bits_id),
  .Queue_15_io_deq_valid (_Queue_15_io_deq_valid),
  .Queue_14_io_deq_valid (_Queue_14_io_deq_valid),
  .Queue_13_io_deq_valid (_Queue_13_io_deq_valid),
  .Queue_12_io_deq_valid (_Queue_12_io_deq_valid),
  .Queue_11_io_deq_valid (_Queue_11_io_deq_valid),
  .Queue_10_io_deq_valid (_Queue_10_io_deq_valid),
  .Queue_9_io_deq_valid  (_Queue_9_io_deq_valid),
  .Queue_8_io_deq_valid  (_Queue_8_io_deq_valid),
  .Queue_7_io_deq_valid  (_Queue_7_io_deq_valid),
  .Queue_6_io_deq_valid  (_Queue_6_io_deq_valid),
  .Queue_5_io_deq_valid  (_Queue_5_io_deq_valid),
  .Queue_4_io_deq_valid  (_Queue_4_io_deq_valid),
  .Queue_3_io_deq_valid  (_Queue_3_io_deq_valid),
  .Queue_2_io_deq_valid  (_Queue_2_io_deq_valid),
  .Queue_1_io_deq_valid  (_Queue_1_io_deq_valid),
  .Queue_io_deq_valid    (_Queue_io_deq_valid),
  .auto_out_r_valid      (auto_out_r_valid),
  .auto_out_b_bits_id    (auto_out_b_bits_id),
  .Queue_31_io_deq_valid (_Queue_31_io_deq_valid),
  .Queue_30_io_deq_valid (_Queue_30_io_deq_valid),
  .Queue_29_io_deq_valid (_Queue_29_io_deq_valid),
  .Queue_28_io_deq_valid (_Queue_28_io_deq_valid),
  .Queue_27_io_deq_valid (_Queue_27_io_deq_valid),
  .Queue_26_io_deq_valid (_Queue_26_io_deq_valid),
  .Queue_25_io_deq_valid (_Queue_25_io_deq_valid),
  .Queue_24_io_deq_valid (_Queue_24_io_deq_valid),
  .Queue_23_io_deq_valid (_Queue_23_io_deq_valid),
  .Queue_22_io_deq_valid (_Queue_22_io_deq_valid),
  .Queue_21_io_deq_valid (_Queue_21_io_deq_valid),
  .Queue_20_io_deq_valid (_Queue_20_io_deq_valid),
  .Queue_19_io_deq_valid (_Queue_19_io_deq_valid),
  .Queue_18_io_deq_valid (_Queue_18_io_deq_valid),
  .Queue_17_io_deq_valid (_Queue_17_io_deq_valid),
  .Queue_16_io_deq_valid (_Queue_16_io_deq_valid),
  .auto_out_b_valid      (auto_out_b_valid),
  .reset                 (reset),
  .clock                 (clock)
);
bind TLToAXI4 TLMonitor_34_assert TLMonitor_34_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_source  (nodeIn_d_bits_source),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_d_bits_corrupt (nodeIn_d_bits_corrupt),
  .io_in_d_bits_denied  (nodeIn_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLToAXI4 TLToAXI4_assert TLToAXI4_assert (
  .count_1  (count_1),
  .dec      (dec),
  .inc      (inc),
  .count_2  (count_2),
  .dec_1    (dec_1),
  .inc_1    (inc_1),
  .count_3  (count_3),
  .dec_2    (dec_2),
  .inc_2    (inc_2),
  .count_4  (count_4),
  .dec_3    (dec_3),
  .inc_3    (inc_3),
  .count_5  (count_5),
  .dec_4    (dec_4),
  .inc_4    (inc_4),
  .count_6  (count_6),
  .dec_5    (dec_5),
  .inc_5    (inc_5),
  .count_7  (count_7),
  .dec_6    (dec_6),
  .inc_6    (inc_6),
  .count_8  (count_8),
  .dec_7    (dec_7),
  .inc_7    (inc_7),
  .count_9  (count_9),
  .dec_8    (dec_8),
  .inc_8    (inc_8),
  .count_10 (count_10),
  .dec_9    (dec_9),
  .inc_9    (inc_9),
  .count_11 (count_11),
  .dec_10   (dec_10),
  .inc_10   (inc_10),
  .count_12 (count_12),
  .dec_11   (dec_11),
  .inc_11   (inc_11),
  .count_13 (count_13),
  .dec_12   (dec_12),
  .inc_12   (inc_12),
  .count_14 (count_14),
  .dec_13   (dec_13),
  .inc_13   (inc_13),
  .count_15 (count_15),
  .dec_14   (dec_14),
  .inc_14   (inc_14),
  .count_16 (count_16),
  .dec_15   (dec_15),
  .inc_15   (inc_15),
  .count_17 (count_17),
  .dec_16   (dec_16),
  .inc_16   (inc_16),
  .count_18 (count_18),
  .dec_17   (dec_17),
  .inc_17   (inc_17),
  .count_19 (count_19),
  .dec_18   (dec_18),
  .inc_18   (inc_18),
  .count_20 (count_20),
  .dec_19   (dec_19),
  .inc_19   (inc_19),
  .reset    (reset),
  .clock    (clock)
);
bind InclusiveCacheControl TLMonitor_35_assert TLMonitor_35_assert (
  .io_in_a_bits_source  (auto_ctrl_in_a_bits_source),
  .io_in_a_bits_size    (auto_ctrl_in_a_bits_size),
  .io_in_a_bits_address (auto_ctrl_in_a_bits_address),
  .io_in_a_bits_param   (auto_ctrl_in_a_bits_param),
  .io_in_a_bits_mask    (auto_ctrl_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_ctrl_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN_3),
  .io_in_d_bits_source  (_out_back_q_io_deq_bits_extra_tlrr_extra_source),
  .io_in_d_bits_size    (_out_back_q_io_deq_bits_extra_tlrr_extra_size),
  .io_in_a_bits_opcode  (auto_ctrl_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (in_ready),
  .io_in_a_valid        (auto_ctrl_in_a_valid),
  .io_in_d_ready        (auto_ctrl_in_d_ready),
  .io_in_d_valid        (out_valid)
);
bind InclusiveCache TLMonitor_36_assert TLMonitor_36_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_inclusive_cache_bank_sched_io_in_d_bits_opcode),
  .io_in_d_bits_source  (_inclusive_cache_bank_sched_io_in_d_bits_source),
  .io_in_d_bits_size    (_inclusive_cache_bank_sched_io_in_d_bits_size),
  .io_in_d_bits_param   (_inclusive_cache_bank_sched_io_in_d_bits_param),
  .io_in_d_bits_corrupt (_inclusive_cache_bank_sched_io_in_d_bits_corrupt),
  .io_in_d_bits_denied  (_inclusive_cache_bank_sched_io_in_d_bits_denied),
  .io_in_d_bits_sink    (_inclusive_cache_bank_sched_io_in_d_bits_sink),
  .io_in_b_bits_address (nodeIn_b_bits_address),
  .io_in_b_bits_param   (_inclusive_cache_bank_sched_io_in_b_bits_param),
  .io_in_c_bits_address (auto_in_c_bits_address),
  .io_in_c_bits_source  (auto_in_c_bits_source),
  .io_in_c_bits_size    (auto_in_c_bits_size),
  .io_in_c_bits_param   (auto_in_c_bits_param),
  .io_in_c_bits_corrupt (auto_in_c_bits_corrupt),
  .io_in_e_bits_sink    (auto_in_e_bits_sink),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_inclusive_cache_bank_sched_io_in_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_inclusive_cache_bank_sched_io_in_d_valid),
  .io_in_b_ready        (auto_in_b_ready),
  .io_in_b_valid        (_inclusive_cache_bank_sched_io_in_b_valid),
  .io_in_c_bits_opcode  (auto_in_c_bits_opcode),
  .io_in_c_ready        (_inclusive_cache_bank_sched_io_in_c_ready),
  .io_in_c_valid        (auto_in_c_valid),
  .io_in_e_valid        (auto_in_e_valid)
);
bind SourceB SourceB_assert SourceB_assert (
  .io_req_bits_clients (io_req_bits_clients),
  .io_req_valid        (io_req_valid),
  .reset               (reset),
  .clock               (clock)
);
bind SourceC SourceC_assert SourceC_assert (
  .room               (room),
  .queue_io_count     (_queue_io_count),
  .queue_io_enq_ready (_queue_io_enq_ready),
  .c_valid            (c_valid),
  .reset              (reset),
  .clock              (clock)
);
bind SourceD SourceD_assert SourceD_assert (
  .queue_io_enq_ready       (_queue_io_enq_ready),
  .queue_io_enq_valid_REG_1 (queue_io_enq_valid_REG_1),
  ._io_grant_safe_T_11      (~s3_full),
  .queue_io_deq_valid       (_queue_io_deq_valid),
  .s3_need_r                (s3_need_r),
  .s4_full                  (s4_full),
  .clock                    (clock),
  .s4_latch                 (s4_latch),
  .s3_latch                 (s3_latch),
  .s2_valid_pb              (s2_valid_pb),
  .s2_req_prio_0            (s2_req_prio_0),
  .io_pb_beat_corrupt       (io_pb_beat_corrupt),
  .io_rel_beat_corrupt      (io_rel_beat_corrupt),
  .s3_need_pb               (s3_need_pb),
  .reset                    (reset)
);
bind ListBuffer ListBuffer_assert ListBuffer_assert (
  .valid        (valid),
  .io_pop_bits  (io_pop_bits),
  .io_pop_valid (io_pop_valid),
  .reset        (reset),
  .clock        (clock)
);
bind ListBuffer_1 ListBuffer_1_assert ListBuffer_1_assert (
  .valid        (valid),
  ._GEN         (_GEN_0),
  .io_pop_valid (io_pop_valid),
  .reset        (reset),
  .clock        (clock)
);
bind SinkC SinkC_assert SinkC_assert (
  .c_q_io_deq_valid        (_c_q_io_deq_valid),
  .c_q_io_deq_bits_corrupt (_c_q_io_deq_bits_corrupt),
  .reset                   (reset),
  .clock                   (clock)
);
bind SinkD SinkD_assert SinkD_assert (
  .d_q_io_deq_valid        (_d_q_io_deq_valid),
  .d_q_io_deq_bits_corrupt (_d_q_io_deq_bits_corrupt),
  .d_q_io_deq_bits_denied  (_d_q_io_deq_bits_denied),
  .reset                   (reset),
  .clock                   (clock)
);
bind Directory Directory_assert Directory_assert (
  .wipeDone                 (wipeCount[10]),
  ._q_io_deq_ready_T        (~io_read_valid),
  ._victimLTE_T_7           (_victimLTE_T_7),
  ._victimLTE_T_6           (_victimLTE_T_6),
  ._victimLTE_T_5           (_victimLTE_T_5),
  .victimLFSR_prng_io_out_9 (_victimLFSR_prng_io_out_9),
  ._victimLTE_T_3           (_victimLTE_T_3),
  ._victimLTE_T_2           (|_GEN_3),
  ._victimLTE_T_1           (|_GEN_2),
  .io_read_valid            (io_read_valid),
  .clock                    (clock),
  .reset                    (reset),
  ._view__T_76              (_view__T_76),
  ._view__T_75              (_view__T_75),
  ._view__T_74              (_view__T_74),
  ._view__T_73              (_view__T_73),
  ._view__T_72              (_view__T_72),
  ._view__T_71              (_view__T_71),
  ._GEN                     (~(|_GEN_2))
);
bind ListBuffer_2 ListBuffer_2_assert ListBuffer_2_assert (
  .valid        (valid),
  .io_pop_bits  (io_pop_bits),
  .io_pop_valid (io_pop_valid),
  .reset        (reset),
  .clock        (clock)
);
bind MSHR MSHR_assert MSHR_assert (
  .evict_c                           (evict_c),
  .meta_dirty                        (meta_dirty),
  ._io_status_bits_blockC_output     (~meta_valid),
  ._io_status_bits_nestC_T_3         (~w_grantfirst),
  .w_pprobeacklast                   (w_pprobeacklast),
  .w_rprobeacklast                   (w_rprobeacklast),
  .w_releaseack                      (w_releaseack),
  .meta_valid                        (meta_valid),
  ._io_status_bits_nestC_output      (_io_status_bits_nestC_output),
  ._io_schedule_bits_c_bits_param_T  (_io_schedule_bits_c_bits_param_T),
  .meta_hit                          (meta_hit),
  .meta_state                        (meta_state),
  ._GEN                              (|meta_state),
  .final_meta_writeback_state        (final_meta_writeback_state),
  .after_c                           (after_c),
  .final_meta_writeback_dirty        (final_meta_writeback_dirty),
  .no_wait                           (no_wait),
  .io_schedule_ready                 (io_schedule_ready),
  ._io_schedule_valid_output         (_io_schedule_valid_output),
  .request_valid                     (request_valid),
  .new_meta_hit                      (new_meta_hit),
  .reset                             (reset),
  .clock                             (clock),
  ._final_meta_writeback_state_T_1   (_final_meta_writeback_state_T_1),
  .bad_grant                         (bad_grant),
  ._io_schedule_bits_dir_bits_data_T (~s_release),
  .w_rprobeackfirst                  (w_rprobeackfirst),
  ._io_schedule_bits_dir_valid_T_2   (~s_writeback),
  ._new_meta_T                       (_new_meta_T),
  .io_allocate_valid                 (io_allocate_valid),
  ._GEN_0                            (~new_meta_hit),
  ._GEN_1                            (_GEN_0),
  .new_request_prio_2                (new_request_prio_2)
);
bind InclusiveCacheBankScheduler InclusiveCacheBankScheduler_assert InclusiveCacheBankScheduler_assert (
  .sinkC_io_req_valid  (_sinkC_io_req_valid),
  ._GEN                (_GEN_57),
  .reset               (reset),
  .clock               (clock),
  .request_bits_prio_0 (~_sinkC_io_req_valid)
);
bind TLBuffer_11 TLMonitor_37_assert TLMonitor_37_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink),
  .io_in_b_bits_address (auto_out_b_bits_address),
  .io_in_b_bits_param   (auto_out_b_bits_param),
  .io_in_c_bits_address (auto_in_c_bits_address),
  .io_in_c_bits_source  (auto_in_c_bits_source),
  .io_in_c_bits_size    (auto_in_c_bits_size),
  .io_in_c_bits_param   (auto_in_c_bits_param),
  .io_in_c_bits_corrupt (auto_in_c_bits_corrupt),
  .io_in_e_bits_sink    (auto_in_e_bits_sink),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_b_ready        (auto_in_b_ready),
  .io_in_b_valid        (auto_out_b_valid),
  .io_in_c_bits_opcode  (auto_in_c_bits_opcode),
  .io_in_c_ready        (auto_out_c_ready),
  .io_in_c_valid        (auto_in_c_valid),
  .io_in_e_valid        (auto_in_e_valid)
);
bind TLCacheCork TLMonitor_38_assert TLMonitor_38_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (in_d_bits_opcode),
  .io_in_d_bits_source  (in_d_bits_source),
  .io_in_d_bits_size    (in_d_bits_size),
  .io_in_d_bits_param   (in_d_bits_param),
  .io_in_d_bits_corrupt (in_d_bits_corrupt),
  .io_in_d_bits_denied  (in_d_bits_denied),
  .io_in_c_bits_address (auto_in_c_bits_address),
  .io_in_c_bits_source  (auto_in_c_bits_source),
  .io_in_c_bits_size    (auto_in_c_bits_size),
  .io_in_c_bits_param   (auto_in_c_bits_param),
  .io_in_c_bits_corrupt (auto_in_c_bits_corrupt),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (nodeIn_d_bits_sink),
  .io_in_c_bits_opcode  (auto_in_c_bits_opcode),
  .io_in_c_ready        (nodeIn_c_ready),
  .io_in_c_valid        (auto_in_c_valid),
  .io_in_e_valid        (auto_in_e_valid),
  .io_in_e_bits_sink    (auto_in_e_bits_sink)
);
bind IDPool IDPool_assert IDPool_assert (
  ._GEN          (_GEN),
  .bitmap        (bitmap),
  ._bitmap1_T    (~taken),
  .io_free_valid (io_free_valid),
  .valid         (valid),
  ._valid1_T     (|bitmap),
  .select        (select),
  ._valid1_T_1   (bitmap[0]),
  ._valid1_T_2   (bitmap[1]),
  ._valid1_T_3   (bitmap[2]),
  ._valid1_T_4   (bitmap[3]),
  ._valid1_T_5   (bitmap[4]),
  ._valid1_T_6   (bitmap[5]),
  ._valid1_T_7   (bitmap[6]),
  .reset         (reset),
  .clock         (clock),
  ._GEN_0        (_GEN_0)
);
bind TLCacheCork TLCacheCork_assert TLCacheCork_assert (
  ._nodeIn_c_ready_T  (_nodeIn_c_ready_T),
  ._c_a_valid_T       (&auto_in_c_bits_opcode),
  .auto_in_c_valid    (auto_in_c_valid),
  .winner__1          (winner__1),
  .c_a_valid          (c_a_valid),
  ._nodeOut_a_valid_T (_nodeOut_a_valid_T),
  .winner_1_2         (winner_1_2),
  .auto_out_d_valid   (auto_out_d_valid),
  .winner_1_1         (winner_1_1),
  ._in_d_valid_T      (_in_d_valid_T),
  .q_1_io_deq_valid   (_q_1_io_deq_valid),
  .reset              (reset),
  .clock              (clock)
);
bind BankBinder TLMonitor_39_assert TLMonitor_39_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_out_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_out_d_valid)
);
bind TLXbar_8 TLMonitor_40_assert TLMonitor_40_assert (
  .io_in_a_bits_address (auto_in_0_a_bits_address),
  .io_in_a_bits_size    (auto_in_0_a_bits_size),
  .io_in_a_bits_source  (auto_in_0_a_bits_source),
  .io_in_a_bits_param   (auto_in_0_a_bits_param),
  .io_in_a_bits_mask    (auto_in_0_a_bits_mask),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[3:0]),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .io_in_b_bits_opcode  (auto_out_b_bits_opcode),
  .io_in_b_bits_address (auto_out_b_bits_address),
  .io_in_b_bits_size    (auto_out_b_bits_size),
  .io_in_b_bits_source  (auto_out_b_bits_source[3:0]),
  .io_in_b_bits_param   (auto_out_b_bits_param),
  .io_in_b_bits_mask    (auto_out_b_bits_mask),
  .io_in_b_bits_corrupt (auto_out_b_bits_corrupt),
  .io_in_c_bits_address (auto_in_0_c_bits_address),
  .io_in_c_bits_source  (auto_in_0_c_bits_source),
  .io_in_c_bits_size    (auto_in_0_c_bits_size),
  .io_in_c_bits_param   (auto_in_0_c_bits_param),
  .io_in_a_bits_opcode  (auto_in_0_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_0_a_valid),
  .io_in_d_ready        (auto_in_0_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink),
  .io_in_b_ready        (auto_in_0_b_ready),
  .io_in_b_valid        (nodeIn_b_valid),
  .io_in_c_bits_opcode  (auto_in_0_c_bits_opcode),
  .io_in_c_ready        (auto_out_c_ready),
  .io_in_c_valid        (auto_in_0_c_valid),
  .io_in_e_bits_sink    (auto_in_0_e_bits_sink),
  .io_in_e_ready        (auto_out_e_ready),
  .io_in_e_valid        (auto_in_0_e_valid)
);
bind TLXbar_8 TLMonitor_41_assert TLMonitor_41_assert (
  .io_in_a_bits_address (auto_in_1_a_bits_address),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_size    (auto_out_d_bits_size),
  .io_in_d_bits_param   (auto_out_d_bits_param),
  .io_in_d_bits_corrupt (auto_out_d_bits_corrupt),
  .io_in_d_bits_denied  (auto_out_d_bits_denied),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (in_1_a_ready),
  .io_in_a_valid        (auto_in_1_a_valid),
  .io_in_d_valid        (in_1_d_valid),
  .io_in_d_bits_sink    (auto_out_d_bits_sink)
);
bind TLXbar_8 TLXbar_8_assert TLXbar_8_assert (
  .winner_1         (winner_1),
  .winner_0         (winner_0),
  ._out_0_a_valid_T (_out_0_a_valid_T),
  .reset            (reset),
  .clock            (clock)
);
bind BoomMSHR BoomMSHR_assert BoomMSHR_assert (
  ._io_way_valid_T           (~(|state)),
  .rpq_io_empty              (_rpq_io_empty),
  .rpq_io_enq_ready          (_rpq_io_enq_ready),
  ._state_T_157              (_state_T_157),
  ._state_T_158              (_state_T_158),
  ._state_T_160              (_state_T_160),
  ._state_T_162              (_state_T_162),
  ._state_T_163              (_state_T_163),
  ._state_T_164              (_state_T_164),
  ._state_T_165              (_state_T_165),
  ._state_T_169              (_state_T_169),
  ._state_T_170              (_state_T_170),
  ._state_T_171              (_state_T_171),
  ._state_T_172              (_state_T_172),
  ._state_T_173              (_state_T_173),
  .clock                     (clock),
  .reset                     (reset),
  ._GEN                      (|state),
  ._rpq_io_enq_valid_T       (_rpq_io_enq_valid_T),
  .io_req_old_meta_coh_state (io_req_old_meta_coh_state),
  ._GEN_0                    (_GEN_28),
  ._GEN_1                    (_GEN_18),
  ._GEN_423                  (_GEN_423),
  .grant_had_data            (grant_had_data),
  ._GEN_2                    (_GEN_13),
  .io_req_tag_match          (io_req_tag_match),
  .state_is_hit              (state_is_hit),
  ._io_probe_rdy_T_3         (_io_probe_rdy_T_3),
  .refill_done               (refill_done),
  ._GEN_3026                 (_GEN_3026),
  ._GEN_3                    (_GEN_11),
  ._GEN_4                    (_GEN_12),
  ._GEN_1000                 (_GEN_1000),
  ._GEN_5                    (_GEN_10),
  ._GEN_1398                 (_GEN_1398),
  ._GEN_6                    (_GEN_9),
  ._GEN_7                    (_GEN_8),
  ._GEN_8                    (_GEN_7),
  ._io_probe_rdy_T_8         (_io_probe_rdy_T_8),
  ._io_probe_rdy_T_4         (_io_probe_rdy_T_4),
  ._rpq_io_enq_valid_T_1     (_rpq_io_enq_valid_T_1),
  ._GEN_9                    (_GEN_15),
  ._sec_rdy_T_6              (_sec_rdy_T_6),
  ._sec_rdy_T_5              (_sec_rdy_T_5),
  ._GEN_707                  (_GEN_707),
  .state_is_hit_1            (state_is_hit_1)
);
bind BoomIOMSHR BoomIOMSHR_assert BoomIOMSHR_assert (
  ._io_req_ready_output (_io_req_ready_output),
  .req_uop_mem_cmd      (req_uop_mem_cmd),
  .reset                (reset),
  .clock                (clock)
);
bind BoomMSHRFile BoomMSHRFile_assert BoomMSHRFile_assert (
  .winner__8                    (winner__8),
  .winner__7                    (winner__7),
  .winner__6                    (winner__6),
  .winner__5                    (winner__5),
  .winner__4                    (winner__4),
  .winner__3                    (winner__3),
  .winner__2                    (winner__2),
  .mshrs_0_io_mem_acquire_valid (_mshrs_0_io_mem_acquire_valid),
  .winner__1                    (winner__1),
  ._io_mem_acquire_valid_T      (_io_mem_acquire_valid_T),
  .mshrs_2_io_mem_acquire_valid (_mshrs_2_io_mem_acquire_valid),
  .mshrs_3_io_mem_acquire_valid (_mshrs_3_io_mem_acquire_valid),
  .mshrs_4_io_mem_acquire_valid (_mshrs_4_io_mem_acquire_valid),
  .mshrs_5_io_mem_acquire_valid (_mshrs_5_io_mem_acquire_valid),
  .mshrs_6_io_mem_acquire_valid (_mshrs_6_io_mem_acquire_valid),
  .mshrs_7_io_mem_acquire_valid (_mshrs_7_io_mem_acquire_valid),
  .mmios_0_io_mem_access_valid  (_mmios_0_io_mem_access_valid),
  .winner_1_7                   (winner_1_7),
  .winner_1_6                   (winner_1_6),
  .winner_1_5                   (winner_1_5),
  .winner_1_4                   (winner_1_4),
  .winner_1_3                   (winner_1_3),
  .winner_1_2                   (winner_1_2),
  .mshrs_0_io_mem_finish_valid  (_mshrs_0_io_mem_finish_valid),
  .winner_1_1                   (winner_1_1),
  ._io_mem_finish_valid_T       (_io_mem_finish_valid_T),
  .mshrs_2_io_mem_finish_valid  (_mshrs_2_io_mem_finish_valid),
  .mshrs_3_io_mem_finish_valid  (_mshrs_3_io_mem_finish_valid),
  .mshrs_4_io_mem_finish_valid  (_mshrs_4_io_mem_finish_valid),
  .mshrs_5_io_mem_finish_valid  (_mshrs_5_io_mem_finish_valid),
  .mshrs_6_io_mem_finish_valid  (_mshrs_6_io_mem_finish_valid),
  .mshrs_7_io_mem_finish_valid  (_mshrs_7_io_mem_finish_valid),
  .reset                        (reset),
  .clock                        (clock)
);
bind BoomNonBlockingDCache BoomNonBlockingDCache_assert BoomNonBlockingDCache_assert (
  ._wb_fire_T                  (_wb_fire_T),
  ._wb_fire_T_1                (_wb_fire_T_1),
  .io_lsu_s1_kill_0            (io_lsu_s1_kill_0),
  .io_lsu_req_bits_0_valid     (io_lsu_req_bits_0_valid),
  .clock                       (clock),
  ._s1_valid_T_19              (_s1_valid_T_19),
  .io_lsu_s1_kill_1            (io_lsu_s1_kill_1),
  .io_lsu_req_bits_1_valid     (io_lsu_req_bits_1_valid),
  ._s2_sc_T_2                  (~(|s2_type)),
  ._mshrs_io_req_0_valid_T     (~s2_hit_0),
  ._s2_hit_T_15                (_s2_hit_T_15),
  .reset                       (reset),
  .s2_valid_0                  (s2_valid_0),
  .s2_sc_fail                  (s2_sc_fail),
  .s2_sc                       (s2_sc),
  .s2_req_0_addr               (s2_req_0_addr),
  .s2_send_resp_0              (s2_send_resp_0),
  .s2_send_nack_0              (s2_send_nack_0),
  .s2_send_resp_1              (s2_send_resp_1),
  .s2_send_nack_1              (s2_send_nack_1),
  ._mshrs_io_req_0_valid_T_74  (_mshrs_io_req_0_valid_T_74),
  ._mshrs_io_req_1_valid_T_74  (_mshrs_io_req_1_valid_T_74),
  .winner_1                    (winner_1),
  .wb_io_release_valid         (_wb_io_release_valid),
  ._nodeOut_c_valid_T          (_nodeOut_c_valid_T),
  ._io_lsu_nack_0_valid_output (_io_lsu_nack_0_valid_output),
  .s2_type                     (s2_type),
  ._io_lsu_nack_1_valid_output (_io_lsu_nack_1_valid_output),
  ._s2_nack_victim_T_2         (_s2_nack_victim_T_2),
  ._s3_valid_T_25              (~s2_sc_fail),
  .s2_nack_1                   (s2_nack_1),
  ._mshrs_io_req_1_valid_T_50  (_mshrs_io_req_1_valid_T_50),
  ._mshrs_io_req_1_valid_T_51  (_mshrs_io_req_1_valid_T_51),
  ._mshrs_io_req_1_valid_T_53  (_mshrs_io_req_1_valid_T_53),
  ._mshrs_io_req_1_valid_T_55  (_mshrs_io_req_1_valid_T_55),
  ._mshrs_io_req_1_valid_T_56  (_mshrs_io_req_1_valid_T_56),
  ._mshrs_io_req_1_valid_T_57  (_mshrs_io_req_1_valid_T_57),
  ._mshrs_io_req_1_valid_T_58  (_mshrs_io_req_1_valid_T_58),
  ._mshrs_io_req_1_valid_T_62  (_mshrs_io_req_1_valid_T_62),
  ._mshrs_io_req_1_valid_T_63  (_mshrs_io_req_1_valid_T_63),
  ._mshrs_io_req_1_valid_T_64  (_mshrs_io_req_1_valid_T_64),
  ._mshrs_io_req_1_valid_T_65  (_mshrs_io_req_1_valid_T_65),
  ._mshrs_io_req_1_valid_T_66  (_mshrs_io_req_1_valid_T_66)
);
bind ICache ICache_assert ICache_assert (
  .s1_valid     (s1_valid),
  .s1_tag_hit_7 (s1_tag_hit_7),
  .s1_tag_hit_6 (s1_tag_hit_6),
  .s1_tag_hit_5 (s1_tag_hit_5),
  .s1_tag_hit_4 (s1_tag_hit_4),
  .s1_tag_hit_3 (s1_tag_hit_3),
  .s1_tag_hit_2 (s1_tag_hit_2),
  .s1_tag_hit_1 (s1_tag_hit_1),
  .s1_tag_hit_0 (s1_tag_hit_0),
  .reset        (reset),
  .clock        (clock)
);
bind BranchPredictor BranchPredictor_assert BranchPredictor_assert (
  .io_update_bits_br_mask       (io_update_bits_br_mask),
  .io_update_bits_cfi_idx_bits  (io_update_bits_cfi_idx_bits),
  .io_update_valid              (io_update_valid),
  .io_update_bits_cfi_is_br     (io_update_bits_cfi_is_br),
  .io_update_bits_cfi_idx_valid (io_update_bits_cfi_idx_valid),
  .reset                        (reset),
  .clock                        (clock)
);
bind TLB TLB_assert TLB_assert (
  .vpn                 (io_req_bits_vaddr[38:12]),
  .io_sfence_bits_addr (io_sfence_bits_addr),
  .io_sfence_bits_rs1  (io_sfence_bits_rs1),
  .io_sfence_valid     (io_sfence_valid),
  .reset               (reset),
  .clock               (clock)
);
bind BoomFrontend BoomFrontend_assert BoomFrontend_assert (
  .f3_bpd_resp_io_deq_bits_pc         (_f3_bpd_resp_io_deq_bits_pc),
  .f3_io_deq_bits_pc                  (_f3_io_deq_bits_pc),
  ._f4_btb_corrections_io_enq_valid_T (_f4_btb_corrections_io_enq_valid_T),
  ._GEN                               (~reset),
  .clock                              (clock)
);
bind MemAddrCalcUnit MemAddrCalcUnit_assert MemAddrCalcUnit_assert (
  .io_req_bits_rs2_data        (io_req_bits_rs2_data),
  .io_req_valid                (io_req_valid),
  .io_req_bits_uop_ctrl_is_std (io_req_bits_uop_ctrl_is_std),
  .io_req_bits_uop_fp_val      (io_req_bits_uop_fp_val),
  .io_req_bits_uop_uopc        (io_req_bits_uop_uopc),
  .ma_ld                       (ma_ld),
  .ma_st                       (ma_st),
  .reset                       (reset),
  .clock                       (clock)
);
bind IntToFPUnit IntToFPUnit_assert IntToFPUnit_assert (
  .io_req_valid                 (io_req_valid),
  .fp_decoder_io_sigs_fromint   (_fp_decoder_io_sigs_fromint),
  .io_req_bits_rs1_data         (io_req_bits_rs1_data),
  .fp_decoder_io_sigs_typeTagIn (_fp_decoder_io_sigs_typeTagIn),
  .reset                        (reset),
  .clock                        (clock)
);
bind ALUExeUnit_2 ALUExeUnit_2_assert ALUExeUnit_2_assert (
  .queue_io_enq_ready (_queue_io_enq_ready),
  .reset              (reset),
  .clock              (clock)
);
bind ALUUnit_1 ALUUnit_1_assert ALUUnit_1_assert (
  .pc_sel       (pc_sel),
  .brinfo_valid (brinfo_valid),
  .reset        (reset),
  .clock        (clock)
);
bind ALUUnit_2 ALUUnit_2_assert ALUUnit_2_assert (
  .pc_sel       (pc_sel),
  .brinfo_valid (brinfo_valid),
  .reset        (reset),
  .clock        (clock)
);
bind ALUExeUnit_4 ALUExeUnit_4_assert ALUExeUnit_4_assert (
  .PipelinedMulUnit_io_resp_valid (_PipelinedMulUnit_io_resp_valid),
  .ALUUnit_io_resp_valid          (_ALUUnit_io_resp_valid),
  .reset                          (reset),
  .clock                          (clock)
);
bind ALUExeUnit_5 ALUExeUnit_5_assert ALUExeUnit_5_assert (
  .DivUnit_io_resp_valid (_DivUnit_io_resp_valid),
  .ALUUnit_io_resp_valid (_ALUUnit_io_resp_valid),
  .reset                 (reset),
  .clock                 (clock)
);
bind FDivSqrtUnit FDivSqrtUnit_assert FDivSqrtUnit_assert (
  .r_buffer_val        (r_buffer_val),
  .io_req_valid        (io_req_valid),
  .r_divsqrt_val       (r_divsqrt_val),
  .r_out_val           (r_out_val),
  ._GEN                (_GEN),
  .reset               (reset),
  .clock               (clock),
  ._may_fire_input_T_2 (~r_divsqrt_val)
);
bind FPUExeUnit FPUExeUnit_assert FPUExeUnit_assert (
  .queue_io_enq_ready       (_queue_io_enq_ready),
  ._fp_sdq_io_enq_valid_T_5 (_fp_sdq_io_enq_valid_T_5),
  .fp_sdq_io_enq_ready      (_fp_sdq_io_enq_ready),
  .reset                    (reset),
  .clock                    (clock)
);
bind IssueSlot IssueSlot_assert IssueSlot_assert (
  .io_clear        (io_clear),
  .io_kill         (io_kill),
  .state           (state),
  .io_in_uop_valid (io_in_uop_valid),
  .reset           (reset),
  .clock           (clock)
);
bind IssueUnitCollapsing IssueUnitCollapsing_assert IssueUnitCollapsing_assert (
  .issue_slots_31_grant (issue_slots_31_grant),
  .issue_slots_30_grant (issue_slots_30_grant),
  .issue_slots_29_grant (issue_slots_29_grant),
  .issue_slots_28_grant (issue_slots_28_grant),
  .issue_slots_27_grant (issue_slots_27_grant),
  .issue_slots_26_grant (issue_slots_26_grant),
  .issue_slots_25_grant (issue_slots_25_grant),
  .issue_slots_24_grant (issue_slots_24_grant),
  .issue_slots_23_grant (issue_slots_23_grant),
  .issue_slots_22_grant (issue_slots_22_grant),
  .issue_slots_21_grant (issue_slots_21_grant),
  .issue_slots_20_grant (issue_slots_20_grant),
  .issue_slots_19_grant (issue_slots_19_grant),
  .issue_slots_18_grant (issue_slots_18_grant),
  .issue_slots_17_grant (issue_slots_17_grant),
  .issue_slots_16_grant (issue_slots_16_grant),
  .issue_slots_15_grant (issue_slots_15_grant),
  .issue_slots_14_grant (issue_slots_14_grant),
  .issue_slots_13_grant (issue_slots_13_grant),
  .issue_slots_12_grant (issue_slots_12_grant),
  .issue_slots_11_grant (issue_slots_11_grant),
  .issue_slots_10_grant (issue_slots_10_grant),
  .issue_slots_9_grant  (issue_slots_9_grant),
  .issue_slots_8_grant  (issue_slots_8_grant),
  .issue_slots_7_grant  (issue_slots_7_grant),
  .issue_slots_6_grant  (issue_slots_6_grant),
  .issue_slots_5_grant  (issue_slots_5_grant),
  .issue_slots_4_grant  (issue_slots_4_grant),
  .issue_slots_3_grant  (issue_slots_3_grant),
  .issue_slots_2_grant  (issue_slots_2_grant),
  .issue_slots_1_grant  (issue_slots_1_grant),
  .issue_slots_0_grant  (issue_slots_0_grant),
  .reset                (reset),
  .clock                (clock)
);
bind RegisterFileSynthesizable RegisterFileSynthesizable_assert RegisterFileSynthesizable_assert (
  .io_write_ports_0_bits_addr (io_write_ports_0_bits_addr),
  .io_write_ports_1_bits_addr (io_write_ports_1_bits_addr),
  .io_write_ports_1_valid     (io_write_ports_1_valid),
  .io_write_ports_0_valid     (io_write_ports_0_valid),
  .io_write_ports_2_bits_addr (io_write_ports_2_bits_addr),
  .io_write_ports_2_valid     (io_write_ports_2_valid),
  .io_write_ports_3_bits_addr (io_write_ports_3_bits_addr),
  .io_write_ports_3_valid     (io_write_ports_3_valid),
  .reset                      (reset),
  .clock                      (clock)
);
bind FpPipeline FpPipeline_assert FpPipeline_assert (
  .ll_wbarb_io_in_0_ready                    (_ll_wbarb_io_in_0_ready),
  .io_from_int_bits_uop_dst_rtype            (io_from_int_bits_uop_dst_rtype),
  ._fregfile_io_write_ports_2_valid_T        (_fregfile_io_write_ports_2_valid_T),
  ._io_wakeups_2_valid_T                     (_io_wakeups_2_valid_T),
  ._fregfile_io_write_ports_3_valid_T        (_fregfile_io_write_ports_3_valid_T),
  ._io_wakeups_3_valid_T                     (_io_wakeups_3_valid_T),
  .fpu_exe_unit_io_fresp_valid               (_fpu_exe_unit_io_fresp_valid),
  .fpu_exe_unit_io_fresp_bits_uop_uses_ldq   (_fpu_exe_unit_io_fresp_bits_uop_uses_ldq),
  .fpu_exe_unit_io_fresp_bits_uop_uses_stq   (_fpu_exe_unit_io_fresp_bits_uop_uses_stq),
  .fpu_exe_unit_io_fresp_bits_uop_is_amo     (_fpu_exe_unit_io_fresp_bits_uop_is_amo),
  .fpu_exe_unit_1_io_fresp_valid             (_fpu_exe_unit_1_io_fresp_valid),
  .fpu_exe_unit_1_io_fresp_bits_uop_uses_ldq (_fpu_exe_unit_1_io_fresp_bits_uop_uses_ldq),
  .fpu_exe_unit_1_io_fresp_bits_uop_uses_stq (_fpu_exe_unit_1_io_fresp_bits_uop_uses_stq),
  .fpu_exe_unit_1_io_fresp_bits_uop_is_amo   (_fpu_exe_unit_1_io_fresp_bits_uop_is_amo),
  .reset                                     (reset),
  .clock                                     (clock),
  .io_from_int_valid                         (io_from_int_valid)
);
bind RenameMapTable RenameMapTable_assert RenameMapTable_assert (
  .io_rollback           (io_rollback),
  .io_remap_reqs_0_pdst  (io_remap_reqs_0_pdst),
  .map_table_31          (map_table_31),
  .map_table_30          (map_table_30),
  .map_table_29          (map_table_29),
  .map_table_28          (map_table_28),
  .map_table_27          (map_table_27),
  .map_table_26          (map_table_26),
  .map_table_25          (map_table_25),
  .map_table_24          (map_table_24),
  .map_table_23          (map_table_23),
  .map_table_22          (map_table_22),
  .map_table_21          (map_table_21),
  .map_table_20          (map_table_20),
  .map_table_19          (map_table_19),
  .map_table_18          (map_table_18),
  .map_table_17          (map_table_17),
  .map_table_16          (map_table_16),
  .map_table_15          (map_table_15),
  .map_table_14          (map_table_14),
  .map_table_13          (map_table_13),
  .map_table_12          (map_table_12),
  .map_table_11          (map_table_11),
  .map_table_10          (map_table_10),
  .map_table_9           (map_table_9),
  .map_table_8           (map_table_8),
  .map_table_7           (map_table_7),
  .map_table_6           (map_table_6),
  .map_table_5           (map_table_5),
  .map_table_4           (map_table_4),
  .map_table_3           (map_table_3),
  .map_table_2           (map_table_2),
  .map_table_1           (map_table_1),
  .map_table_0           (map_table_0),
  .io_remap_reqs_0_valid (io_remap_reqs_0_valid),
  .io_remap_reqs_1_pdst  (io_remap_reqs_1_pdst),
  .io_remap_reqs_1_valid (io_remap_reqs_1_valid),
  .io_remap_reqs_2_pdst  (io_remap_reqs_2_pdst),
  .io_remap_reqs_2_valid (io_remap_reqs_2_valid),
  .io_remap_reqs_3_pdst  (io_remap_reqs_3_pdst),
  .io_remap_reqs_3_valid (io_remap_reqs_3_valid),
  .reset                 (reset),
  .clock                 (clock)
);
bind RenameFreeList RenameFreeList_assert RenameFreeList_assert (
  .dealloc_mask            (dealloc_mask),
  .free_list               (free_list),
  .allocs_3                (allocs_3),
  .r_valid_3               (r_valid_3),
  .allocs_2                (allocs_2),
  .r_valid_2               (r_valid_2),
  .allocs_1                (allocs_1),
  .r_valid_1               (r_valid_1),
  .allocs_0                (allocs_0),
  .r_valid                 (r_valid),
  .io_debug_pipeline_empty (io_debug_pipeline_empty),
  .reset                   (reset),
  .clock                   (clock)
);
bind RenameStage RenameStage_assert RenameStage_assert (
  .freelist_io_alloc_pregs_3_bits      (_freelist_io_alloc_pregs_3_bits),
  .ren2_alloc_reqs_3                   (ren2_alloc_reqs_3),
  .freelist_io_alloc_pregs_2_bits      (_freelist_io_alloc_pregs_2_bits),
  .ren2_alloc_reqs_2                   (ren2_alloc_reqs_2),
  .freelist_io_alloc_pregs_1_bits      (_freelist_io_alloc_pregs_1_bits),
  .ren2_alloc_reqs_1                   (ren2_alloc_reqs_1),
  .freelist_io_alloc_pregs_0_bits      (_freelist_io_alloc_pregs_0_bits),
  .ren2_alloc_reqs_0                   (ren2_alloc_reqs_0),
  .io_wakeups_9_valid                  (io_wakeups_9_valid),
  .io_wakeups_9_bits_uop_dst_rtype     (io_wakeups_9_bits_uop_dst_rtype),
  .io_wakeups_8_valid                  (io_wakeups_8_valid),
  .io_wakeups_8_bits_uop_dst_rtype     (io_wakeups_8_bits_uop_dst_rtype),
  .io_wakeups_7_valid                  (io_wakeups_7_valid),
  .io_wakeups_7_bits_uop_dst_rtype     (io_wakeups_7_bits_uop_dst_rtype),
  .io_wakeups_6_valid                  (io_wakeups_6_valid),
  .io_wakeups_6_bits_uop_dst_rtype     (io_wakeups_6_bits_uop_dst_rtype),
  .io_wakeups_5_valid                  (io_wakeups_5_valid),
  .io_wakeups_5_bits_uop_dst_rtype     (io_wakeups_5_bits_uop_dst_rtype),
  .io_wakeups_4_valid                  (io_wakeups_4_valid),
  .io_wakeups_4_bits_uop_dst_rtype     (io_wakeups_4_bits_uop_dst_rtype),
  .io_wakeups_3_valid                  (io_wakeups_3_valid),
  .io_wakeups_3_bits_uop_dst_rtype     (io_wakeups_3_bits_uop_dst_rtype),
  .io_wakeups_2_valid                  (io_wakeups_2_valid),
  .io_wakeups_2_bits_uop_dst_rtype     (io_wakeups_2_bits_uop_dst_rtype),
  .io_wakeups_1_valid                  (io_wakeups_1_valid),
  .io_wakeups_1_bits_uop_dst_rtype     (io_wakeups_1_bits_uop_dst_rtype),
  .io_wakeups_0_valid                  (io_wakeups_0_valid),
  .io_wakeups_0_bits_uop_dst_rtype     (io_wakeups_0_bits_uop_dst_rtype),
  .r_valid                             (r_valid),
  .busytable_io_busy_resps_0_prs1_busy (_busytable_io_busy_resps_0_prs1_busy),
  .r_uop_lrs1                          (r_uop_lrs1),
  .busytable_io_busy_resps_0_prs2_busy (_busytable_io_busy_resps_0_prs2_busy),
  .r_uop_lrs2                          (r_uop_lrs2),
  .r_valid_1                           (r_valid_1),
  .busytable_io_busy_resps_1_prs1_busy (_busytable_io_busy_resps_1_prs1_busy),
  .r_uop_1_lrs1                        (r_uop_1_lrs1),
  .busytable_io_busy_resps_1_prs2_busy (_busytable_io_busy_resps_1_prs2_busy),
  .r_uop_1_lrs2                        (r_uop_1_lrs2),
  .r_valid_2                           (r_valid_2),
  .busytable_io_busy_resps_2_prs1_busy (_busytable_io_busy_resps_2_prs1_busy),
  .r_uop_2_lrs1                        (r_uop_2_lrs1),
  .busytable_io_busy_resps_2_prs2_busy (_busytable_io_busy_resps_2_prs2_busy),
  .r_uop_2_lrs2                        (r_uop_2_lrs2),
  .r_valid_3                           (r_valid_3),
  .busytable_io_busy_resps_3_prs1_busy (_busytable_io_busy_resps_3_prs1_busy),
  .r_uop_3_lrs1                        (r_uop_3_lrs1),
  .busytable_io_busy_resps_3_prs2_busy (_busytable_io_busy_resps_3_prs2_busy),
  .r_uop_3_lrs2                        (r_uop_3_lrs2),
  .reset                               (reset),
  .clock                               (clock)
);
bind RenameMapTable_1 RenameMapTable_1_assert RenameMapTable_1_assert (
  .io_rollback           (io_rollback),
  .io_remap_reqs_0_pdst  (io_remap_reqs_0_pdst),
  .map_table_31          (map_table_31),
  .map_table_30          (map_table_30),
  .map_table_29          (map_table_29),
  .map_table_28          (map_table_28),
  .map_table_27          (map_table_27),
  .map_table_26          (map_table_26),
  .map_table_25          (map_table_25),
  .map_table_24          (map_table_24),
  .map_table_23          (map_table_23),
  .map_table_22          (map_table_22),
  .map_table_21          (map_table_21),
  .map_table_20          (map_table_20),
  .map_table_19          (map_table_19),
  .map_table_18          (map_table_18),
  .map_table_17          (map_table_17),
  .map_table_16          (map_table_16),
  .map_table_15          (map_table_15),
  .map_table_14          (map_table_14),
  .map_table_13          (map_table_13),
  .map_table_12          (map_table_12),
  .map_table_11          (map_table_11),
  .map_table_10          (map_table_10),
  .map_table_9           (map_table_9),
  .map_table_8           (map_table_8),
  .map_table_7           (map_table_7),
  .map_table_6           (map_table_6),
  .map_table_5           (map_table_5),
  .map_table_4           (map_table_4),
  .map_table_3           (map_table_3),
  .map_table_2           (map_table_2),
  .map_table_1           (map_table_1),
  .map_table_0           (map_table_0),
  .io_remap_reqs_0_valid (io_remap_reqs_0_valid),
  .io_remap_reqs_1_pdst  (io_remap_reqs_1_pdst),
  .io_remap_reqs_1_valid (io_remap_reqs_1_valid),
  .io_remap_reqs_2_pdst  (io_remap_reqs_2_pdst),
  .io_remap_reqs_2_valid (io_remap_reqs_2_valid),
  .io_remap_reqs_3_pdst  (io_remap_reqs_3_pdst),
  .io_remap_reqs_3_valid (io_remap_reqs_3_valid),
  .reset                 (reset),
  .clock                 (clock)
);
bind RenameFreeList_1 RenameFreeList_1_assert RenameFreeList_1_assert (
  .dealloc_mask            (dealloc_mask),
  .free_list               (free_list),
  .allocs_3                (allocs_3),
  .r_valid_3               (r_valid_3),
  .allocs_2                (allocs_2),
  .r_valid_2               (r_valid_2),
  .allocs_1                (allocs_1),
  .r_valid_1               (r_valid_1),
  .allocs_0                (allocs_0),
  .r_valid                 (r_valid),
  .io_debug_pipeline_empty (io_debug_pipeline_empty),
  .reset                   (reset),
  .clock                   (clock)
);
bind RenameStage_1 RenameStage_1_assert RenameStage_1_assert (
  .freelist_io_alloc_pregs_3_bits  (_freelist_io_alloc_pregs_3_bits),
  .ren2_alloc_reqs_3               (ren2_alloc_reqs_3),
  .freelist_io_alloc_pregs_2_bits  (_freelist_io_alloc_pregs_2_bits),
  .ren2_alloc_reqs_2               (ren2_alloc_reqs_2),
  .freelist_io_alloc_pregs_1_bits  (_freelist_io_alloc_pregs_1_bits),
  .ren2_alloc_reqs_1               (ren2_alloc_reqs_1),
  .freelist_io_alloc_pregs_0_bits  (_freelist_io_alloc_pregs_0_bits),
  .ren2_alloc_reqs_0               (ren2_alloc_reqs_0),
  .io_wakeups_3_valid              (io_wakeups_3_valid),
  .io_wakeups_3_bits_uop_dst_rtype (io_wakeups_3_bits_uop_dst_rtype),
  .io_wakeups_2_valid              (io_wakeups_2_valid),
  .io_wakeups_2_bits_uop_dst_rtype (io_wakeups_2_bits_uop_dst_rtype),
  .io_wakeups_1_valid              (io_wakeups_1_valid),
  .io_wakeups_1_bits_uop_dst_rtype (io_wakeups_1_bits_uop_dst_rtype),
  .io_wakeups_0_valid              (io_wakeups_0_valid),
  .io_wakeups_0_bits_uop_dst_rtype (io_wakeups_0_bits_uop_dst_rtype),
  .reset                           (reset),
  .clock                           (clock)
);
bind IssueSlot_32 IssueSlot_32_assert IssueSlot_32_assert (
  .io_clear                  (io_clear),
  .io_kill                   (io_kill),
  .state                     (state),
  .next_uop_prs1             (next_uop_prs1),
  .next_uop_prs2             (next_uop_prs2),
  .io_spec_ld_wakeup_0_valid (io_spec_ld_wakeup_0_valid),
  .io_spec_ld_wakeup_0_bits  (io_spec_ld_wakeup_0_bits),
  .io_spec_ld_wakeup_1_valid (io_spec_ld_wakeup_1_valid),
  .io_spec_ld_wakeup_1_bits  (io_spec_ld_wakeup_1_bits),
  .next_p1_poisoned          (next_p1_poisoned),
  .next_p2_poisoned          (next_p2_poisoned),
  .io_in_uop_valid           (io_in_uop_valid),
  .reset                     (reset),
  .clock                     (clock),
  ._GEN                      (_GEN_7),
  ._GEN_0                    (_GEN_8),
  ._GEN_140                  (_GEN_140),
  ._GEN_142                  (_GEN_142),
  ._GEN_1                    (_GEN_11),
  ._GEN_2                    (_GEN_12)
);
bind IssueUnitCollapsing_1 IssueUnitCollapsing_1_assert IssueUnitCollapsing_1_assert (
  .issue_slots_23_grant (issue_slots_23_grant),
  .issue_slots_22_grant (issue_slots_22_grant),
  .issue_slots_21_grant (issue_slots_21_grant),
  .issue_slots_20_grant (issue_slots_20_grant),
  .issue_slots_19_grant (issue_slots_19_grant),
  .issue_slots_18_grant (issue_slots_18_grant),
  .issue_slots_17_grant (issue_slots_17_grant),
  .issue_slots_16_grant (issue_slots_16_grant),
  .issue_slots_15_grant (issue_slots_15_grant),
  .issue_slots_14_grant (issue_slots_14_grant),
  .issue_slots_13_grant (issue_slots_13_grant),
  .issue_slots_12_grant (issue_slots_12_grant),
  .issue_slots_11_grant (issue_slots_11_grant),
  .issue_slots_10_grant (issue_slots_10_grant),
  .issue_slots_9_grant  (issue_slots_9_grant),
  .issue_slots_8_grant  (issue_slots_8_grant),
  .issue_slots_7_grant  (issue_slots_7_grant),
  .issue_slots_6_grant  (issue_slots_6_grant),
  .issue_slots_5_grant  (issue_slots_5_grant),
  .issue_slots_4_grant  (issue_slots_4_grant),
  .issue_slots_3_grant  (issue_slots_3_grant),
  .issue_slots_2_grant  (issue_slots_2_grant),
  .issue_slots_1_grant  (issue_slots_1_grant),
  .issue_slots_0_grant  (issue_slots_0_grant),
  .reset                (reset),
  .clock                (clock)
);
bind IssueUnitCollapsing_2 IssueUnitCollapsing_2_assert IssueUnitCollapsing_2_assert (
  .issue_slots_39_grant (issue_slots_39_grant),
  .issue_slots_38_grant (issue_slots_38_grant),
  .issue_slots_37_grant (issue_slots_37_grant),
  .issue_slots_36_grant (issue_slots_36_grant),
  .issue_slots_35_grant (issue_slots_35_grant),
  .issue_slots_34_grant (issue_slots_34_grant),
  .issue_slots_33_grant (issue_slots_33_grant),
  .issue_slots_32_grant (issue_slots_32_grant),
  .issue_slots_31_grant (issue_slots_31_grant),
  .issue_slots_30_grant (issue_slots_30_grant),
  .issue_slots_29_grant (issue_slots_29_grant),
  .issue_slots_28_grant (issue_slots_28_grant),
  .issue_slots_27_grant (issue_slots_27_grant),
  .issue_slots_26_grant (issue_slots_26_grant),
  .issue_slots_25_grant (issue_slots_25_grant),
  .issue_slots_24_grant (issue_slots_24_grant),
  .issue_slots_23_grant (issue_slots_23_grant),
  .issue_slots_22_grant (issue_slots_22_grant),
  .issue_slots_21_grant (issue_slots_21_grant),
  .issue_slots_20_grant (issue_slots_20_grant),
  .issue_slots_19_grant (issue_slots_19_grant),
  .issue_slots_18_grant (issue_slots_18_grant),
  .issue_slots_17_grant (issue_slots_17_grant),
  .issue_slots_16_grant (issue_slots_16_grant),
  .issue_slots_15_grant (issue_slots_15_grant),
  .issue_slots_14_grant (issue_slots_14_grant),
  .issue_slots_13_grant (issue_slots_13_grant),
  .issue_slots_12_grant (issue_slots_12_grant),
  .issue_slots_11_grant (issue_slots_11_grant),
  .issue_slots_10_grant (issue_slots_10_grant),
  .issue_slots_9_grant  (issue_slots_9_grant),
  .issue_slots_8_grant  (issue_slots_8_grant),
  .issue_slots_7_grant  (issue_slots_7_grant),
  .issue_slots_6_grant  (issue_slots_6_grant),
  .issue_slots_5_grant  (issue_slots_5_grant),
  .issue_slots_4_grant  (issue_slots_4_grant),
  .issue_slots_3_grant  (issue_slots_3_grant),
  .issue_slots_2_grant  (issue_slots_2_grant),
  .issue_slots_1_grant  (issue_slots_1_grant),
  .issue_slots_0_grant  (issue_slots_0_grant),
  .reset                (reset),
  .clock                (clock)
);
bind RegisterFileSynthesizable_1 RegisterFileSynthesizable_1_assert RegisterFileSynthesizable_1_assert (
  .io_write_ports_0_bits_addr (io_write_ports_0_bits_addr),
  .io_write_ports_1_bits_addr (io_write_ports_1_bits_addr),
  .io_write_ports_1_valid     (io_write_ports_1_valid),
  .io_write_ports_0_valid     (io_write_ports_0_valid),
  .io_write_ports_2_bits_addr (io_write_ports_2_bits_addr),
  .io_write_ports_2_valid     (io_write_ports_2_valid),
  .io_write_ports_3_bits_addr (io_write_ports_3_bits_addr),
  .io_write_ports_3_valid     (io_write_ports_3_valid),
  .io_write_ports_4_bits_addr (io_write_ports_4_bits_addr),
  .io_write_ports_4_valid     (io_write_ports_4_valid),
  .io_write_ports_5_bits_addr (io_write_ports_5_bits_addr),
  .io_write_ports_5_valid     (io_write_ports_5_valid),
  .reset                      (reset),
  .clock                      (clock)
);
bind Rob Rob_assert Rob_assert (
  .rob_tail                          (rob_tail),
  .rob_val__31                       (rob_val__31),
  .rob_val__30                       (rob_val__30),
  .rob_val__29                       (rob_val__29),
  .rob_val__28                       (rob_val__28),
  .rob_val__27                       (rob_val__27),
  .rob_val__26                       (rob_val__26),
  .rob_val__25                       (rob_val__25),
  .rob_val__24                       (rob_val__24),
  .rob_val__23                       (rob_val__23),
  .rob_val__22                       (rob_val__22),
  .rob_val__21                       (rob_val__21),
  .rob_val__20                       (rob_val__20),
  .rob_val__19                       (rob_val__19),
  .rob_val__18                       (rob_val__18),
  .rob_val__17                       (rob_val__17),
  .rob_val__16                       (rob_val__16),
  .rob_val__15                       (rob_val__15),
  .rob_val__14                       (rob_val__14),
  .rob_val__13                       (rob_val__13),
  .rob_val__12                       (rob_val__12),
  .rob_val__11                       (rob_val__11),
  .rob_val__10                       (rob_val__10),
  .rob_val__9                        (rob_val__9),
  .rob_val__8                        (rob_val__8),
  .rob_val__7                        (rob_val__7),
  .rob_val__6                        (rob_val__6),
  .rob_val__5                        (rob_val__5),
  .rob_val__4                        (rob_val__4),
  .rob_val__3                        (rob_val__3),
  .rob_val__2                        (rob_val__2),
  .rob_val__1                        (rob_val__1),
  .rob_val__0                        (rob_val__0),
  .io_enq_uops_0_rob_idx             (io_enq_uops_0_rob_idx),
  ._GEN                              (io_lsu_clr_bsy_0_bits[6:2]),
  .rob_bsy__31                       (rob_bsy__31),
  .rob_bsy__30                       (rob_bsy__30),
  .rob_bsy__29                       (rob_bsy__29),
  .rob_bsy__28                       (rob_bsy__28),
  .rob_bsy__27                       (rob_bsy__27),
  .rob_bsy__26                       (rob_bsy__26),
  .rob_bsy__25                       (rob_bsy__25),
  .rob_bsy__24                       (rob_bsy__24),
  .rob_bsy__23                       (rob_bsy__23),
  .rob_bsy__22                       (rob_bsy__22),
  .rob_bsy__21                       (rob_bsy__21),
  .rob_bsy__20                       (rob_bsy__20),
  .rob_bsy__19                       (rob_bsy__19),
  .rob_bsy__18                       (rob_bsy__18),
  .rob_bsy__17                       (rob_bsy__17),
  .rob_bsy__16                       (rob_bsy__16),
  .rob_bsy__15                       (rob_bsy__15),
  .rob_bsy__14                       (rob_bsy__14),
  .rob_bsy__13                       (rob_bsy__13),
  .rob_bsy__12                       (rob_bsy__12),
  .rob_bsy__11                       (rob_bsy__11),
  .rob_bsy__10                       (rob_bsy__10),
  .rob_bsy__9                        (rob_bsy__9),
  .rob_bsy__8                        (rob_bsy__8),
  .rob_bsy__7                        (rob_bsy__7),
  .rob_bsy__6                        (rob_bsy__6),
  .rob_bsy__5                        (rob_bsy__5),
  .rob_bsy__4                        (rob_bsy__4),
  .rob_bsy__3                        (rob_bsy__3),
  .rob_bsy__2                        (rob_bsy__2),
  .rob_bsy__1                        (rob_bsy__1),
  .rob_bsy__0                        (rob_bsy__0),
  ._GEN_0                            (io_lsu_clr_bsy_1_bits[6:2]),
  ._GEN_1                            (io_lsu_clr_bsy_2_bits[6:2]),
  ._GEN_2                            (io_lxcpt_bits_uop_rob_idx[6:2]),
  .clock                             (clock),
  ._GEN_3                            (_GEN_769),
  ._GEN_4                            (_GEN_641),
  ._GEN_5                            (_GEN_513),
  ._GEN_6                            (_GEN_385),
  ._GEN_7                            (_GEN_257),
  ._GEN_8                            (_GEN_129),
  ._GEN_9                            (_GEN_33),
  .io_enq_uops_0_uses_ldq            (io_enq_uops_0_uses_ldq),
  .io_enq_uops_0_is_br               (io_enq_uops_0_is_br),
  .io_enq_uops_0_is_jalr             (io_enq_uops_0_is_jalr),
  .io_enq_uops_0_uses_stq            (io_enq_uops_0_uses_stq),
  .io_enq_uops_0_is_fence            (io_enq_uops_0_is_fence),
  ._GEN_10                           (_GEN_97),
  ._GEN_11                           (_GEN_131),
  ._GEN_12                           (_GEN_225),
  ._GEN_13                           (_GEN_259),
  ._GEN_14                           (_GEN_353),
  ._GEN_15                           (_GEN_387),
  ._GEN_16                           (_GEN_481),
  ._GEN_17                           (_GEN_515),
  ._GEN_18                           (_GEN_609),
  ._GEN_19                           (_GEN_643),
  ._GEN_20                           (_GEN_737),
  ._GEN_21                           (_GEN_771),
  ._GEN_22                           (_GEN_865),
  ._GEN_23                           (_GEN_34),
  ._GEN_24                           (_GEN_98),
  ._GEN_25                           (_GEN_133),
  ._GEN_26                           (_GEN_226),
  ._GEN_27                           (_GEN_261),
  ._GEN_28                           (_GEN_354),
  ._GEN_29                           (_GEN_389),
  ._GEN_30                           (_GEN_482),
  ._GEN_31                           (_GEN_517),
  ._GEN_32                           (_GEN_610),
  ._GEN_33                           (_GEN_645),
  ._GEN_34                           (_GEN_738),
  ._GEN_35                           (_GEN_773),
  ._GEN_36                           (_GEN_866),
  ._GEN_37                           (_GEN_35),
  ._GEN_38                           (_GEN_99),
  ._GEN_39                           (_GEN_135),
  ._GEN_40                           (_GEN_227),
  ._GEN_41                           (_GEN_263),
  ._GEN_42                           (_GEN_355),
  ._GEN_43                           (_GEN_391),
  ._GEN_44                           (_GEN_483),
  ._GEN_45                           (_GEN_519),
  ._GEN_46                           (_GEN_611),
  ._GEN_47                           (_GEN_647),
  ._GEN_48                           (_GEN_739),
  ._GEN_49                           (_GEN_775),
  ._GEN_50                           (_GEN_867),
  ._GEN_51                           (_GEN_36),
  ._GEN_52                           (_GEN_100),
  ._GEN_53                           (_GEN_137),
  ._GEN_54                           (_GEN_228),
  ._GEN_55                           (_GEN_265),
  ._GEN_56                           (_GEN_356),
  ._GEN_57                           (_GEN_393),
  ._GEN_58                           (_GEN_484),
  ._GEN_59                           (_GEN_521),
  ._GEN_60                           (_GEN_612),
  ._GEN_61                           (_GEN_649),
  ._GEN_62                           (_GEN_740),
  ._GEN_63                           (_GEN_777),
  ._GEN_64                           (_GEN_868),
  ._GEN_65                           (_GEN_37),
  ._GEN_66                           (_GEN_101),
  ._GEN_67                           (_GEN_139),
  ._GEN_68                           (_GEN_229),
  ._GEN_69                           (_GEN_267),
  ._GEN_70                           (_GEN_357),
  ._GEN_71                           (_GEN_395),
  ._GEN_72                           (_GEN_485),
  ._GEN_73                           (_GEN_523),
  ._GEN_74                           (_GEN_613),
  ._GEN_75                           (_GEN_651),
  ._GEN_76                           (_GEN_741),
  ._GEN_77                           (_GEN_779),
  ._GEN_78                           (_GEN_869),
  ._GEN_79                           (_GEN_38),
  ._GEN_80                           (_GEN_102),
  ._GEN_81                           (_GEN_141),
  ._GEN_82                           (_GEN_230),
  ._GEN_83                           (_GEN_269),
  ._GEN_84                           (_GEN_358),
  ._GEN_85                           (_GEN_397),
  ._GEN_86                           (_GEN_486),
  ._GEN_87                           (_GEN_525),
  ._GEN_88                           (_GEN_614),
  ._GEN_89                           (_GEN_653),
  ._GEN_90                           (_GEN_742),
  ._GEN_91                           (_GEN_781),
  ._GEN_92                           (_GEN_870),
  ._GEN_93                           (_GEN_39),
  ._GEN_94                           (_GEN_103),
  ._GEN_95                           (_GEN_143),
  ._GEN_96                           (_GEN_231),
  ._GEN_97                           (_GEN_271),
  ._GEN_98                           (_GEN_359),
  ._GEN_99                           (_GEN_399),
  ._GEN_100                          (_GEN_487),
  ._GEN_101                          (_GEN_527),
  ._GEN_102                          (_GEN_615),
  ._GEN_103                          (_GEN_655),
  ._GEN_104                          (_GEN_743),
  ._GEN_105                          (_GEN_783),
  ._GEN_106                          (_GEN_871),
  ._GEN_107                          (_GEN_40),
  ._GEN_108                          (_GEN_104),
  ._GEN_109                          (_GEN_145),
  ._GEN_110                          (_GEN_232),
  ._GEN_111                          (_GEN_273),
  ._GEN_112                          (_GEN_360),
  ._GEN_113                          (_GEN_401),
  ._GEN_114                          (_GEN_488),
  ._GEN_115                          (_GEN_529),
  ._GEN_116                          (_GEN_616),
  ._GEN_117                          (_GEN_657),
  ._GEN_118                          (_GEN_744),
  ._GEN_119                          (_GEN_785),
  ._GEN_120                          (_GEN_872),
  ._GEN_121                          (_GEN_41),
  ._GEN_122                          (_GEN_105),
  ._GEN_123                          (_GEN_147),
  ._GEN_124                          (_GEN_233),
  ._GEN_125                          (_GEN_275),
  ._GEN_126                          (_GEN_361),
  ._GEN_127                          (_GEN_403),
  ._GEN_128                          (_GEN_489),
  ._GEN_129                          (_GEN_531),
  ._GEN_130                          (_GEN_617),
  ._GEN_131                          (_GEN_659),
  ._GEN_132                          (_GEN_745),
  ._GEN_133                          (_GEN_787),
  ._GEN_134                          (_GEN_873),
  ._GEN_135                          (_GEN_42),
  ._GEN_136                          (_GEN_106),
  ._GEN_137                          (_GEN_149),
  ._GEN_138                          (_GEN_234),
  ._GEN_139                          (_GEN_277),
  ._GEN_140                          (_GEN_362),
  ._GEN_141                          (_GEN_405),
  ._GEN_142                          (_GEN_490),
  ._GEN_143                          (_GEN_533),
  ._GEN_144                          (_GEN_618),
  ._GEN_145                          (_GEN_661),
  ._GEN_146                          (_GEN_746),
  ._GEN_147                          (_GEN_789),
  ._GEN_148                          (_GEN_874),
  ._GEN_149                          (_GEN_43),
  ._GEN_150                          (_GEN_107),
  ._GEN_151                          (_GEN_151),
  ._GEN_152                          (_GEN_235),
  ._GEN_153                          (_GEN_279),
  ._GEN_154                          (_GEN_363),
  ._GEN_155                          (_GEN_407),
  ._GEN_156                          (_GEN_491),
  ._GEN_157                          (_GEN_535),
  ._GEN_158                          (_GEN_619),
  ._GEN_159                          (_GEN_663),
  ._GEN_160                          (_GEN_747),
  ._GEN_161                          (_GEN_791),
  ._GEN_162                          (_GEN_875),
  ._GEN_163                          (_GEN_44),
  ._GEN_164                          (_GEN_108),
  ._GEN_165                          (_GEN_153),
  ._GEN_166                          (_GEN_236),
  ._GEN_167                          (_GEN_281),
  ._GEN_168                          (_GEN_364),
  ._GEN_169                          (_GEN_409),
  ._GEN_170                          (_GEN_492),
  ._GEN_171                          (_GEN_537),
  ._GEN_172                          (_GEN_620),
  ._GEN_173                          (_GEN_665),
  ._GEN_174                          (_GEN_748),
  ._GEN_175                          (_GEN_793),
  ._GEN_176                          (_GEN_876),
  ._GEN_177                          (_GEN_45),
  ._GEN_178                          (_GEN_109),
  ._GEN_179                          (_GEN_155),
  ._GEN_180                          (_GEN_237),
  ._GEN_181                          (_GEN_283),
  ._GEN_182                          (_GEN_365),
  ._GEN_183                          (_GEN_411),
  ._GEN_184                          (_GEN_493),
  ._GEN_185                          (_GEN_539),
  ._GEN_186                          (_GEN_621),
  ._GEN_187                          (_GEN_667),
  ._GEN_188                          (_GEN_749),
  ._GEN_189                          (_GEN_795),
  ._GEN_190                          (_GEN_877),
  ._GEN_191                          (_GEN_46),
  ._GEN_192                          (_GEN_110),
  ._GEN_193                          (_GEN_157),
  ._GEN_194                          (_GEN_238),
  ._GEN_195                          (_GEN_285),
  ._GEN_196                          (_GEN_366),
  ._GEN_197                          (_GEN_413),
  ._GEN_198                          (_GEN_494),
  ._GEN_199                          (_GEN_541),
  ._GEN_200                          (_GEN_622),
  ._GEN_201                          (_GEN_669),
  ._GEN_202                          (_GEN_750),
  ._GEN_203                          (_GEN_797),
  ._GEN_204                          (_GEN_878),
  ._GEN_205                          (_GEN_47),
  ._GEN_206                          (_GEN_111),
  ._GEN_207                          (_GEN_159),
  ._GEN_208                          (_GEN_239),
  ._GEN_209                          (_GEN_287),
  ._GEN_210                          (_GEN_367),
  ._GEN_211                          (_GEN_415),
  ._GEN_212                          (_GEN_495),
  ._GEN_213                          (_GEN_543),
  ._GEN_214                          (_GEN_623),
  ._GEN_215                          (_GEN_671),
  ._GEN_216                          (_GEN_751),
  ._GEN_217                          (_GEN_799),
  ._GEN_218                          (_GEN_879),
  ._GEN_219                          (_GEN_48),
  ._GEN_220                          (_GEN_112),
  ._GEN_221                          (_GEN_161),
  ._GEN_222                          (_GEN_240),
  ._GEN_223                          (_GEN_289),
  ._GEN_224                          (_GEN_368),
  ._GEN_225                          (_GEN_417),
  ._GEN_226                          (_GEN_496),
  ._GEN_227                          (_GEN_545),
  ._GEN_228                          (_GEN_624),
  ._GEN_229                          (_GEN_673),
  ._GEN_230                          (_GEN_752),
  ._GEN_231                          (_GEN_801),
  ._GEN_232                          (_GEN_880),
  ._GEN_233                          (_GEN_49),
  ._GEN_234                          (_GEN_113),
  ._GEN_235                          (_GEN_163),
  ._GEN_236                          (_GEN_241),
  ._GEN_237                          (_GEN_291),
  ._GEN_238                          (_GEN_369),
  ._GEN_239                          (_GEN_419),
  ._GEN_240                          (_GEN_497),
  ._GEN_241                          (_GEN_547),
  ._GEN_242                          (_GEN_625),
  ._GEN_243                          (_GEN_675),
  ._GEN_244                          (_GEN_753),
  ._GEN_245                          (_GEN_803),
  ._GEN_246                          (_GEN_881),
  ._GEN_247                          (_GEN_50),
  ._GEN_248                          (_GEN_114),
  ._GEN_249                          (_GEN_165),
  ._GEN_250                          (_GEN_242),
  ._GEN_251                          (_GEN_293),
  ._GEN_252                          (_GEN_370),
  ._GEN_253                          (_GEN_421),
  ._GEN_254                          (_GEN_498),
  ._GEN_255                          (_GEN_549),
  ._GEN_256                          (_GEN_626),
  ._GEN_257                          (_GEN_677),
  ._GEN_258                          (_GEN_754),
  ._GEN_259                          (_GEN_805),
  ._GEN_260                          (_GEN_882),
  ._GEN_261                          (_GEN_51),
  ._GEN_262                          (_GEN_115),
  ._GEN_263                          (_GEN_167),
  ._GEN_264                          (_GEN_243),
  ._GEN_265                          (_GEN_295),
  ._GEN_266                          (_GEN_371),
  ._GEN_267                          (_GEN_423),
  ._GEN_268                          (_GEN_499),
  ._GEN_269                          (_GEN_551),
  ._GEN_270                          (_GEN_627),
  ._GEN_271                          (_GEN_679),
  ._GEN_272                          (_GEN_755),
  ._GEN_273                          (_GEN_807),
  ._GEN_274                          (_GEN_883),
  ._GEN_275                          (_GEN_52),
  ._GEN_276                          (_GEN_116),
  ._GEN_277                          (_GEN_169),
  ._GEN_278                          (_GEN_244),
  ._GEN_279                          (_GEN_297),
  ._GEN_280                          (_GEN_372),
  ._GEN_281                          (_GEN_425),
  ._GEN_282                          (_GEN_500),
  ._GEN_283                          (_GEN_553),
  ._GEN_284                          (_GEN_628),
  ._GEN_285                          (_GEN_681),
  ._GEN_286                          (_GEN_756),
  ._GEN_287                          (_GEN_809),
  ._GEN_288                          (_GEN_884),
  ._GEN_289                          (_GEN_53),
  ._GEN_290                          (_GEN_117),
  ._GEN_291                          (_GEN_171),
  ._GEN_292                          (_GEN_245),
  ._GEN_293                          (_GEN_299),
  ._GEN_294                          (_GEN_373),
  ._GEN_295                          (_GEN_427),
  ._GEN_296                          (_GEN_501),
  ._GEN_297                          (_GEN_555),
  ._GEN_298                          (_GEN_629),
  ._GEN_299                          (_GEN_683),
  ._GEN_300                          (_GEN_757),
  ._GEN_301                          (_GEN_811),
  ._GEN_302                          (_GEN_885),
  ._GEN_303                          (_GEN_54),
  ._GEN_304                          (_GEN_118),
  ._GEN_305                          (_GEN_173),
  ._GEN_306                          (_GEN_246),
  ._GEN_307                          (_GEN_301),
  ._GEN_308                          (_GEN_374),
  ._GEN_309                          (_GEN_429),
  ._GEN_310                          (_GEN_502),
  ._GEN_311                          (_GEN_557),
  ._GEN_312                          (_GEN_630),
  ._GEN_313                          (_GEN_685),
  ._GEN_314                          (_GEN_758),
  ._GEN_315                          (_GEN_813),
  ._GEN_316                          (_GEN_886),
  ._GEN_317                          (_GEN_55),
  ._GEN_318                          (_GEN_119),
  ._GEN_319                          (_GEN_175),
  ._GEN_320                          (_GEN_247),
  ._GEN_321                          (_GEN_303),
  ._GEN_322                          (_GEN_375),
  ._GEN_323                          (_GEN_431),
  ._GEN_324                          (_GEN_503),
  ._GEN_325                          (_GEN_559),
  ._GEN_326                          (_GEN_631),
  ._GEN_327                          (_GEN_687),
  ._GEN_328                          (_GEN_759),
  ._GEN_329                          (_GEN_815),
  ._GEN_330                          (_GEN_887),
  ._GEN_331                          (_GEN_56),
  ._GEN_332                          (_GEN_120),
  ._GEN_333                          (_GEN_177),
  ._GEN_334                          (_GEN_248),
  ._GEN_335                          (_GEN_305),
  ._GEN_336                          (_GEN_376),
  ._GEN_337                          (_GEN_433),
  ._GEN_338                          (_GEN_504),
  ._GEN_339                          (_GEN_561),
  ._GEN_340                          (_GEN_632),
  ._GEN_341                          (_GEN_689),
  ._GEN_342                          (_GEN_760),
  ._GEN_343                          (_GEN_817),
  ._GEN_344                          (_GEN_888),
  ._GEN_345                          (_GEN_57),
  ._GEN_346                          (_GEN_121),
  ._GEN_347                          (_GEN_179),
  ._GEN_348                          (_GEN_249),
  ._GEN_349                          (_GEN_307),
  ._GEN_350                          (_GEN_377),
  ._GEN_351                          (_GEN_435),
  ._GEN_352                          (_GEN_505),
  ._GEN_353                          (_GEN_563),
  ._GEN_354                          (_GEN_633),
  ._GEN_355                          (_GEN_691),
  ._GEN_356                          (_GEN_761),
  ._GEN_357                          (_GEN_819),
  ._GEN_358                          (_GEN_889),
  ._GEN_359                          (_GEN_58),
  ._GEN_360                          (_GEN_122),
  ._GEN_361                          (_GEN_181),
  ._GEN_362                          (_GEN_250),
  ._GEN_363                          (_GEN_309),
  ._GEN_364                          (_GEN_378),
  ._GEN_365                          (_GEN_437),
  ._GEN_366                          (_GEN_506),
  ._GEN_367                          (_GEN_565),
  ._GEN_368                          (_GEN_634),
  ._GEN_369                          (_GEN_693),
  ._GEN_370                          (_GEN_762),
  ._GEN_371                          (_GEN_821),
  ._GEN_372                          (_GEN_890),
  ._GEN_373                          (_GEN_59),
  ._GEN_374                          (_GEN_123),
  ._GEN_375                          (_GEN_183),
  ._GEN_376                          (_GEN_251),
  ._GEN_377                          (_GEN_311),
  ._GEN_378                          (_GEN_379),
  ._GEN_379                          (_GEN_439),
  ._GEN_380                          (_GEN_507),
  ._GEN_381                          (_GEN_567),
  ._GEN_382                          (_GEN_635),
  ._GEN_383                          (_GEN_695),
  ._GEN_384                          (_GEN_763),
  ._GEN_385                          (_GEN_823),
  ._GEN_386                          (_GEN_891),
  ._GEN_387                          (_GEN_60),
  ._GEN_388                          (_GEN_124),
  ._GEN_389                          (_GEN_185),
  ._GEN_390                          (_GEN_252),
  ._GEN_391                          (_GEN_313),
  ._GEN_392                          (_GEN_380),
  ._GEN_393                          (_GEN_441),
  ._GEN_394                          (_GEN_508),
  ._GEN_395                          (_GEN_569),
  ._GEN_396                          (_GEN_636),
  ._GEN_397                          (_GEN_697),
  ._GEN_398                          (_GEN_764),
  ._GEN_399                          (_GEN_825),
  ._GEN_400                          (_GEN_892),
  ._GEN_401                          (_GEN_61),
  ._GEN_402                          (_GEN_125),
  ._GEN_403                          (_GEN_187),
  ._GEN_404                          (_GEN_253),
  ._GEN_405                          (_GEN_315),
  ._GEN_406                          (_GEN_381),
  ._GEN_407                          (_GEN_443),
  ._GEN_408                          (_GEN_509),
  ._GEN_409                          (_GEN_571),
  ._GEN_410                          (_GEN_637),
  ._GEN_411                          (_GEN_699),
  ._GEN_412                          (_GEN_765),
  ._GEN_413                          (_GEN_827),
  ._GEN_414                          (_GEN_893),
  ._GEN_415                          (_GEN_62),
  ._GEN_416                          (_GEN_126),
  ._GEN_417                          (_GEN_189),
  ._GEN_418                          (_GEN_254),
  ._GEN_419                          (_GEN_317),
  ._GEN_420                          (_GEN_382),
  ._GEN_421                          (_GEN_445),
  ._GEN_422                          (_GEN_510),
  ._GEN_423                          (_GEN_573),
  ._GEN_424                          (_GEN_638),
  ._GEN_425                          (_GEN_701),
  ._GEN_426                          (_GEN_766),
  ._GEN_427                          (_GEN_829),
  ._GEN_428                          (_GEN_894),
  ._GEN_429                          (_GEN_63),
  ._GEN_430                          (_GEN_127),
  ._GEN_431                          (_GEN_191),
  ._GEN_432                          (_GEN_255),
  ._GEN_433                          (_GEN_319),
  ._GEN_434                          (_GEN_383),
  ._GEN_435                          (_GEN_447),
  ._GEN_436                          (_GEN_511),
  ._GEN_437                          (_GEN_575),
  ._GEN_438                          (_GEN_639),
  ._GEN_439                          (_GEN_703),
  ._GEN_440                          (_GEN_767),
  ._GEN_441                          (_GEN_831),
  ._GEN_442                          (_GEN_895),
  ._GEN_443                          (_GEN_64),
  ._GEN_444                          (_GEN_128),
  ._GEN_445                          (_GEN_192),
  ._GEN_446                          (_GEN_256),
  ._GEN_447                          (_GEN_320),
  ._GEN_448                          (_GEN_384),
  ._GEN_449                          (_GEN_448),
  ._GEN_450                          (_GEN_512),
  ._GEN_451                          (_GEN_576),
  ._GEN_452                          (_GEN_640),
  ._GEN_453                          (_GEN_704),
  ._GEN_454                          (_GEN_768),
  ._GEN_455                          (_GEN_832),
  ._GEN_456                          (_GEN_896),
  ._io_commit_rbk_valids_0_output    (_io_commit_rbk_valids_0_output),
  ._io_commit_rbk_valids_1_output    (_io_commit_rbk_valids_1_output),
  ._io_commit_rbk_valids_2_output    (_io_commit_rbk_valids_2_output),
  ._io_commit_rbk_valids_3_output    (_io_commit_rbk_valids_3_output),
  ._io_commit_valids_0_output        (_io_commit_valids_0_output),
  ._io_commit_valids_1_output        (_io_commit_valids_1_output),
  ._io_commit_valids_2_output        (_io_commit_valids_2_output),
  ._io_commit_valids_3_output        (_io_commit_valids_3_output),
  ._GEN_457                          (_GEN_65),
  ._temp_uop_T_61                    (io_wb_resps_0_bits_uop_rob_idx[6:2]),
  .io_wb_resps_0_bits_uop_pdst       (io_wb_resps_0_bits_uop_pdst),
  .rob_uop__31_pdst                  (rob_uop__31_pdst),
  .rob_uop__30_pdst                  (rob_uop__30_pdst),
  .rob_uop__29_pdst                  (rob_uop__29_pdst),
  .rob_uop__28_pdst                  (rob_uop__28_pdst),
  .rob_uop__27_pdst                  (rob_uop__27_pdst),
  .rob_uop__26_pdst                  (rob_uop__26_pdst),
  .rob_uop__25_pdst                  (rob_uop__25_pdst),
  .rob_uop__24_pdst                  (rob_uop__24_pdst),
  .rob_uop__23_pdst                  (rob_uop__23_pdst),
  .rob_uop__22_pdst                  (rob_uop__22_pdst),
  .rob_uop__21_pdst                  (rob_uop__21_pdst),
  .rob_uop__20_pdst                  (rob_uop__20_pdst),
  .rob_uop__19_pdst                  (rob_uop__19_pdst),
  .rob_uop__18_pdst                  (rob_uop__18_pdst),
  .rob_uop__17_pdst                  (rob_uop__17_pdst),
  .rob_uop__16_pdst                  (rob_uop__16_pdst),
  .rob_uop__15_pdst                  (rob_uop__15_pdst),
  .rob_uop__14_pdst                  (rob_uop__14_pdst),
  .rob_uop__13_pdst                  (rob_uop__13_pdst),
  .rob_uop__12_pdst                  (rob_uop__12_pdst),
  .rob_uop__11_pdst                  (rob_uop__11_pdst),
  .rob_uop__10_pdst                  (rob_uop__10_pdst),
  .rob_uop__9_pdst                   (rob_uop__9_pdst),
  .rob_uop__8_pdst                   (rob_uop__8_pdst),
  .rob_uop__7_pdst                   (rob_uop__7_pdst),
  .rob_uop__6_pdst                   (rob_uop__6_pdst),
  .rob_uop__5_pdst                   (rob_uop__5_pdst),
  .rob_uop__4_pdst                   (rob_uop__4_pdst),
  .rob_uop__3_pdst                   (rob_uop__3_pdst),
  .rob_uop__2_pdst                   (rob_uop__2_pdst),
  .rob_uop__1_pdst                   (rob_uop__1_pdst),
  .rob_uop__0_pdst                   (rob_uop__0_pdst),
  .rob_uop__31_ldst_val              (rob_uop__31_ldst_val),
  .rob_uop__30_ldst_val              (rob_uop__30_ldst_val),
  .rob_uop__29_ldst_val              (rob_uop__29_ldst_val),
  .rob_uop__28_ldst_val              (rob_uop__28_ldst_val),
  .rob_uop__27_ldst_val              (rob_uop__27_ldst_val),
  .rob_uop__26_ldst_val              (rob_uop__26_ldst_val),
  .rob_uop__25_ldst_val              (rob_uop__25_ldst_val),
  .rob_uop__24_ldst_val              (rob_uop__24_ldst_val),
  .rob_uop__23_ldst_val              (rob_uop__23_ldst_val),
  .rob_uop__22_ldst_val              (rob_uop__22_ldst_val),
  .rob_uop__21_ldst_val              (rob_uop__21_ldst_val),
  .rob_uop__20_ldst_val              (rob_uop__20_ldst_val),
  .rob_uop__19_ldst_val              (rob_uop__19_ldst_val),
  .rob_uop__18_ldst_val              (rob_uop__18_ldst_val),
  .rob_uop__17_ldst_val              (rob_uop__17_ldst_val),
  .rob_uop__16_ldst_val              (rob_uop__16_ldst_val),
  .rob_uop__15_ldst_val              (rob_uop__15_ldst_val),
  .rob_uop__14_ldst_val              (rob_uop__14_ldst_val),
  .rob_uop__13_ldst_val              (rob_uop__13_ldst_val),
  .rob_uop__12_ldst_val              (rob_uop__12_ldst_val),
  .rob_uop__11_ldst_val              (rob_uop__11_ldst_val),
  .rob_uop__10_ldst_val              (rob_uop__10_ldst_val),
  .rob_uop__9_ldst_val               (rob_uop__9_ldst_val),
  .rob_uop__8_ldst_val               (rob_uop__8_ldst_val),
  .rob_uop__7_ldst_val               (rob_uop__7_ldst_val),
  .rob_uop__6_ldst_val               (rob_uop__6_ldst_val),
  .rob_uop__5_ldst_val               (rob_uop__5_ldst_val),
  .rob_uop__4_ldst_val               (rob_uop__4_ldst_val),
  .rob_uop__3_ldst_val               (rob_uop__3_ldst_val),
  .rob_uop__2_ldst_val               (rob_uop__2_ldst_val),
  .rob_uop__1_ldst_val               (rob_uop__1_ldst_val),
  .rob_uop__0_ldst_val               (rob_uop__0_ldst_val),
  ._temp_uop_T_63                    (io_wb_resps_1_bits_uop_rob_idx[6:2]),
  .io_wb_resps_1_bits_uop_pdst       (io_wb_resps_1_bits_uop_pdst),
  ._GEN_458                          (_GEN_193),
  ._temp_uop_T_65                    (io_wb_resps_2_bits_uop_rob_idx[6:2]),
  .io_wb_resps_2_bits_uop_pdst       (io_wb_resps_2_bits_uop_pdst),
  ._temp_uop_T_67                    (io_wb_resps_3_bits_uop_rob_idx[6:2]),
  .io_wb_resps_3_bits_uop_pdst       (io_wb_resps_3_bits_uop_pdst),
  ._GEN_459                          (_GEN_321),
  ._temp_uop_T_69                    (io_wb_resps_4_bits_uop_rob_idx[6:2]),
  .io_wb_resps_4_bits_uop_pdst       (io_wb_resps_4_bits_uop_pdst),
  ._temp_uop_T_71                    (io_wb_resps_5_bits_uop_rob_idx[6:2]),
  .io_wb_resps_5_bits_uop_pdst       (io_wb_resps_5_bits_uop_pdst),
  ._GEN_460                          (_GEN_449),
  ._temp_uop_T_73                    (io_wb_resps_6_bits_uop_rob_idx[6:2]),
  .io_wb_resps_6_bits_uop_pdst       (io_wb_resps_6_bits_uop_pdst),
  ._temp_uop_T_75                    (io_wb_resps_7_bits_uop_rob_idx[6:2]),
  .io_wb_resps_7_bits_uop_pdst       (io_wb_resps_7_bits_uop_pdst),
  ._GEN_461                          (_GEN_577),
  ._temp_uop_T_77                    (io_wb_resps_8_bits_uop_rob_idx[6:2]),
  .io_wb_resps_8_bits_uop_pdst       (io_wb_resps_8_bits_uop_pdst),
  ._temp_uop_T_79                    (io_wb_resps_9_bits_uop_rob_idx[6:2]),
  .io_wb_resps_9_bits_uop_pdst       (io_wb_resps_9_bits_uop_pdst),
  .rob_val_1_31                      (rob_val_1_31),
  .rob_val_1_30                      (rob_val_1_30),
  .rob_val_1_29                      (rob_val_1_29),
  .rob_val_1_28                      (rob_val_1_28),
  .rob_val_1_27                      (rob_val_1_27),
  .rob_val_1_26                      (rob_val_1_26),
  .rob_val_1_25                      (rob_val_1_25),
  .rob_val_1_24                      (rob_val_1_24),
  .rob_val_1_23                      (rob_val_1_23),
  .rob_val_1_22                      (rob_val_1_22),
  .rob_val_1_21                      (rob_val_1_21),
  .rob_val_1_20                      (rob_val_1_20),
  .rob_val_1_19                      (rob_val_1_19),
  .rob_val_1_18                      (rob_val_1_18),
  .rob_val_1_17                      (rob_val_1_17),
  .rob_val_1_16                      (rob_val_1_16),
  .rob_val_1_15                      (rob_val_1_15),
  .rob_val_1_14                      (rob_val_1_14),
  .rob_val_1_13                      (rob_val_1_13),
  .rob_val_1_12                      (rob_val_1_12),
  .rob_val_1_11                      (rob_val_1_11),
  .rob_val_1_10                      (rob_val_1_10),
  .rob_val_1_9                       (rob_val_1_9),
  .rob_val_1_8                       (rob_val_1_8),
  .rob_val_1_7                       (rob_val_1_7),
  .rob_val_1_6                       (rob_val_1_6),
  .rob_val_1_5                       (rob_val_1_5),
  .rob_val_1_4                       (rob_val_1_4),
  .rob_val_1_3                       (rob_val_1_3),
  .rob_val_1_2                       (rob_val_1_2),
  .rob_val_1_1                       (rob_val_1_1),
  .rob_val_1_0                       (rob_val_1_0),
  .io_enq_uops_1_rob_idx             (io_enq_uops_1_rob_idx),
  .rob_bsy_1_31                      (rob_bsy_1_31),
  .rob_bsy_1_30                      (rob_bsy_1_30),
  .rob_bsy_1_29                      (rob_bsy_1_29),
  .rob_bsy_1_28                      (rob_bsy_1_28),
  .rob_bsy_1_27                      (rob_bsy_1_27),
  .rob_bsy_1_26                      (rob_bsy_1_26),
  .rob_bsy_1_25                      (rob_bsy_1_25),
  .rob_bsy_1_24                      (rob_bsy_1_24),
  .rob_bsy_1_23                      (rob_bsy_1_23),
  .rob_bsy_1_22                      (rob_bsy_1_22),
  .rob_bsy_1_21                      (rob_bsy_1_21),
  .rob_bsy_1_20                      (rob_bsy_1_20),
  .rob_bsy_1_19                      (rob_bsy_1_19),
  .rob_bsy_1_18                      (rob_bsy_1_18),
  .rob_bsy_1_17                      (rob_bsy_1_17),
  .rob_bsy_1_16                      (rob_bsy_1_16),
  .rob_bsy_1_15                      (rob_bsy_1_15),
  .rob_bsy_1_14                      (rob_bsy_1_14),
  .rob_bsy_1_13                      (rob_bsy_1_13),
  .rob_bsy_1_12                      (rob_bsy_1_12),
  .rob_bsy_1_11                      (rob_bsy_1_11),
  .rob_bsy_1_10                      (rob_bsy_1_10),
  .rob_bsy_1_9                       (rob_bsy_1_9),
  .rob_bsy_1_8                       (rob_bsy_1_8),
  .rob_bsy_1_7                       (rob_bsy_1_7),
  .rob_bsy_1_6                       (rob_bsy_1_6),
  .rob_bsy_1_5                       (rob_bsy_1_5),
  .rob_bsy_1_4                       (rob_bsy_1_4),
  .rob_bsy_1_3                       (rob_bsy_1_3),
  .rob_bsy_1_2                       (rob_bsy_1_2),
  .rob_bsy_1_1                       (rob_bsy_1_1),
  .rob_bsy_1_0                       (rob_bsy_1_0),
  ._GEN_462                          (_GEN_1293),
  ._GEN_463                          (_GEN_1227),
  ._GEN_464                          (_GEN_1161),
  ._GEN_465                          (_GEN_1095),
  ._GEN_466                          (_GEN_1029),
  ._GEN_467                          (_GEN_963),
  ._GEN_468                          (_GEN_898),
  .io_enq_uops_1_uses_ldq            (io_enq_uops_1_uses_ldq),
  .io_enq_uops_1_is_br               (io_enq_uops_1_is_br),
  .io_enq_uops_1_is_jalr             (io_enq_uops_1_is_jalr),
  .io_enq_uops_1_uses_stq            (io_enq_uops_1_uses_stq),
  .io_enq_uops_1_is_fence            (io_enq_uops_1_is_fence),
  ._GEN_469                          (_GEN_931),
  ._GEN_470                          (_GEN_964),
  ._GEN_471                          (_GEN_997),
  ._GEN_472                          (_GEN_1030),
  ._GEN_473                          (_GEN_1063),
  ._GEN_474                          (_GEN_1096),
  ._GEN_475                          (_GEN_1129),
  ._GEN_476                          (_GEN_1162),
  ._GEN_477                          (_GEN_1195),
  ._GEN_478                          (_GEN_1228),
  ._GEN_479                          (_GEN_1261),
  ._GEN_480                          (_GEN_1294),
  ._GEN_481                          (_GEN_1327),
  ._GEN_482                          (_GEN_899),
  ._GEN_483                          (_GEN_932),
  ._GEN_484                          (_GEN_965),
  ._GEN_485                          (_GEN_998),
  ._GEN_486                          (_GEN_1031),
  ._GEN_487                          (_GEN_1064),
  ._GEN_488                          (_GEN_1097),
  ._GEN_489                          (_GEN_1130),
  ._GEN_490                          (_GEN_1163),
  ._GEN_491                          (_GEN_1196),
  ._GEN_492                          (_GEN_1229),
  ._GEN_493                          (_GEN_1262),
  ._GEN_494                          (_GEN_1295),
  ._GEN_495                          (_GEN_1328),
  ._GEN_496                          (_GEN_900),
  ._GEN_497                          (_GEN_933),
  ._GEN_498                          (_GEN_966),
  ._GEN_499                          (_GEN_999),
  ._GEN_500                          (_GEN_1032),
  ._GEN_501                          (_GEN_1065),
  ._GEN_502                          (_GEN_1098),
  ._GEN_503                          (_GEN_1131),
  ._GEN_504                          (_GEN_1164),
  ._GEN_505                          (_GEN_1197),
  ._GEN_506                          (_GEN_1230),
  ._GEN_507                          (_GEN_1263),
  ._GEN_508                          (_GEN_1296),
  ._GEN_509                          (_GEN_1329),
  ._GEN_510                          (_GEN_901),
  ._GEN_511                          (_GEN_934),
  ._GEN_512                          (_GEN_967),
  ._GEN_513                          (_GEN_1000),
  ._GEN_514                          (_GEN_1033),
  ._GEN_515                          (_GEN_1066),
  ._GEN_516                          (_GEN_1099),
  ._GEN_517                          (_GEN_1132),
  ._GEN_518                          (_GEN_1165),
  ._GEN_519                          (_GEN_1198),
  ._GEN_520                          (_GEN_1231),
  ._GEN_521                          (_GEN_1264),
  ._GEN_522                          (_GEN_1297),
  ._GEN_523                          (_GEN_1330),
  ._GEN_524                          (_GEN_902),
  ._GEN_525                          (_GEN_935),
  ._GEN_526                          (_GEN_968),
  ._GEN_527                          (_GEN_1001),
  ._GEN_528                          (_GEN_1034),
  ._GEN_529                          (_GEN_1067),
  ._GEN_530                          (_GEN_1100),
  ._GEN_531                          (_GEN_1133),
  ._GEN_532                          (_GEN_1166),
  ._GEN_533                          (_GEN_1199),
  ._GEN_534                          (_GEN_1232),
  ._GEN_535                          (_GEN_1265),
  ._GEN_536                          (_GEN_1298),
  ._GEN_537                          (_GEN_1331),
  ._GEN_538                          (_GEN_903),
  ._GEN_539                          (_GEN_936),
  ._GEN_540                          (_GEN_969),
  ._GEN_541                          (_GEN_1002),
  ._GEN_542                          (_GEN_1035),
  ._GEN_543                          (_GEN_1068),
  ._GEN_544                          (_GEN_1101),
  ._GEN_545                          (_GEN_1134),
  ._GEN_546                          (_GEN_1167),
  ._GEN_547                          (_GEN_1200),
  ._GEN_548                          (_GEN_1233),
  ._GEN_549                          (_GEN_1266),
  ._GEN_550                          (_GEN_1299),
  ._GEN_551                          (_GEN_1332),
  ._GEN_552                          (_GEN_904),
  ._GEN_553                          (_GEN_937),
  ._GEN_554                          (_GEN_970),
  ._GEN_555                          (_GEN_1003),
  ._GEN_556                          (_GEN_1036),
  ._GEN_557                          (_GEN_1069),
  ._GEN_558                          (_GEN_1102),
  ._GEN_559                          (_GEN_1135),
  ._GEN_560                          (_GEN_1168),
  ._GEN_561                          (_GEN_1201),
  ._GEN_562                          (_GEN_1234),
  ._GEN_563                          (_GEN_1267),
  ._GEN_564                          (_GEN_1300),
  ._GEN_565                          (_GEN_1333),
  ._GEN_566                          (_GEN_905),
  ._GEN_567                          (_GEN_938),
  ._GEN_568                          (_GEN_971),
  ._GEN_569                          (_GEN_1004),
  ._GEN_570                          (_GEN_1037),
  ._GEN_571                          (_GEN_1070),
  ._GEN_572                          (_GEN_1103),
  ._GEN_573                          (_GEN_1136),
  ._GEN_574                          (_GEN_1169),
  ._GEN_575                          (_GEN_1202),
  ._GEN_576                          (_GEN_1235),
  ._GEN_577                          (_GEN_1268),
  ._GEN_578                          (_GEN_1301),
  ._GEN_579                          (_GEN_1334),
  ._GEN_580                          (_GEN_906),
  ._GEN_581                          (_GEN_939),
  ._GEN_582                          (_GEN_972),
  ._GEN_583                          (_GEN_1005),
  ._GEN_584                          (_GEN_1038),
  ._GEN_585                          (_GEN_1071),
  ._GEN_586                          (_GEN_1104),
  ._GEN_587                          (_GEN_1137),
  ._GEN_588                          (_GEN_1170),
  ._GEN_589                          (_GEN_1203),
  ._GEN_590                          (_GEN_1236),
  ._GEN_591                          (_GEN_1269),
  ._GEN_592                          (_GEN_1302),
  ._GEN_593                          (_GEN_1335),
  ._GEN_594                          (_GEN_907),
  ._GEN_595                          (_GEN_940),
  ._GEN_596                          (_GEN_973),
  ._GEN_597                          (_GEN_1006),
  ._GEN_598                          (_GEN_1039),
  ._GEN_599                          (_GEN_1072),
  ._GEN_600                          (_GEN_1105),
  ._GEN_601                          (_GEN_1138),
  ._GEN_602                          (_GEN_1171),
  ._GEN_603                          (_GEN_1204),
  ._GEN_604                          (_GEN_1237),
  ._GEN_605                          (_GEN_1270),
  ._GEN_606                          (_GEN_1303),
  ._GEN_607                          (_GEN_1336),
  ._GEN_608                          (_GEN_908),
  ._GEN_609                          (_GEN_941),
  ._GEN_610                          (_GEN_974),
  ._GEN_611                          (_GEN_1007),
  ._GEN_612                          (_GEN_1040),
  ._GEN_613                          (_GEN_1073),
  ._GEN_614                          (_GEN_1106),
  ._GEN_615                          (_GEN_1139),
  ._GEN_616                          (_GEN_1172),
  ._GEN_617                          (_GEN_1205),
  ._GEN_618                          (_GEN_1238),
  ._GEN_619                          (_GEN_1271),
  ._GEN_620                          (_GEN_1304),
  ._GEN_621                          (_GEN_1337),
  ._GEN_622                          (_GEN_909),
  ._GEN_623                          (_GEN_942),
  ._GEN_624                          (_GEN_975),
  ._GEN_625                          (_GEN_1008),
  ._GEN_626                          (_GEN_1041),
  ._GEN_627                          (_GEN_1074),
  ._GEN_628                          (_GEN_1107),
  ._GEN_629                          (_GEN_1140),
  ._GEN_630                          (_GEN_1173),
  ._GEN_631                          (_GEN_1206),
  ._GEN_632                          (_GEN_1239),
  ._GEN_633                          (_GEN_1272),
  ._GEN_634                          (_GEN_1305),
  ._GEN_635                          (_GEN_1338),
  ._GEN_636                          (_GEN_910),
  ._GEN_637                          (_GEN_943),
  ._GEN_638                          (_GEN_976),
  ._GEN_639                          (_GEN_1009),
  ._GEN_640                          (_GEN_1042),
  ._GEN_641                          (_GEN_1075),
  ._GEN_642                          (_GEN_1108),
  ._GEN_643                          (_GEN_1141),
  ._GEN_644                          (_GEN_1174),
  ._GEN_645                          (_GEN_1207),
  ._GEN_646                          (_GEN_1240),
  ._GEN_647                          (_GEN_1273),
  ._GEN_648                          (_GEN_1306),
  ._GEN_649                          (_GEN_1339),
  ._GEN_650                          (_GEN_911),
  ._GEN_651                          (_GEN_944),
  ._GEN_652                          (_GEN_977),
  ._GEN_653                          (_GEN_1010),
  ._GEN_654                          (_GEN_1043),
  ._GEN_655                          (_GEN_1076),
  ._GEN_656                          (_GEN_1109),
  ._GEN_657                          (_GEN_1142),
  ._GEN_658                          (_GEN_1175),
  ._GEN_659                          (_GEN_1208),
  ._GEN_660                          (_GEN_1241),
  ._GEN_661                          (_GEN_1274),
  ._GEN_662                          (_GEN_1307),
  ._GEN_663                          (_GEN_1340),
  ._GEN_664                          (_GEN_912),
  ._GEN_665                          (_GEN_945),
  ._GEN_666                          (_GEN_978),
  ._GEN_667                          (_GEN_1011),
  ._GEN_668                          (_GEN_1044),
  ._GEN_669                          (_GEN_1077),
  ._GEN_670                          (_GEN_1110),
  ._GEN_671                          (_GEN_1143),
  ._GEN_672                          (_GEN_1176),
  ._GEN_673                          (_GEN_1209),
  ._GEN_674                          (_GEN_1242),
  ._GEN_675                          (_GEN_1275),
  ._GEN_676                          (_GEN_1308),
  ._GEN_677                          (_GEN_1341),
  ._GEN_678                          (_GEN_913),
  ._GEN_679                          (_GEN_946),
  ._GEN_680                          (_GEN_979),
  ._GEN_681                          (_GEN_1012),
  ._GEN_682                          (_GEN_1045),
  ._GEN_683                          (_GEN_1078),
  ._GEN_684                          (_GEN_1111),
  ._GEN_685                          (_GEN_1144),
  ._GEN_686                          (_GEN_1177),
  ._GEN_687                          (_GEN_1210),
  ._GEN_688                          (_GEN_1243),
  ._GEN_689                          (_GEN_1276),
  ._GEN_690                          (_GEN_1309),
  ._GEN_691                          (_GEN_1342),
  ._GEN_692                          (_GEN_914),
  ._GEN_693                          (_GEN_947),
  ._GEN_694                          (_GEN_980),
  ._GEN_695                          (_GEN_1013),
  ._GEN_696                          (_GEN_1046),
  ._GEN_697                          (_GEN_1079),
  ._GEN_698                          (_GEN_1112),
  ._GEN_699                          (_GEN_1145),
  ._GEN_700                          (_GEN_1178),
  ._GEN_701                          (_GEN_1211),
  ._GEN_702                          (_GEN_1244),
  ._GEN_703                          (_GEN_1277),
  ._GEN_704                          (_GEN_1310),
  ._GEN_705                          (_GEN_1343),
  ._GEN_706                          (_GEN_915),
  ._GEN_707                          (_GEN_948),
  ._GEN_708                          (_GEN_981),
  ._GEN_709                          (_GEN_1014),
  ._GEN_710                          (_GEN_1047),
  ._GEN_711                          (_GEN_1080),
  ._GEN_712                          (_GEN_1113),
  ._GEN_713                          (_GEN_1146),
  ._GEN_714                          (_GEN_1179),
  ._GEN_715                          (_GEN_1212),
  ._GEN_716                          (_GEN_1245),
  ._GEN_717                          (_GEN_1278),
  ._GEN_718                          (_GEN_1311),
  ._GEN_719                          (_GEN_1344),
  ._GEN_720                          (_GEN_916),
  ._GEN_721                          (_GEN_949),
  ._GEN_722                          (_GEN_982),
  ._GEN_723                          (_GEN_1015),
  ._GEN_724                          (_GEN_1048),
  ._GEN_725                          (_GEN_1081),
  ._GEN_726                          (_GEN_1114),
  ._GEN_727                          (_GEN_1147),
  ._GEN_728                          (_GEN_1180),
  ._GEN_729                          (_GEN_1213),
  ._GEN_730                          (_GEN_1246),
  ._GEN_731                          (_GEN_1279),
  ._GEN_732                          (_GEN_1312),
  ._GEN_733                          (_GEN_1345),
  ._GEN_734                          (_GEN_917),
  ._GEN_735                          (_GEN_950),
  ._GEN_736                          (_GEN_983),
  ._GEN_737                          (_GEN_1016),
  ._GEN_738                          (_GEN_1049),
  ._GEN_739                          (_GEN_1082),
  ._GEN_740                          (_GEN_1115),
  ._GEN_741                          (_GEN_1148),
  ._GEN_742                          (_GEN_1181),
  ._GEN_743                          (_GEN_1214),
  ._GEN_744                          (_GEN_1247),
  ._GEN_745                          (_GEN_1280),
  ._GEN_746                          (_GEN_1313),
  ._GEN_747                          (_GEN_1346),
  ._GEN_748                          (_GEN_918),
  ._GEN_749                          (_GEN_951),
  ._GEN_750                          (_GEN_984),
  ._GEN_751                          (_GEN_1017),
  ._GEN_752                          (_GEN_1050),
  ._GEN_753                          (_GEN_1083),
  ._GEN_754                          (_GEN_1116),
  ._GEN_755                          (_GEN_1149),
  ._GEN_756                          (_GEN_1182),
  ._GEN_757                          (_GEN_1215),
  ._GEN_758                          (_GEN_1248),
  ._GEN_759                          (_GEN_1281),
  ._GEN_760                          (_GEN_1314),
  ._GEN_761                          (_GEN_1347),
  ._GEN_762                          (_GEN_919),
  ._GEN_763                          (_GEN_952),
  ._GEN_764                          (_GEN_985),
  ._GEN_765                          (_GEN_1018),
  ._GEN_766                          (_GEN_1051),
  ._GEN_767                          (_GEN_1084),
  ._GEN_768                          (_GEN_1117),
  ._GEN_769                          (_GEN_1150),
  ._GEN_770                          (_GEN_1183),
  ._GEN_771                          (_GEN_1216),
  ._GEN_772                          (_GEN_1249),
  ._GEN_773                          (_GEN_1282),
  ._GEN_774                          (_GEN_1315),
  ._GEN_775                          (_GEN_1348),
  ._GEN_776                          (_GEN_920),
  ._GEN_777                          (_GEN_953),
  ._GEN_778                          (_GEN_986),
  ._GEN_779                          (_GEN_1019),
  ._GEN_780                          (_GEN_1052),
  ._GEN_781                          (_GEN_1085),
  ._GEN_782                          (_GEN_1118),
  ._GEN_783                          (_GEN_1151),
  ._GEN_784                          (_GEN_1184),
  ._GEN_785                          (_GEN_1217),
  ._GEN_786                          (_GEN_1250),
  ._GEN_787                          (_GEN_1283),
  ._GEN_788                          (_GEN_1316),
  ._GEN_789                          (_GEN_1349),
  ._GEN_790                          (_GEN_921),
  ._GEN_791                          (_GEN_954),
  ._GEN_792                          (_GEN_987),
  ._GEN_793                          (_GEN_1020),
  ._GEN_794                          (_GEN_1053),
  ._GEN_795                          (_GEN_1086),
  ._GEN_796                          (_GEN_1119),
  ._GEN_797                          (_GEN_1152),
  ._GEN_798                          (_GEN_1185),
  ._GEN_799                          (_GEN_1218),
  ._GEN_800                          (_GEN_1251),
  ._GEN_801                          (_GEN_1284),
  ._GEN_802                          (_GEN_1317),
  ._GEN_803                          (_GEN_1350),
  ._GEN_804                          (_GEN_922),
  ._GEN_805                          (_GEN_955),
  ._GEN_806                          (_GEN_988),
  ._GEN_807                          (_GEN_1021),
  ._GEN_808                          (_GEN_1054),
  ._GEN_809                          (_GEN_1087),
  ._GEN_810                          (_GEN_1120),
  ._GEN_811                          (_GEN_1153),
  ._GEN_812                          (_GEN_1186),
  ._GEN_813                          (_GEN_1219),
  ._GEN_814                          (_GEN_1252),
  ._GEN_815                          (_GEN_1285),
  ._GEN_816                          (_GEN_1318),
  ._GEN_817                          (_GEN_1351),
  ._GEN_818                          (_GEN_923),
  ._GEN_819                          (_GEN_956),
  ._GEN_820                          (_GEN_989),
  ._GEN_821                          (_GEN_1022),
  ._GEN_822                          (_GEN_1055),
  ._GEN_823                          (_GEN_1088),
  ._GEN_824                          (_GEN_1121),
  ._GEN_825                          (_GEN_1154),
  ._GEN_826                          (_GEN_1187),
  ._GEN_827                          (_GEN_1220),
  ._GEN_828                          (_GEN_1253),
  ._GEN_829                          (_GEN_1286),
  ._GEN_830                          (_GEN_1319),
  ._GEN_831                          (_GEN_1352),
  ._GEN_832                          (_GEN_924),
  ._GEN_833                          (_GEN_957),
  ._GEN_834                          (_GEN_990),
  ._GEN_835                          (_GEN_1023),
  ._GEN_836                          (_GEN_1056),
  ._GEN_837                          (_GEN_1089),
  ._GEN_838                          (_GEN_1122),
  ._GEN_839                          (_GEN_1155),
  ._GEN_840                          (_GEN_1188),
  ._GEN_841                          (_GEN_1221),
  ._GEN_842                          (_GEN_1254),
  ._GEN_843                          (_GEN_1287),
  ._GEN_844                          (_GEN_1320),
  ._GEN_845                          (_GEN_1353),
  ._GEN_846                          (_GEN_925),
  ._GEN_847                          (_GEN_958),
  ._GEN_848                          (_GEN_991),
  ._GEN_849                          (_GEN_1024),
  ._GEN_850                          (_GEN_1057),
  ._GEN_851                          (_GEN_1090),
  ._GEN_852                          (_GEN_1123),
  ._GEN_853                          (_GEN_1156),
  ._GEN_854                          (_GEN_1189),
  ._GEN_855                          (_GEN_1222),
  ._GEN_856                          (_GEN_1255),
  ._GEN_857                          (_GEN_1288),
  ._GEN_858                          (_GEN_1321),
  ._GEN_859                          (_GEN_1354),
  ._GEN_860                          (_GEN_926),
  ._GEN_861                          (_GEN_959),
  ._GEN_862                          (_GEN_992),
  ._GEN_863                          (_GEN_1025),
  ._GEN_864                          (_GEN_1058),
  ._GEN_865                          (_GEN_1091),
  ._GEN_866                          (_GEN_1124),
  ._GEN_867                          (_GEN_1157),
  ._GEN_868                          (_GEN_1190),
  ._GEN_869                          (_GEN_1223),
  ._GEN_870                          (_GEN_1256),
  ._GEN_871                          (_GEN_1289),
  ._GEN_872                          (_GEN_1322),
  ._GEN_873                          (_GEN_1355),
  ._GEN_874                          (_GEN_927),
  ._GEN_875                          (_GEN_960),
  ._GEN_876                          (_GEN_993),
  ._GEN_877                          (_GEN_1026),
  ._GEN_878                          (_GEN_1059),
  ._GEN_879                          (_GEN_1092),
  ._GEN_880                          (_GEN_1125),
  ._GEN_881                          (_GEN_1158),
  ._GEN_882                          (_GEN_1191),
  ._GEN_883                          (_GEN_1224),
  ._GEN_884                          (_GEN_1257),
  ._GEN_885                          (_GEN_1290),
  ._GEN_886                          (_GEN_1323),
  ._GEN_887                          (_GEN_1356),
  ._GEN_888                          (_GEN_928),
  ._GEN_889                          (_GEN_961),
  ._GEN_890                          (_GEN_994),
  ._GEN_891                          (_GEN_1027),
  ._GEN_892                          (_GEN_1060),
  ._GEN_893                          (_GEN_1093),
  ._GEN_894                          (_GEN_1126),
  ._GEN_895                          (_GEN_1159),
  ._GEN_896                          (_GEN_1192),
  ._GEN_897                          (_GEN_1225),
  ._GEN_898                          (_GEN_1258),
  ._GEN_899                          (_GEN_1291),
  ._GEN_900                          (_GEN_1324),
  ._GEN_901                          (_GEN_1357),
  ._GEN_902                          (_GEN_929),
  ._GEN_903                          (_GEN_962),
  ._GEN_904                          (_GEN_995),
  ._GEN_905                          (_GEN_1028),
  ._GEN_906                          (_GEN_1061),
  ._GEN_907                          (_GEN_1094),
  ._GEN_908                          (_GEN_1127),
  ._GEN_909                          (_GEN_1160),
  ._GEN_910                          (_GEN_1193),
  ._GEN_911                          (_GEN_1226),
  ._GEN_912                          (_GEN_1259),
  ._GEN_913                          (_GEN_1292),
  ._GEN_914                          (_GEN_1325),
  ._GEN_915                          (_GEN_1358),
  ._GEN_916                          (_GEN_930),
  .rob_uop_1_31_pdst                 (rob_uop_1_31_pdst),
  .rob_uop_1_30_pdst                 (rob_uop_1_30_pdst),
  .rob_uop_1_29_pdst                 (rob_uop_1_29_pdst),
  .rob_uop_1_28_pdst                 (rob_uop_1_28_pdst),
  .rob_uop_1_27_pdst                 (rob_uop_1_27_pdst),
  .rob_uop_1_26_pdst                 (rob_uop_1_26_pdst),
  .rob_uop_1_25_pdst                 (rob_uop_1_25_pdst),
  .rob_uop_1_24_pdst                 (rob_uop_1_24_pdst),
  .rob_uop_1_23_pdst                 (rob_uop_1_23_pdst),
  .rob_uop_1_22_pdst                 (rob_uop_1_22_pdst),
  .rob_uop_1_21_pdst                 (rob_uop_1_21_pdst),
  .rob_uop_1_20_pdst                 (rob_uop_1_20_pdst),
  .rob_uop_1_19_pdst                 (rob_uop_1_19_pdst),
  .rob_uop_1_18_pdst                 (rob_uop_1_18_pdst),
  .rob_uop_1_17_pdst                 (rob_uop_1_17_pdst),
  .rob_uop_1_16_pdst                 (rob_uop_1_16_pdst),
  .rob_uop_1_15_pdst                 (rob_uop_1_15_pdst),
  .rob_uop_1_14_pdst                 (rob_uop_1_14_pdst),
  .rob_uop_1_13_pdst                 (rob_uop_1_13_pdst),
  .rob_uop_1_12_pdst                 (rob_uop_1_12_pdst),
  .rob_uop_1_11_pdst                 (rob_uop_1_11_pdst),
  .rob_uop_1_10_pdst                 (rob_uop_1_10_pdst),
  .rob_uop_1_9_pdst                  (rob_uop_1_9_pdst),
  .rob_uop_1_8_pdst                  (rob_uop_1_8_pdst),
  .rob_uop_1_7_pdst                  (rob_uop_1_7_pdst),
  .rob_uop_1_6_pdst                  (rob_uop_1_6_pdst),
  .rob_uop_1_5_pdst                  (rob_uop_1_5_pdst),
  .rob_uop_1_4_pdst                  (rob_uop_1_4_pdst),
  .rob_uop_1_3_pdst                  (rob_uop_1_3_pdst),
  .rob_uop_1_2_pdst                  (rob_uop_1_2_pdst),
  .rob_uop_1_1_pdst                  (rob_uop_1_1_pdst),
  .rob_uop_1_0_pdst                  (rob_uop_1_0_pdst),
  .rob_uop_1_31_ldst_val             (rob_uop_1_31_ldst_val),
  .rob_uop_1_30_ldst_val             (rob_uop_1_30_ldst_val),
  .rob_uop_1_29_ldst_val             (rob_uop_1_29_ldst_val),
  .rob_uop_1_28_ldst_val             (rob_uop_1_28_ldst_val),
  .rob_uop_1_27_ldst_val             (rob_uop_1_27_ldst_val),
  .rob_uop_1_26_ldst_val             (rob_uop_1_26_ldst_val),
  .rob_uop_1_25_ldst_val             (rob_uop_1_25_ldst_val),
  .rob_uop_1_24_ldst_val             (rob_uop_1_24_ldst_val),
  .rob_uop_1_23_ldst_val             (rob_uop_1_23_ldst_val),
  .rob_uop_1_22_ldst_val             (rob_uop_1_22_ldst_val),
  .rob_uop_1_21_ldst_val             (rob_uop_1_21_ldst_val),
  .rob_uop_1_20_ldst_val             (rob_uop_1_20_ldst_val),
  .rob_uop_1_19_ldst_val             (rob_uop_1_19_ldst_val),
  .rob_uop_1_18_ldst_val             (rob_uop_1_18_ldst_val),
  .rob_uop_1_17_ldst_val             (rob_uop_1_17_ldst_val),
  .rob_uop_1_16_ldst_val             (rob_uop_1_16_ldst_val),
  .rob_uop_1_15_ldst_val             (rob_uop_1_15_ldst_val),
  .rob_uop_1_14_ldst_val             (rob_uop_1_14_ldst_val),
  .rob_uop_1_13_ldst_val             (rob_uop_1_13_ldst_val),
  .rob_uop_1_12_ldst_val             (rob_uop_1_12_ldst_val),
  .rob_uop_1_11_ldst_val             (rob_uop_1_11_ldst_val),
  .rob_uop_1_10_ldst_val             (rob_uop_1_10_ldst_val),
  .rob_uop_1_9_ldst_val              (rob_uop_1_9_ldst_val),
  .rob_uop_1_8_ldst_val              (rob_uop_1_8_ldst_val),
  .rob_uop_1_7_ldst_val              (rob_uop_1_7_ldst_val),
  .rob_uop_1_6_ldst_val              (rob_uop_1_6_ldst_val),
  .rob_uop_1_5_ldst_val              (rob_uop_1_5_ldst_val),
  .rob_uop_1_4_ldst_val              (rob_uop_1_4_ldst_val),
  .rob_uop_1_3_ldst_val              (rob_uop_1_3_ldst_val),
  .rob_uop_1_2_ldst_val              (rob_uop_1_2_ldst_val),
  .rob_uop_1_1_ldst_val              (rob_uop_1_1_ldst_val),
  .rob_uop_1_0_ldst_val              (rob_uop_1_0_ldst_val),
  ._GEN_917                          (_GEN_996),
  ._GEN_918                          (_GEN_1062),
  ._GEN_919                          (_GEN_1128),
  ._GEN_920                          (_GEN_1194),
  .rob_val_2_31                      (rob_val_2_31),
  .rob_val_2_30                      (rob_val_2_30),
  .rob_val_2_29                      (rob_val_2_29),
  .rob_val_2_28                      (rob_val_2_28),
  .rob_val_2_27                      (rob_val_2_27),
  .rob_val_2_26                      (rob_val_2_26),
  .rob_val_2_25                      (rob_val_2_25),
  .rob_val_2_24                      (rob_val_2_24),
  .rob_val_2_23                      (rob_val_2_23),
  .rob_val_2_22                      (rob_val_2_22),
  .rob_val_2_21                      (rob_val_2_21),
  .rob_val_2_20                      (rob_val_2_20),
  .rob_val_2_19                      (rob_val_2_19),
  .rob_val_2_18                      (rob_val_2_18),
  .rob_val_2_17                      (rob_val_2_17),
  .rob_val_2_16                      (rob_val_2_16),
  .rob_val_2_15                      (rob_val_2_15),
  .rob_val_2_14                      (rob_val_2_14),
  .rob_val_2_13                      (rob_val_2_13),
  .rob_val_2_12                      (rob_val_2_12),
  .rob_val_2_11                      (rob_val_2_11),
  .rob_val_2_10                      (rob_val_2_10),
  .rob_val_2_9                       (rob_val_2_9),
  .rob_val_2_8                       (rob_val_2_8),
  .rob_val_2_7                       (rob_val_2_7),
  .rob_val_2_6                       (rob_val_2_6),
  .rob_val_2_5                       (rob_val_2_5),
  .rob_val_2_4                       (rob_val_2_4),
  .rob_val_2_3                       (rob_val_2_3),
  .rob_val_2_2                       (rob_val_2_2),
  .rob_val_2_1                       (rob_val_2_1),
  .rob_val_2_0                       (rob_val_2_0),
  .io_enq_uops_2_rob_idx             (io_enq_uops_2_rob_idx),
  .rob_bsy_2_31                      (rob_bsy_2_31),
  .rob_bsy_2_30                      (rob_bsy_2_30),
  .rob_bsy_2_29                      (rob_bsy_2_29),
  .rob_bsy_2_28                      (rob_bsy_2_28),
  .rob_bsy_2_27                      (rob_bsy_2_27),
  .rob_bsy_2_26                      (rob_bsy_2_26),
  .rob_bsy_2_25                      (rob_bsy_2_25),
  .rob_bsy_2_24                      (rob_bsy_2_24),
  .rob_bsy_2_23                      (rob_bsy_2_23),
  .rob_bsy_2_22                      (rob_bsy_2_22),
  .rob_bsy_2_21                      (rob_bsy_2_21),
  .rob_bsy_2_20                      (rob_bsy_2_20),
  .rob_bsy_2_19                      (rob_bsy_2_19),
  .rob_bsy_2_18                      (rob_bsy_2_18),
  .rob_bsy_2_17                      (rob_bsy_2_17),
  .rob_bsy_2_16                      (rob_bsy_2_16),
  .rob_bsy_2_15                      (rob_bsy_2_15),
  .rob_bsy_2_14                      (rob_bsy_2_14),
  .rob_bsy_2_13                      (rob_bsy_2_13),
  .rob_bsy_2_12                      (rob_bsy_2_12),
  .rob_bsy_2_11                      (rob_bsy_2_11),
  .rob_bsy_2_10                      (rob_bsy_2_10),
  .rob_bsy_2_9                       (rob_bsy_2_9),
  .rob_bsy_2_8                       (rob_bsy_2_8),
  .rob_bsy_2_7                       (rob_bsy_2_7),
  .rob_bsy_2_6                       (rob_bsy_2_6),
  .rob_bsy_2_5                       (rob_bsy_2_5),
  .rob_bsy_2_4                       (rob_bsy_2_4),
  .rob_bsy_2_3                       (rob_bsy_2_3),
  .rob_bsy_2_2                       (rob_bsy_2_2),
  .rob_bsy_2_1                       (rob_bsy_2_1),
  .rob_bsy_2_0                       (rob_bsy_2_0),
  ._GEN_921                          (_GEN_1755),
  ._GEN_922                          (_GEN_1689),
  ._GEN_923                          (_GEN_1623),
  ._GEN_924                          (_GEN_1557),
  ._GEN_925                          (_GEN_1491),
  ._GEN_926                          (_GEN_1425),
  ._GEN_927                          (_GEN_1360),
  .io_enq_uops_2_uses_ldq            (io_enq_uops_2_uses_ldq),
  .io_enq_uops_2_is_br               (io_enq_uops_2_is_br),
  .io_enq_uops_2_is_jalr             (io_enq_uops_2_is_jalr),
  .io_enq_uops_2_uses_stq            (io_enq_uops_2_uses_stq),
  .io_enq_uops_2_is_fence            (io_enq_uops_2_is_fence),
  ._GEN_928                          (_GEN_1393),
  ._GEN_929                          (_GEN_1426),
  ._GEN_930                          (_GEN_1459),
  ._GEN_931                          (_GEN_1492),
  ._GEN_932                          (_GEN_1525),
  ._GEN_933                          (_GEN_1558),
  ._GEN_934                          (_GEN_1591),
  ._GEN_935                          (_GEN_1624),
  ._GEN_936                          (_GEN_1657),
  ._GEN_937                          (_GEN_1690),
  ._GEN_938                          (_GEN_1723),
  ._GEN_939                          (_GEN_1756),
  ._GEN_940                          (_GEN_1789),
  ._GEN_941                          (_GEN_1361),
  ._GEN_942                          (_GEN_1394),
  ._GEN_943                          (_GEN_1427),
  ._GEN_944                          (_GEN_1460),
  ._GEN_945                          (_GEN_1493),
  ._GEN_946                          (_GEN_1526),
  ._GEN_947                          (_GEN_1559),
  ._GEN_948                          (_GEN_1592),
  ._GEN_949                          (_GEN_1625),
  ._GEN_950                          (_GEN_1658),
  ._GEN_951                          (_GEN_1691),
  ._GEN_952                          (_GEN_1724),
  ._GEN_953                          (_GEN_1757),
  ._GEN_954                          (_GEN_1790),
  ._GEN_955                          (_GEN_1362),
  ._GEN_956                          (_GEN_1395),
  ._GEN_957                          (_GEN_1428),
  ._GEN_958                          (_GEN_1461),
  ._GEN_959                          (_GEN_1494),
  ._GEN_960                          (_GEN_1527),
  ._GEN_961                          (_GEN_1560),
  ._GEN_962                          (_GEN_1593),
  ._GEN_963                          (_GEN_1626),
  ._GEN_964                          (_GEN_1659),
  ._GEN_965                          (_GEN_1692),
  ._GEN_966                          (_GEN_1725),
  ._GEN_967                          (_GEN_1758),
  ._GEN_968                          (_GEN_1791),
  ._GEN_969                          (_GEN_1363),
  ._GEN_970                          (_GEN_1396),
  ._GEN_971                          (_GEN_1429),
  ._GEN_972                          (_GEN_1462),
  ._GEN_973                          (_GEN_1495),
  ._GEN_974                          (_GEN_1528),
  ._GEN_975                          (_GEN_1561),
  ._GEN_976                          (_GEN_1594),
  ._GEN_977                          (_GEN_1627),
  ._GEN_978                          (_GEN_1660),
  ._GEN_979                          (_GEN_1693),
  ._GEN_980                          (_GEN_1726),
  ._GEN_981                          (_GEN_1759),
  ._GEN_982                          (_GEN_1792),
  ._GEN_983                          (_GEN_1364),
  ._GEN_984                          (_GEN_1397),
  ._GEN_985                          (_GEN_1430),
  ._GEN_986                          (_GEN_1463),
  ._GEN_987                          (_GEN_1496),
  ._GEN_988                          (_GEN_1529),
  ._GEN_989                          (_GEN_1562),
  ._GEN_990                          (_GEN_1595),
  ._GEN_991                          (_GEN_1628),
  ._GEN_992                          (_GEN_1661),
  ._GEN_993                          (_GEN_1694),
  ._GEN_994                          (_GEN_1727),
  ._GEN_995                          (_GEN_1760),
  ._GEN_996                          (_GEN_1793),
  ._GEN_997                          (_GEN_1365),
  ._GEN_998                          (_GEN_1398),
  ._GEN_999                          (_GEN_1431),
  ._GEN_1000                         (_GEN_1464),
  ._GEN_1001                         (_GEN_1497),
  ._GEN_1002                         (_GEN_1530),
  ._GEN_1003                         (_GEN_1563),
  ._GEN_1004                         (_GEN_1596),
  ._GEN_1005                         (_GEN_1629),
  ._GEN_1006                         (_GEN_1662),
  ._GEN_1007                         (_GEN_1695),
  ._GEN_1008                         (_GEN_1728),
  ._GEN_1009                         (_GEN_1761),
  ._GEN_1010                         (_GEN_1794),
  ._GEN_1011                         (_GEN_1366),
  ._GEN_1012                         (_GEN_1399),
  ._GEN_1013                         (_GEN_1432),
  ._GEN_1014                         (_GEN_1465),
  ._GEN_1015                         (_GEN_1498),
  ._GEN_1016                         (_GEN_1531),
  ._GEN_1017                         (_GEN_1564),
  ._GEN_1018                         (_GEN_1597),
  ._GEN_1019                         (_GEN_1630),
  ._GEN_1020                         (_GEN_1663),
  ._GEN_1021                         (_GEN_1696),
  ._GEN_1022                         (_GEN_1729),
  ._GEN_1023                         (_GEN_1762),
  ._GEN_1024                         (_GEN_1795),
  ._GEN_1025                         (_GEN_1367),
  ._GEN_1026                         (_GEN_1400),
  ._GEN_1027                         (_GEN_1433),
  ._GEN_1028                         (_GEN_1466),
  ._GEN_1029                         (_GEN_1499),
  ._GEN_1030                         (_GEN_1532),
  ._GEN_1031                         (_GEN_1565),
  ._GEN_1032                         (_GEN_1598),
  ._GEN_1033                         (_GEN_1631),
  ._GEN_1034                         (_GEN_1664),
  ._GEN_1035                         (_GEN_1697),
  ._GEN_1036                         (_GEN_1730),
  ._GEN_1037                         (_GEN_1763),
  ._GEN_1038                         (_GEN_1796),
  ._GEN_1039                         (_GEN_1368),
  ._GEN_1040                         (_GEN_1401),
  ._GEN_1041                         (_GEN_1434),
  ._GEN_1042                         (_GEN_1467),
  ._GEN_1043                         (_GEN_1500),
  ._GEN_1044                         (_GEN_1533),
  ._GEN_1045                         (_GEN_1566),
  ._GEN_1046                         (_GEN_1599),
  ._GEN_1047                         (_GEN_1632),
  ._GEN_1048                         (_GEN_1665),
  ._GEN_1049                         (_GEN_1698),
  ._GEN_1050                         (_GEN_1731),
  ._GEN_1051                         (_GEN_1764),
  ._GEN_1052                         (_GEN_1797),
  ._GEN_1053                         (_GEN_1369),
  ._GEN_1054                         (_GEN_1402),
  ._GEN_1055                         (_GEN_1435),
  ._GEN_1056                         (_GEN_1468),
  ._GEN_1057                         (_GEN_1501),
  ._GEN_1058                         (_GEN_1534),
  ._GEN_1059                         (_GEN_1567),
  ._GEN_1060                         (_GEN_1600),
  ._GEN_1061                         (_GEN_1633),
  ._GEN_1062                         (_GEN_1666),
  ._GEN_1063                         (_GEN_1699),
  ._GEN_1064                         (_GEN_1732),
  ._GEN_1065                         (_GEN_1765),
  ._GEN_1066                         (_GEN_1798),
  ._GEN_1067                         (_GEN_1370),
  ._GEN_1068                         (_GEN_1403),
  ._GEN_1069                         (_GEN_1436),
  ._GEN_1070                         (_GEN_1469),
  ._GEN_1071                         (_GEN_1502),
  ._GEN_1072                         (_GEN_1535),
  ._GEN_1073                         (_GEN_1568),
  ._GEN_1074                         (_GEN_1601),
  ._GEN_1075                         (_GEN_1634),
  ._GEN_1076                         (_GEN_1667),
  ._GEN_1077                         (_GEN_1700),
  ._GEN_1078                         (_GEN_1733),
  ._GEN_1079                         (_GEN_1766),
  ._GEN_1080                         (_GEN_1799),
  ._GEN_1081                         (_GEN_1371),
  ._GEN_1082                         (_GEN_1404),
  ._GEN_1083                         (_GEN_1437),
  ._GEN_1084                         (_GEN_1470),
  ._GEN_1085                         (_GEN_1503),
  ._GEN_1086                         (_GEN_1536),
  ._GEN_1087                         (_GEN_1569),
  ._GEN_1088                         (_GEN_1602),
  ._GEN_1089                         (_GEN_1635),
  ._GEN_1090                         (_GEN_1668),
  ._GEN_1091                         (_GEN_1701),
  ._GEN_1092                         (_GEN_1734),
  ._GEN_1093                         (_GEN_1767),
  ._GEN_1094                         (_GEN_1800),
  ._GEN_1095                         (_GEN_1372),
  ._GEN_1096                         (_GEN_1405),
  ._GEN_1097                         (_GEN_1438),
  ._GEN_1098                         (_GEN_1471),
  ._GEN_1099                         (_GEN_1504),
  ._GEN_1100                         (_GEN_1537),
  ._GEN_1101                         (_GEN_1570),
  ._GEN_1102                         (_GEN_1603),
  ._GEN_1103                         (_GEN_1636),
  ._GEN_1104                         (_GEN_1669),
  ._GEN_1105                         (_GEN_1702),
  ._GEN_1106                         (_GEN_1735),
  ._GEN_1107                         (_GEN_1768),
  ._GEN_1108                         (_GEN_1801),
  ._GEN_1109                         (_GEN_1373),
  ._GEN_1110                         (_GEN_1406),
  ._GEN_1111                         (_GEN_1439),
  ._GEN_1112                         (_GEN_1472),
  ._GEN_1113                         (_GEN_1505),
  ._GEN_1114                         (_GEN_1538),
  ._GEN_1115                         (_GEN_1571),
  ._GEN_1116                         (_GEN_1604),
  ._GEN_1117                         (_GEN_1637),
  ._GEN_1118                         (_GEN_1670),
  ._GEN_1119                         (_GEN_1703),
  ._GEN_1120                         (_GEN_1736),
  ._GEN_1121                         (_GEN_1769),
  ._GEN_1122                         (_GEN_1802),
  ._GEN_1123                         (_GEN_1374),
  ._GEN_1124                         (_GEN_1407),
  ._GEN_1125                         (_GEN_1440),
  ._GEN_1126                         (_GEN_1473),
  ._GEN_1127                         (_GEN_1506),
  ._GEN_1128                         (_GEN_1539),
  ._GEN_1129                         (_GEN_1572),
  ._GEN_1130                         (_GEN_1605),
  ._GEN_1131                         (_GEN_1638),
  ._GEN_1132                         (_GEN_1671),
  ._GEN_1133                         (_GEN_1704),
  ._GEN_1134                         (_GEN_1737),
  ._GEN_1135                         (_GEN_1770),
  ._GEN_1136                         (_GEN_1803),
  ._GEN_1137                         (_GEN_1375),
  ._GEN_1138                         (_GEN_1408),
  ._GEN_1139                         (_GEN_1441),
  ._GEN_1140                         (_GEN_1474),
  ._GEN_1141                         (_GEN_1507),
  ._GEN_1142                         (_GEN_1540),
  ._GEN_1143                         (_GEN_1573),
  ._GEN_1144                         (_GEN_1606),
  ._GEN_1145                         (_GEN_1639),
  ._GEN_1146                         (_GEN_1672),
  ._GEN_1147                         (_GEN_1705),
  ._GEN_1148                         (_GEN_1738),
  ._GEN_1149                         (_GEN_1771),
  ._GEN_1150                         (_GEN_1804),
  ._GEN_1151                         (_GEN_1376),
  ._GEN_1152                         (_GEN_1409),
  ._GEN_1153                         (_GEN_1442),
  ._GEN_1154                         (_GEN_1475),
  ._GEN_1155                         (_GEN_1508),
  ._GEN_1156                         (_GEN_1541),
  ._GEN_1157                         (_GEN_1574),
  ._GEN_1158                         (_GEN_1607),
  ._GEN_1159                         (_GEN_1640),
  ._GEN_1160                         (_GEN_1673),
  ._GEN_1161                         (_GEN_1706),
  ._GEN_1162                         (_GEN_1739),
  ._GEN_1163                         (_GEN_1772),
  ._GEN_1164                         (_GEN_1805),
  ._GEN_1165                         (_GEN_1377),
  ._GEN_1166                         (_GEN_1410),
  ._GEN_1167                         (_GEN_1443),
  ._GEN_1168                         (_GEN_1476),
  ._GEN_1169                         (_GEN_1509),
  ._GEN_1170                         (_GEN_1542),
  ._GEN_1171                         (_GEN_1575),
  ._GEN_1172                         (_GEN_1608),
  ._GEN_1173                         (_GEN_1641),
  ._GEN_1174                         (_GEN_1674),
  ._GEN_1175                         (_GEN_1707),
  ._GEN_1176                         (_GEN_1740),
  ._GEN_1177                         (_GEN_1773),
  ._GEN_1178                         (_GEN_1806),
  ._GEN_1179                         (_GEN_1378),
  ._GEN_1180                         (_GEN_1411),
  ._GEN_1181                         (_GEN_1444),
  ._GEN_1182                         (_GEN_1477),
  ._GEN_1183                         (_GEN_1510),
  ._GEN_1184                         (_GEN_1543),
  ._GEN_1185                         (_GEN_1576),
  ._GEN_1186                         (_GEN_1609),
  ._GEN_1187                         (_GEN_1642),
  ._GEN_1188                         (_GEN_1675),
  ._GEN_1189                         (_GEN_1708),
  ._GEN_1190                         (_GEN_1741),
  ._GEN_1191                         (_GEN_1774),
  ._GEN_1192                         (_GEN_1807),
  ._GEN_1193                         (_GEN_1379),
  ._GEN_1194                         (_GEN_1412),
  ._GEN_1195                         (_GEN_1445),
  ._GEN_1196                         (_GEN_1478),
  ._GEN_1197                         (_GEN_1511),
  ._GEN_1198                         (_GEN_1544),
  ._GEN_1199                         (_GEN_1577),
  ._GEN_1200                         (_GEN_1610),
  ._GEN_1201                         (_GEN_1643),
  ._GEN_1202                         (_GEN_1676),
  ._GEN_1203                         (_GEN_1709),
  ._GEN_1204                         (_GEN_1742),
  ._GEN_1205                         (_GEN_1775),
  ._GEN_1206                         (_GEN_1808),
  ._GEN_1207                         (_GEN_1380),
  ._GEN_1208                         (_GEN_1413),
  ._GEN_1209                         (_GEN_1446),
  ._GEN_1210                         (_GEN_1479),
  ._GEN_1211                         (_GEN_1512),
  ._GEN_1212                         (_GEN_1545),
  ._GEN_1213                         (_GEN_1578),
  ._GEN_1214                         (_GEN_1611),
  ._GEN_1215                         (_GEN_1644),
  ._GEN_1216                         (_GEN_1677),
  ._GEN_1217                         (_GEN_1710),
  ._GEN_1218                         (_GEN_1743),
  ._GEN_1219                         (_GEN_1776),
  ._GEN_1220                         (_GEN_1809),
  ._GEN_1221                         (_GEN_1381),
  ._GEN_1222                         (_GEN_1414),
  ._GEN_1223                         (_GEN_1447),
  ._GEN_1224                         (_GEN_1480),
  ._GEN_1225                         (_GEN_1513),
  ._GEN_1226                         (_GEN_1546),
  ._GEN_1227                         (_GEN_1579),
  ._GEN_1228                         (_GEN_1612),
  ._GEN_1229                         (_GEN_1645),
  ._GEN_1230                         (_GEN_1678),
  ._GEN_1231                         (_GEN_1711),
  ._GEN_1232                         (_GEN_1744),
  ._GEN_1233                         (_GEN_1777),
  ._GEN_1234                         (_GEN_1810),
  ._GEN_1235                         (_GEN_1382),
  ._GEN_1236                         (_GEN_1415),
  ._GEN_1237                         (_GEN_1448),
  ._GEN_1238                         (_GEN_1481),
  ._GEN_1239                         (_GEN_1514),
  ._GEN_1240                         (_GEN_1547),
  ._GEN_1241                         (_GEN_1580),
  ._GEN_1242                         (_GEN_1613),
  ._GEN_1243                         (_GEN_1646),
  ._GEN_1244                         (_GEN_1679),
  ._GEN_1245                         (_GEN_1712),
  ._GEN_1246                         (_GEN_1745),
  ._GEN_1247                         (_GEN_1778),
  ._GEN_1248                         (_GEN_1811),
  ._GEN_1249                         (_GEN_1383),
  ._GEN_1250                         (_GEN_1416),
  ._GEN_1251                         (_GEN_1449),
  ._GEN_1252                         (_GEN_1482),
  ._GEN_1253                         (_GEN_1515),
  ._GEN_1254                         (_GEN_1548),
  ._GEN_1255                         (_GEN_1581),
  ._GEN_1256                         (_GEN_1614),
  ._GEN_1257                         (_GEN_1647),
  ._GEN_1258                         (_GEN_1680),
  ._GEN_1259                         (_GEN_1713),
  ._GEN_1260                         (_GEN_1746),
  ._GEN_1261                         (_GEN_1779),
  ._GEN_1262                         (_GEN_1812),
  ._GEN_1263                         (_GEN_1384),
  ._GEN_1264                         (_GEN_1417),
  ._GEN_1265                         (_GEN_1450),
  ._GEN_1266                         (_GEN_1483),
  ._GEN_1267                         (_GEN_1516),
  ._GEN_1268                         (_GEN_1549),
  ._GEN_1269                         (_GEN_1582),
  ._GEN_1270                         (_GEN_1615),
  ._GEN_1271                         (_GEN_1648),
  ._GEN_1272                         (_GEN_1681),
  ._GEN_1273                         (_GEN_1714),
  ._GEN_1274                         (_GEN_1747),
  ._GEN_1275                         (_GEN_1780),
  ._GEN_1276                         (_GEN_1813),
  ._GEN_1277                         (_GEN_1385),
  ._GEN_1278                         (_GEN_1418),
  ._GEN_1279                         (_GEN_1451),
  ._GEN_1280                         (_GEN_1484),
  ._GEN_1281                         (_GEN_1517),
  ._GEN_1282                         (_GEN_1550),
  ._GEN_1283                         (_GEN_1583),
  ._GEN_1284                         (_GEN_1616),
  ._GEN_1285                         (_GEN_1649),
  ._GEN_1286                         (_GEN_1682),
  ._GEN_1287                         (_GEN_1715),
  ._GEN_1288                         (_GEN_1748),
  ._GEN_1289                         (_GEN_1781),
  ._GEN_1290                         (_GEN_1814),
  ._GEN_1291                         (_GEN_1386),
  ._GEN_1292                         (_GEN_1419),
  ._GEN_1293                         (_GEN_1452),
  ._GEN_1294                         (_GEN_1485),
  ._GEN_1295                         (_GEN_1518),
  ._GEN_1296                         (_GEN_1551),
  ._GEN_1297                         (_GEN_1584),
  ._GEN_1298                         (_GEN_1617),
  ._GEN_1299                         (_GEN_1650),
  ._GEN_1300                         (_GEN_1683),
  ._GEN_1301                         (_GEN_1716),
  ._GEN_1302                         (_GEN_1749),
  ._GEN_1303                         (_GEN_1782),
  ._GEN_1304                         (_GEN_1815),
  ._GEN_1305                         (_GEN_1387),
  ._GEN_1306                         (_GEN_1420),
  ._GEN_1307                         (_GEN_1453),
  ._GEN_1308                         (_GEN_1486),
  ._GEN_1309                         (_GEN_1519),
  ._GEN_1310                         (_GEN_1552),
  ._GEN_1311                         (_GEN_1585),
  ._GEN_1312                         (_GEN_1618),
  ._GEN_1313                         (_GEN_1651),
  ._GEN_1314                         (_GEN_1684),
  ._GEN_1315                         (_GEN_1717),
  ._GEN_1316                         (_GEN_1750),
  ._GEN_1317                         (_GEN_1783),
  ._GEN_1318                         (_GEN_1816),
  ._GEN_1319                         (_GEN_1388),
  ._GEN_1320                         (_GEN_1421),
  ._GEN_1321                         (_GEN_1454),
  ._GEN_1322                         (_GEN_1487),
  ._GEN_1323                         (_GEN_1520),
  ._GEN_1324                         (_GEN_1553),
  ._GEN_1325                         (_GEN_1586),
  ._GEN_1326                         (_GEN_1619),
  ._GEN_1327                         (_GEN_1652),
  ._GEN_1328                         (_GEN_1685),
  ._GEN_1329                         (_GEN_1718),
  ._GEN_1330                         (_GEN_1751),
  ._GEN_1331                         (_GEN_1784),
  ._GEN_1332                         (_GEN_1817),
  ._GEN_1333                         (_GEN_1389),
  ._GEN_1334                         (_GEN_1422),
  ._GEN_1335                         (_GEN_1455),
  ._GEN_1336                         (_GEN_1488),
  ._GEN_1337                         (_GEN_1521),
  ._GEN_1338                         (_GEN_1554),
  ._GEN_1339                         (_GEN_1587),
  ._GEN_1340                         (_GEN_1620),
  ._GEN_1341                         (_GEN_1653),
  ._GEN_1342                         (_GEN_1686),
  ._GEN_1343                         (_GEN_1719),
  ._GEN_1344                         (_GEN_1752),
  ._GEN_1345                         (_GEN_1785),
  ._GEN_1346                         (_GEN_1818),
  ._GEN_1347                         (_GEN_1390),
  ._GEN_1348                         (_GEN_1423),
  ._GEN_1349                         (_GEN_1456),
  ._GEN_1350                         (_GEN_1489),
  ._GEN_1351                         (_GEN_1522),
  ._GEN_1352                         (_GEN_1555),
  ._GEN_1353                         (_GEN_1588),
  ._GEN_1354                         (_GEN_1621),
  ._GEN_1355                         (_GEN_1654),
  ._GEN_1356                         (_GEN_1687),
  ._GEN_1357                         (_GEN_1720),
  ._GEN_1358                         (_GEN_1753),
  ._GEN_1359                         (_GEN_1786),
  ._GEN_1360                         (_GEN_1819),
  ._GEN_1361                         (_GEN_1391),
  ._GEN_1362                         (_GEN_1424),
  ._GEN_1363                         (_GEN_1457),
  ._GEN_1364                         (_GEN_1490),
  ._GEN_1365                         (_GEN_1523),
  ._GEN_1366                         (_GEN_1556),
  ._GEN_1367                         (_GEN_1589),
  ._GEN_1368                         (_GEN_1622),
  ._GEN_1369                         (_GEN_1655),
  ._GEN_1370                         (_GEN_1688),
  ._GEN_1371                         (_GEN_1721),
  ._GEN_1372                         (_GEN_1754),
  ._GEN_1373                         (_GEN_1787),
  ._GEN_1374                         (_GEN_1820),
  ._GEN_1375                         (_GEN_1392),
  .rob_uop_2_31_pdst                 (rob_uop_2_31_pdst),
  .rob_uop_2_30_pdst                 (rob_uop_2_30_pdst),
  .rob_uop_2_29_pdst                 (rob_uop_2_29_pdst),
  .rob_uop_2_28_pdst                 (rob_uop_2_28_pdst),
  .rob_uop_2_27_pdst                 (rob_uop_2_27_pdst),
  .rob_uop_2_26_pdst                 (rob_uop_2_26_pdst),
  .rob_uop_2_25_pdst                 (rob_uop_2_25_pdst),
  .rob_uop_2_24_pdst                 (rob_uop_2_24_pdst),
  .rob_uop_2_23_pdst                 (rob_uop_2_23_pdst),
  .rob_uop_2_22_pdst                 (rob_uop_2_22_pdst),
  .rob_uop_2_21_pdst                 (rob_uop_2_21_pdst),
  .rob_uop_2_20_pdst                 (rob_uop_2_20_pdst),
  .rob_uop_2_19_pdst                 (rob_uop_2_19_pdst),
  .rob_uop_2_18_pdst                 (rob_uop_2_18_pdst),
  .rob_uop_2_17_pdst                 (rob_uop_2_17_pdst),
  .rob_uop_2_16_pdst                 (rob_uop_2_16_pdst),
  .rob_uop_2_15_pdst                 (rob_uop_2_15_pdst),
  .rob_uop_2_14_pdst                 (rob_uop_2_14_pdst),
  .rob_uop_2_13_pdst                 (rob_uop_2_13_pdst),
  .rob_uop_2_12_pdst                 (rob_uop_2_12_pdst),
  .rob_uop_2_11_pdst                 (rob_uop_2_11_pdst),
  .rob_uop_2_10_pdst                 (rob_uop_2_10_pdst),
  .rob_uop_2_9_pdst                  (rob_uop_2_9_pdst),
  .rob_uop_2_8_pdst                  (rob_uop_2_8_pdst),
  .rob_uop_2_7_pdst                  (rob_uop_2_7_pdst),
  .rob_uop_2_6_pdst                  (rob_uop_2_6_pdst),
  .rob_uop_2_5_pdst                  (rob_uop_2_5_pdst),
  .rob_uop_2_4_pdst                  (rob_uop_2_4_pdst),
  .rob_uop_2_3_pdst                  (rob_uop_2_3_pdst),
  .rob_uop_2_2_pdst                  (rob_uop_2_2_pdst),
  .rob_uop_2_1_pdst                  (rob_uop_2_1_pdst),
  .rob_uop_2_0_pdst                  (rob_uop_2_0_pdst),
  .rob_uop_2_31_ldst_val             (rob_uop_2_31_ldst_val),
  .rob_uop_2_30_ldst_val             (rob_uop_2_30_ldst_val),
  .rob_uop_2_29_ldst_val             (rob_uop_2_29_ldst_val),
  .rob_uop_2_28_ldst_val             (rob_uop_2_28_ldst_val),
  .rob_uop_2_27_ldst_val             (rob_uop_2_27_ldst_val),
  .rob_uop_2_26_ldst_val             (rob_uop_2_26_ldst_val),
  .rob_uop_2_25_ldst_val             (rob_uop_2_25_ldst_val),
  .rob_uop_2_24_ldst_val             (rob_uop_2_24_ldst_val),
  .rob_uop_2_23_ldst_val             (rob_uop_2_23_ldst_val),
  .rob_uop_2_22_ldst_val             (rob_uop_2_22_ldst_val),
  .rob_uop_2_21_ldst_val             (rob_uop_2_21_ldst_val),
  .rob_uop_2_20_ldst_val             (rob_uop_2_20_ldst_val),
  .rob_uop_2_19_ldst_val             (rob_uop_2_19_ldst_val),
  .rob_uop_2_18_ldst_val             (rob_uop_2_18_ldst_val),
  .rob_uop_2_17_ldst_val             (rob_uop_2_17_ldst_val),
  .rob_uop_2_16_ldst_val             (rob_uop_2_16_ldst_val),
  .rob_uop_2_15_ldst_val             (rob_uop_2_15_ldst_val),
  .rob_uop_2_14_ldst_val             (rob_uop_2_14_ldst_val),
  .rob_uop_2_13_ldst_val             (rob_uop_2_13_ldst_val),
  .rob_uop_2_12_ldst_val             (rob_uop_2_12_ldst_val),
  .rob_uop_2_11_ldst_val             (rob_uop_2_11_ldst_val),
  .rob_uop_2_10_ldst_val             (rob_uop_2_10_ldst_val),
  .rob_uop_2_9_ldst_val              (rob_uop_2_9_ldst_val),
  .rob_uop_2_8_ldst_val              (rob_uop_2_8_ldst_val),
  .rob_uop_2_7_ldst_val              (rob_uop_2_7_ldst_val),
  .rob_uop_2_6_ldst_val              (rob_uop_2_6_ldst_val),
  .rob_uop_2_5_ldst_val              (rob_uop_2_5_ldst_val),
  .rob_uop_2_4_ldst_val              (rob_uop_2_4_ldst_val),
  .rob_uop_2_3_ldst_val              (rob_uop_2_3_ldst_val),
  .rob_uop_2_2_ldst_val              (rob_uop_2_2_ldst_val),
  .rob_uop_2_1_ldst_val              (rob_uop_2_1_ldst_val),
  .rob_uop_2_0_ldst_val              (rob_uop_2_0_ldst_val),
  ._GEN_1376                         (_GEN_1458),
  ._GEN_1377                         (_GEN_1524),
  ._GEN_1378                         (_GEN_1590),
  ._GEN_1379                         (_GEN_1656),
  .rob_val_3_31                      (rob_val_3_31),
  .rob_val_3_30                      (rob_val_3_30),
  .rob_val_3_29                      (rob_val_3_29),
  .rob_val_3_28                      (rob_val_3_28),
  .rob_val_3_27                      (rob_val_3_27),
  .rob_val_3_26                      (rob_val_3_26),
  .rob_val_3_25                      (rob_val_3_25),
  .rob_val_3_24                      (rob_val_3_24),
  .rob_val_3_23                      (rob_val_3_23),
  .rob_val_3_22                      (rob_val_3_22),
  .rob_val_3_21                      (rob_val_3_21),
  .rob_val_3_20                      (rob_val_3_20),
  .rob_val_3_19                      (rob_val_3_19),
  .rob_val_3_18                      (rob_val_3_18),
  .rob_val_3_17                      (rob_val_3_17),
  .rob_val_3_16                      (rob_val_3_16),
  .rob_val_3_15                      (rob_val_3_15),
  .rob_val_3_14                      (rob_val_3_14),
  .rob_val_3_13                      (rob_val_3_13),
  .rob_val_3_12                      (rob_val_3_12),
  .rob_val_3_11                      (rob_val_3_11),
  .rob_val_3_10                      (rob_val_3_10),
  .rob_val_3_9                       (rob_val_3_9),
  .rob_val_3_8                       (rob_val_3_8),
  .rob_val_3_7                       (rob_val_3_7),
  .rob_val_3_6                       (rob_val_3_6),
  .rob_val_3_5                       (rob_val_3_5),
  .rob_val_3_4                       (rob_val_3_4),
  .rob_val_3_3                       (rob_val_3_3),
  .rob_val_3_2                       (rob_val_3_2),
  .rob_val_3_1                       (rob_val_3_1),
  .rob_val_3_0                       (rob_val_3_0),
  .io_enq_uops_3_rob_idx             (io_enq_uops_3_rob_idx),
  .rob_bsy_3_31                      (rob_bsy_3_31),
  .rob_bsy_3_30                      (rob_bsy_3_30),
  .rob_bsy_3_29                      (rob_bsy_3_29),
  .rob_bsy_3_28                      (rob_bsy_3_28),
  .rob_bsy_3_27                      (rob_bsy_3_27),
  .rob_bsy_3_26                      (rob_bsy_3_26),
  .rob_bsy_3_25                      (rob_bsy_3_25),
  .rob_bsy_3_24                      (rob_bsy_3_24),
  .rob_bsy_3_23                      (rob_bsy_3_23),
  .rob_bsy_3_22                      (rob_bsy_3_22),
  .rob_bsy_3_21                      (rob_bsy_3_21),
  .rob_bsy_3_20                      (rob_bsy_3_20),
  .rob_bsy_3_19                      (rob_bsy_3_19),
  .rob_bsy_3_18                      (rob_bsy_3_18),
  .rob_bsy_3_17                      (rob_bsy_3_17),
  .rob_bsy_3_16                      (rob_bsy_3_16),
  .rob_bsy_3_15                      (rob_bsy_3_15),
  .rob_bsy_3_14                      (rob_bsy_3_14),
  .rob_bsy_3_13                      (rob_bsy_3_13),
  .rob_bsy_3_12                      (rob_bsy_3_12),
  .rob_bsy_3_11                      (rob_bsy_3_11),
  .rob_bsy_3_10                      (rob_bsy_3_10),
  .rob_bsy_3_9                       (rob_bsy_3_9),
  .rob_bsy_3_8                       (rob_bsy_3_8),
  .rob_bsy_3_7                       (rob_bsy_3_7),
  .rob_bsy_3_6                       (rob_bsy_3_6),
  .rob_bsy_3_5                       (rob_bsy_3_5),
  .rob_bsy_3_4                       (rob_bsy_3_4),
  .rob_bsy_3_3                       (rob_bsy_3_3),
  .rob_bsy_3_2                       (rob_bsy_3_2),
  .rob_bsy_3_1                       (rob_bsy_3_1),
  .rob_bsy_3_0                       (rob_bsy_3_0),
  ._GEN_1380                         (_GEN_2217),
  ._GEN_1381                         (_GEN_2151),
  ._GEN_1382                         (_GEN_2085),
  ._GEN_1383                         (_GEN_2019),
  ._GEN_1384                         (_GEN_1953),
  ._GEN_1385                         (_GEN_1887),
  ._GEN_1386                         (_GEN_1822),
  .io_enq_uops_3_uses_ldq            (io_enq_uops_3_uses_ldq),
  .io_enq_uops_3_is_br               (io_enq_uops_3_is_br),
  .io_enq_uops_3_is_jalr             (io_enq_uops_3_is_jalr),
  .io_enq_uops_3_uses_stq            (io_enq_uops_3_uses_stq),
  .io_enq_uops_3_is_fence            (io_enq_uops_3_is_fence),
  ._GEN_1387                         (_GEN_1855),
  ._GEN_1388                         (_GEN_1888),
  ._GEN_1389                         (_GEN_1921),
  ._GEN_1390                         (_GEN_1954),
  ._GEN_1391                         (_GEN_1987),
  ._GEN_1392                         (_GEN_2020),
  ._GEN_1393                         (_GEN_2053),
  ._GEN_1394                         (_GEN_2086),
  ._GEN_1395                         (_GEN_2119),
  ._GEN_1396                         (_GEN_2152),
  ._GEN_1397                         (_GEN_2185),
  ._GEN_1398                         (_GEN_2218),
  ._GEN_1399                         (_GEN_2251),
  ._GEN_1400                         (_GEN_1823),
  ._GEN_1401                         (_GEN_1856),
  ._GEN_1402                         (_GEN_1889),
  ._GEN_1403                         (_GEN_1922),
  ._GEN_1404                         (_GEN_1955),
  ._GEN_1405                         (_GEN_1988),
  ._GEN_1406                         (_GEN_2021),
  ._GEN_1407                         (_GEN_2054),
  ._GEN_1408                         (_GEN_2087),
  ._GEN_1409                         (_GEN_2120),
  ._GEN_1410                         (_GEN_2153),
  ._GEN_1411                         (_GEN_2186),
  ._GEN_1412                         (_GEN_2219),
  ._GEN_1413                         (_GEN_2252),
  ._GEN_1414                         (_GEN_1824),
  ._GEN_1415                         (_GEN_1857),
  ._GEN_1416                         (_GEN_1890),
  ._GEN_1417                         (_GEN_1923),
  ._GEN_1418                         (_GEN_1956),
  ._GEN_1419                         (_GEN_1989),
  ._GEN_1420                         (_GEN_2022),
  ._GEN_1421                         (_GEN_2055),
  ._GEN_1422                         (_GEN_2088),
  ._GEN_1423                         (_GEN_2121),
  ._GEN_1424                         (_GEN_2154),
  ._GEN_1425                         (_GEN_2187),
  ._GEN_1426                         (_GEN_2220),
  ._GEN_1427                         (_GEN_2253),
  ._GEN_1428                         (_GEN_1825),
  ._GEN_1429                         (_GEN_1858),
  ._GEN_1430                         (_GEN_1891),
  ._GEN_1431                         (_GEN_1924),
  ._GEN_1432                         (_GEN_1957),
  ._GEN_1433                         (_GEN_1990),
  ._GEN_1434                         (_GEN_2023),
  ._GEN_1435                         (_GEN_2056),
  ._GEN_1436                         (_GEN_2089),
  ._GEN_1437                         (_GEN_2122),
  ._GEN_1438                         (_GEN_2155),
  ._GEN_1439                         (_GEN_2188),
  ._GEN_1440                         (_GEN_2221),
  ._GEN_1441                         (_GEN_2254),
  ._GEN_1442                         (_GEN_1826),
  ._GEN_1443                         (_GEN_1859),
  ._GEN_1444                         (_GEN_1892),
  ._GEN_1445                         (_GEN_1925),
  ._GEN_1446                         (_GEN_1958),
  ._GEN_1447                         (_GEN_1991),
  ._GEN_1448                         (_GEN_2024),
  ._GEN_1449                         (_GEN_2057),
  ._GEN_1450                         (_GEN_2090),
  ._GEN_1451                         (_GEN_2123),
  ._GEN_1452                         (_GEN_2156),
  ._GEN_1453                         (_GEN_2189),
  ._GEN_1454                         (_GEN_2222),
  ._GEN_1455                         (_GEN_2255),
  ._GEN_1456                         (_GEN_1827),
  ._GEN_1457                         (_GEN_1860),
  ._GEN_1458                         (_GEN_1893),
  ._GEN_1459                         (_GEN_1926),
  ._GEN_1460                         (_GEN_1959),
  ._GEN_1461                         (_GEN_1992),
  ._GEN_1462                         (_GEN_2025),
  ._GEN_1463                         (_GEN_2058),
  ._GEN_1464                         (_GEN_2091),
  ._GEN_1465                         (_GEN_2124),
  ._GEN_1466                         (_GEN_2157),
  ._GEN_1467                         (_GEN_2190),
  ._GEN_1468                         (_GEN_2223),
  ._GEN_1469                         (_GEN_2256),
  ._GEN_1470                         (_GEN_1828),
  ._GEN_1471                         (_GEN_1861),
  ._GEN_1472                         (_GEN_1894),
  ._GEN_1473                         (_GEN_1927),
  ._GEN_1474                         (_GEN_1960),
  ._GEN_1475                         (_GEN_1993),
  ._GEN_1476                         (_GEN_2026),
  ._GEN_1477                         (_GEN_2059),
  ._GEN_1478                         (_GEN_2092),
  ._GEN_1479                         (_GEN_2125),
  ._GEN_1480                         (_GEN_2158),
  ._GEN_1481                         (_GEN_2191),
  ._GEN_1482                         (_GEN_2224),
  ._GEN_1483                         (_GEN_2257),
  ._GEN_1484                         (_GEN_1829),
  ._GEN_1485                         (_GEN_1862),
  ._GEN_1486                         (_GEN_1895),
  ._GEN_1487                         (_GEN_1928),
  ._GEN_1488                         (_GEN_1961),
  ._GEN_1489                         (_GEN_1994),
  ._GEN_1490                         (_GEN_2027),
  ._GEN_1491                         (_GEN_2060),
  ._GEN_1492                         (_GEN_2093),
  ._GEN_1493                         (_GEN_2126),
  ._GEN_1494                         (_GEN_2159),
  ._GEN_1495                         (_GEN_2192),
  ._GEN_1496                         (_GEN_2225),
  ._GEN_1497                         (_GEN_2258),
  ._GEN_1498                         (_GEN_1830),
  ._GEN_1499                         (_GEN_1863),
  ._GEN_1500                         (_GEN_1896),
  ._GEN_1501                         (_GEN_1929),
  ._GEN_1502                         (_GEN_1962),
  ._GEN_1503                         (_GEN_1995),
  ._GEN_1504                         (_GEN_2028),
  ._GEN_1505                         (_GEN_2061),
  ._GEN_1506                         (_GEN_2094),
  ._GEN_1507                         (_GEN_2127),
  ._GEN_1508                         (_GEN_2160),
  ._GEN_1509                         (_GEN_2193),
  ._GEN_1510                         (_GEN_2226),
  ._GEN_1511                         (_GEN_2259),
  ._GEN_1512                         (_GEN_1831),
  ._GEN_1513                         (_GEN_1864),
  ._GEN_1514                         (_GEN_1897),
  ._GEN_1515                         (_GEN_1930),
  ._GEN_1516                         (_GEN_1963),
  ._GEN_1517                         (_GEN_1996),
  ._GEN_1518                         (_GEN_2029),
  ._GEN_1519                         (_GEN_2062),
  ._GEN_1520                         (_GEN_2095),
  ._GEN_1521                         (_GEN_2128),
  ._GEN_1522                         (_GEN_2161),
  ._GEN_1523                         (_GEN_2194),
  ._GEN_1524                         (_GEN_2227),
  ._GEN_1525                         (_GEN_2260),
  ._GEN_1526                         (_GEN_1832),
  ._GEN_1527                         (_GEN_1865),
  ._GEN_1528                         (_GEN_1898),
  ._GEN_1529                         (_GEN_1931),
  ._GEN_1530                         (_GEN_1964),
  ._GEN_1531                         (_GEN_1997),
  ._GEN_1532                         (_GEN_2030),
  ._GEN_1533                         (_GEN_2063),
  ._GEN_1534                         (_GEN_2096),
  ._GEN_1535                         (_GEN_2129),
  ._GEN_1536                         (_GEN_2162),
  ._GEN_1537                         (_GEN_2195),
  ._GEN_1538                         (_GEN_2228),
  ._GEN_1539                         (_GEN_2261),
  ._GEN_1540                         (_GEN_1833),
  ._GEN_1541                         (_GEN_1866),
  ._GEN_1542                         (_GEN_1899),
  ._GEN_1543                         (_GEN_1932),
  ._GEN_1544                         (_GEN_1965),
  ._GEN_1545                         (_GEN_1998),
  ._GEN_1546                         (_GEN_2031),
  ._GEN_1547                         (_GEN_2064),
  ._GEN_1548                         (_GEN_2097),
  ._GEN_1549                         (_GEN_2130),
  ._GEN_1550                         (_GEN_2163),
  ._GEN_1551                         (_GEN_2196),
  ._GEN_1552                         (_GEN_2229),
  ._GEN_1553                         (_GEN_2262),
  ._GEN_1554                         (_GEN_1834),
  ._GEN_1555                         (_GEN_1867),
  ._GEN_1556                         (_GEN_1900),
  ._GEN_1557                         (_GEN_1933),
  ._GEN_1558                         (_GEN_1966),
  ._GEN_1559                         (_GEN_1999),
  ._GEN_1560                         (_GEN_2032),
  ._GEN_1561                         (_GEN_2065),
  ._GEN_1562                         (_GEN_2098),
  ._GEN_1563                         (_GEN_2131),
  ._GEN_1564                         (_GEN_2164),
  ._GEN_1565                         (_GEN_2197),
  ._GEN_1566                         (_GEN_2230),
  ._GEN_1567                         (_GEN_2263),
  ._GEN_1568                         (_GEN_1835),
  ._GEN_1569                         (_GEN_1868),
  ._GEN_1570                         (_GEN_1901),
  ._GEN_1571                         (_GEN_1934),
  ._GEN_1572                         (_GEN_1967),
  ._GEN_1573                         (_GEN_2000),
  ._GEN_1574                         (_GEN_2033),
  ._GEN_1575                         (_GEN_2066),
  ._GEN_1576                         (_GEN_2099),
  ._GEN_1577                         (_GEN_2132),
  ._GEN_1578                         (_GEN_2165),
  ._GEN_1579                         (_GEN_2198),
  ._GEN_1580                         (_GEN_2231),
  ._GEN_1581                         (_GEN_2264),
  ._GEN_1582                         (_GEN_1836),
  ._GEN_1583                         (_GEN_1869),
  ._GEN_1584                         (_GEN_1902),
  ._GEN_1585                         (_GEN_1935),
  ._GEN_1586                         (_GEN_1968),
  ._GEN_1587                         (_GEN_2001),
  ._GEN_1588                         (_GEN_2034),
  ._GEN_1589                         (_GEN_2067),
  ._GEN_1590                         (_GEN_2100),
  ._GEN_1591                         (_GEN_2133),
  ._GEN_1592                         (_GEN_2166),
  ._GEN_1593                         (_GEN_2199),
  ._GEN_1594                         (_GEN_2232),
  ._GEN_1595                         (_GEN_2265),
  ._GEN_1596                         (_GEN_1837),
  ._GEN_1597                         (_GEN_1870),
  ._GEN_1598                         (_GEN_1903),
  ._GEN_1599                         (_GEN_1936),
  ._GEN_1600                         (_GEN_1969),
  ._GEN_1601                         (_GEN_2002),
  ._GEN_1602                         (_GEN_2035),
  ._GEN_1603                         (_GEN_2068),
  ._GEN_1604                         (_GEN_2101),
  ._GEN_1605                         (_GEN_2134),
  ._GEN_1606                         (_GEN_2167),
  ._GEN_1607                         (_GEN_2200),
  ._GEN_1608                         (_GEN_2233),
  ._GEN_1609                         (_GEN_2266),
  ._GEN_1610                         (_GEN_1838),
  ._GEN_1611                         (_GEN_1871),
  ._GEN_1612                         (_GEN_1904),
  ._GEN_1613                         (_GEN_1937),
  ._GEN_1614                         (_GEN_1970),
  ._GEN_1615                         (_GEN_2003),
  ._GEN_1616                         (_GEN_2036),
  ._GEN_1617                         (_GEN_2069),
  ._GEN_1618                         (_GEN_2102),
  ._GEN_1619                         (_GEN_2135),
  ._GEN_1620                         (_GEN_2168),
  ._GEN_1621                         (_GEN_2201),
  ._GEN_1622                         (_GEN_2234),
  ._GEN_1623                         (_GEN_2267),
  ._GEN_1624                         (_GEN_1839),
  ._GEN_1625                         (_GEN_1872),
  ._GEN_1626                         (_GEN_1905),
  ._GEN_1627                         (_GEN_1938),
  ._GEN_1628                         (_GEN_1971),
  ._GEN_1629                         (_GEN_2004),
  ._GEN_1630                         (_GEN_2037),
  ._GEN_1631                         (_GEN_2070),
  ._GEN_1632                         (_GEN_2103),
  ._GEN_1633                         (_GEN_2136),
  ._GEN_1634                         (_GEN_2169),
  ._GEN_1635                         (_GEN_2202),
  ._GEN_1636                         (_GEN_2235),
  ._GEN_1637                         (_GEN_2268),
  ._GEN_1638                         (_GEN_1840),
  ._GEN_1639                         (_GEN_1873),
  ._GEN_1640                         (_GEN_1906),
  ._GEN_1641                         (_GEN_1939),
  ._GEN_1642                         (_GEN_1972),
  ._GEN_1643                         (_GEN_2005),
  ._GEN_1644                         (_GEN_2038),
  ._GEN_1645                         (_GEN_2071),
  ._GEN_1646                         (_GEN_2104),
  ._GEN_1647                         (_GEN_2137),
  ._GEN_1648                         (_GEN_2170),
  ._GEN_1649                         (_GEN_2203),
  ._GEN_1650                         (_GEN_2236),
  ._GEN_1651                         (_GEN_2269),
  ._GEN_1652                         (_GEN_1841),
  ._GEN_1653                         (_GEN_1874),
  ._GEN_1654                         (_GEN_1907),
  ._GEN_1655                         (_GEN_1940),
  ._GEN_1656                         (_GEN_1973),
  ._GEN_1657                         (_GEN_2006),
  ._GEN_1658                         (_GEN_2039),
  ._GEN_1659                         (_GEN_2072),
  ._GEN_1660                         (_GEN_2105),
  ._GEN_1661                         (_GEN_2138),
  ._GEN_1662                         (_GEN_2171),
  ._GEN_1663                         (_GEN_2204),
  ._GEN_1664                         (_GEN_2237),
  ._GEN_1665                         (_GEN_2270),
  ._GEN_1666                         (_GEN_1842),
  ._GEN_1667                         (_GEN_1875),
  ._GEN_1668                         (_GEN_1908),
  ._GEN_1669                         (_GEN_1941),
  ._GEN_1670                         (_GEN_1974),
  ._GEN_1671                         (_GEN_2007),
  ._GEN_1672                         (_GEN_2040),
  ._GEN_1673                         (_GEN_2073),
  ._GEN_1674                         (_GEN_2106),
  ._GEN_1675                         (_GEN_2139),
  ._GEN_1676                         (_GEN_2172),
  ._GEN_1677                         (_GEN_2205),
  ._GEN_1678                         (_GEN_2238),
  ._GEN_1679                         (_GEN_2271),
  ._GEN_1680                         (_GEN_1843),
  ._GEN_1681                         (_GEN_1876),
  ._GEN_1682                         (_GEN_1909),
  ._GEN_1683                         (_GEN_1942),
  ._GEN_1684                         (_GEN_1975),
  ._GEN_1685                         (_GEN_2008),
  ._GEN_1686                         (_GEN_2041),
  ._GEN_1687                         (_GEN_2074),
  ._GEN_1688                         (_GEN_2107),
  ._GEN_1689                         (_GEN_2140),
  ._GEN_1690                         (_GEN_2173),
  ._GEN_1691                         (_GEN_2206),
  ._GEN_1692                         (_GEN_2239),
  ._GEN_1693                         (_GEN_2272),
  ._GEN_1694                         (_GEN_1844),
  ._GEN_1695                         (_GEN_1877),
  ._GEN_1696                         (_GEN_1910),
  ._GEN_1697                         (_GEN_1943),
  ._GEN_1698                         (_GEN_1976),
  ._GEN_1699                         (_GEN_2009),
  ._GEN_1700                         (_GEN_2042),
  ._GEN_1701                         (_GEN_2075),
  ._GEN_1702                         (_GEN_2108),
  ._GEN_1703                         (_GEN_2141),
  ._GEN_1704                         (_GEN_2174),
  ._GEN_1705                         (_GEN_2207),
  ._GEN_1706                         (_GEN_2240),
  ._GEN_1707                         (_GEN_2273),
  ._GEN_1708                         (_GEN_1845),
  ._GEN_1709                         (_GEN_1878),
  ._GEN_1710                         (_GEN_1911),
  ._GEN_1711                         (_GEN_1944),
  ._GEN_1712                         (_GEN_1977),
  ._GEN_1713                         (_GEN_2010),
  ._GEN_1714                         (_GEN_2043),
  ._GEN_1715                         (_GEN_2076),
  ._GEN_1716                         (_GEN_2109),
  ._GEN_1717                         (_GEN_2142),
  ._GEN_1718                         (_GEN_2175),
  ._GEN_1719                         (_GEN_2208),
  ._GEN_1720                         (_GEN_2241),
  ._GEN_1721                         (_GEN_2274),
  ._GEN_1722                         (_GEN_1846),
  ._GEN_1723                         (_GEN_1879),
  ._GEN_1724                         (_GEN_1912),
  ._GEN_1725                         (_GEN_1945),
  ._GEN_1726                         (_GEN_1978),
  ._GEN_1727                         (_GEN_2011),
  ._GEN_1728                         (_GEN_2044),
  ._GEN_1729                         (_GEN_2077),
  ._GEN_1730                         (_GEN_2110),
  ._GEN_1731                         (_GEN_2143),
  ._GEN_1732                         (_GEN_2176),
  ._GEN_1733                         (_GEN_2209),
  ._GEN_1734                         (_GEN_2242),
  ._GEN_1735                         (_GEN_2275),
  ._GEN_1736                         (_GEN_1847),
  ._GEN_1737                         (_GEN_1880),
  ._GEN_1738                         (_GEN_1913),
  ._GEN_1739                         (_GEN_1946),
  ._GEN_1740                         (_GEN_1979),
  ._GEN_1741                         (_GEN_2012),
  ._GEN_1742                         (_GEN_2045),
  ._GEN_1743                         (_GEN_2078),
  ._GEN_1744                         (_GEN_2111),
  ._GEN_1745                         (_GEN_2144),
  ._GEN_1746                         (_GEN_2177),
  ._GEN_1747                         (_GEN_2210),
  ._GEN_1748                         (_GEN_2243),
  ._GEN_1749                         (_GEN_2276),
  ._GEN_1750                         (_GEN_1848),
  ._GEN_1751                         (_GEN_1881),
  ._GEN_1752                         (_GEN_1914),
  ._GEN_1753                         (_GEN_1947),
  ._GEN_1754                         (_GEN_1980),
  ._GEN_1755                         (_GEN_2013),
  ._GEN_1756                         (_GEN_2046),
  ._GEN_1757                         (_GEN_2079),
  ._GEN_1758                         (_GEN_2112),
  ._GEN_1759                         (_GEN_2145),
  ._GEN_1760                         (_GEN_2178),
  ._GEN_1761                         (_GEN_2211),
  ._GEN_1762                         (_GEN_2244),
  ._GEN_1763                         (_GEN_2277),
  ._GEN_1764                         (_GEN_1849),
  ._GEN_1765                         (_GEN_1882),
  ._GEN_1766                         (_GEN_1915),
  ._GEN_1767                         (_GEN_1948),
  ._GEN_1768                         (_GEN_1981),
  ._GEN_1769                         (_GEN_2014),
  ._GEN_1770                         (_GEN_2047),
  ._GEN_1771                         (_GEN_2080),
  ._GEN_1772                         (_GEN_2113),
  ._GEN_1773                         (_GEN_2146),
  ._GEN_1774                         (_GEN_2179),
  ._GEN_1775                         (_GEN_2212),
  ._GEN_1776                         (_GEN_2245),
  ._GEN_1777                         (_GEN_2278),
  ._GEN_1778                         (_GEN_1850),
  ._GEN_1779                         (_GEN_1883),
  ._GEN_1780                         (_GEN_1916),
  ._GEN_1781                         (_GEN_1949),
  ._GEN_1782                         (_GEN_1982),
  ._GEN_1783                         (_GEN_2015),
  ._GEN_1784                         (_GEN_2048),
  ._GEN_1785                         (_GEN_2081),
  ._GEN_1786                         (_GEN_2114),
  ._GEN_1787                         (_GEN_2147),
  ._GEN_1788                         (_GEN_2180),
  ._GEN_1789                         (_GEN_2213),
  ._GEN_1790                         (_GEN_2246),
  ._GEN_1791                         (_GEN_2279),
  ._GEN_1792                         (_GEN_1851),
  ._GEN_1793                         (_GEN_1884),
  ._GEN_1794                         (_GEN_1917),
  ._GEN_1795                         (_GEN_1950),
  ._GEN_1796                         (_GEN_1983),
  ._GEN_1797                         (_GEN_2016),
  ._GEN_1798                         (_GEN_2049),
  ._GEN_1799                         (_GEN_2082),
  ._GEN_1800                         (_GEN_2115),
  ._GEN_1801                         (_GEN_2148),
  ._GEN_1802                         (_GEN_2181),
  ._GEN_1803                         (_GEN_2214),
  ._GEN_1804                         (_GEN_2247),
  ._GEN_1805                         (_GEN_2280),
  ._GEN_1806                         (_GEN_1852),
  ._GEN_1807                         (_GEN_1885),
  ._GEN_1808                         (_GEN_1918),
  ._GEN_1809                         (_GEN_1951),
  ._GEN_1810                         (_GEN_1984),
  ._GEN_1811                         (_GEN_2017),
  ._GEN_1812                         (_GEN_2050),
  ._GEN_1813                         (_GEN_2083),
  ._GEN_1814                         (_GEN_2116),
  ._GEN_1815                         (_GEN_2149),
  ._GEN_1816                         (_GEN_2182),
  ._GEN_1817                         (_GEN_2215),
  ._GEN_1818                         (_GEN_2248),
  ._GEN_1819                         (_GEN_2281),
  ._GEN_1820                         (_GEN_1853),
  ._GEN_1821                         (_GEN_1886),
  ._GEN_1822                         (_GEN_1919),
  ._GEN_1823                         (_GEN_1952),
  ._GEN_1824                         (_GEN_1985),
  ._GEN_1825                         (_GEN_2018),
  ._GEN_1826                         (_GEN_2051),
  ._GEN_1827                         (_GEN_2084),
  ._GEN_1828                         (_GEN_2117),
  ._GEN_1829                         (_GEN_2150),
  ._GEN_1830                         (_GEN_2183),
  ._GEN_1831                         (_GEN_2216),
  ._GEN_1832                         (_GEN_2249),
  ._GEN_1833                         (_GEN_2282),
  ._GEN_1834                         (_GEN_1854),
  .rob_uop_3_31_pdst                 (rob_uop_3_31_pdst),
  .rob_uop_3_30_pdst                 (rob_uop_3_30_pdst),
  .rob_uop_3_29_pdst                 (rob_uop_3_29_pdst),
  .rob_uop_3_28_pdst                 (rob_uop_3_28_pdst),
  .rob_uop_3_27_pdst                 (rob_uop_3_27_pdst),
  .rob_uop_3_26_pdst                 (rob_uop_3_26_pdst),
  .rob_uop_3_25_pdst                 (rob_uop_3_25_pdst),
  .rob_uop_3_24_pdst                 (rob_uop_3_24_pdst),
  .rob_uop_3_23_pdst                 (rob_uop_3_23_pdst),
  .rob_uop_3_22_pdst                 (rob_uop_3_22_pdst),
  .rob_uop_3_21_pdst                 (rob_uop_3_21_pdst),
  .rob_uop_3_20_pdst                 (rob_uop_3_20_pdst),
  .rob_uop_3_19_pdst                 (rob_uop_3_19_pdst),
  .rob_uop_3_18_pdst                 (rob_uop_3_18_pdst),
  .rob_uop_3_17_pdst                 (rob_uop_3_17_pdst),
  .rob_uop_3_16_pdst                 (rob_uop_3_16_pdst),
  .rob_uop_3_15_pdst                 (rob_uop_3_15_pdst),
  .rob_uop_3_14_pdst                 (rob_uop_3_14_pdst),
  .rob_uop_3_13_pdst                 (rob_uop_3_13_pdst),
  .rob_uop_3_12_pdst                 (rob_uop_3_12_pdst),
  .rob_uop_3_11_pdst                 (rob_uop_3_11_pdst),
  .rob_uop_3_10_pdst                 (rob_uop_3_10_pdst),
  .rob_uop_3_9_pdst                  (rob_uop_3_9_pdst),
  .rob_uop_3_8_pdst                  (rob_uop_3_8_pdst),
  .rob_uop_3_7_pdst                  (rob_uop_3_7_pdst),
  .rob_uop_3_6_pdst                  (rob_uop_3_6_pdst),
  .rob_uop_3_5_pdst                  (rob_uop_3_5_pdst),
  .rob_uop_3_4_pdst                  (rob_uop_3_4_pdst),
  .rob_uop_3_3_pdst                  (rob_uop_3_3_pdst),
  .rob_uop_3_2_pdst                  (rob_uop_3_2_pdst),
  .rob_uop_3_1_pdst                  (rob_uop_3_1_pdst),
  .rob_uop_3_0_pdst                  (rob_uop_3_0_pdst),
  .rob_uop_3_31_ldst_val             (rob_uop_3_31_ldst_val),
  .rob_uop_3_30_ldst_val             (rob_uop_3_30_ldst_val),
  .rob_uop_3_29_ldst_val             (rob_uop_3_29_ldst_val),
  .rob_uop_3_28_ldst_val             (rob_uop_3_28_ldst_val),
  .rob_uop_3_27_ldst_val             (rob_uop_3_27_ldst_val),
  .rob_uop_3_26_ldst_val             (rob_uop_3_26_ldst_val),
  .rob_uop_3_25_ldst_val             (rob_uop_3_25_ldst_val),
  .rob_uop_3_24_ldst_val             (rob_uop_3_24_ldst_val),
  .rob_uop_3_23_ldst_val             (rob_uop_3_23_ldst_val),
  .rob_uop_3_22_ldst_val             (rob_uop_3_22_ldst_val),
  .rob_uop_3_21_ldst_val             (rob_uop_3_21_ldst_val),
  .rob_uop_3_20_ldst_val             (rob_uop_3_20_ldst_val),
  .rob_uop_3_19_ldst_val             (rob_uop_3_19_ldst_val),
  .rob_uop_3_18_ldst_val             (rob_uop_3_18_ldst_val),
  .rob_uop_3_17_ldst_val             (rob_uop_3_17_ldst_val),
  .rob_uop_3_16_ldst_val             (rob_uop_3_16_ldst_val),
  .rob_uop_3_15_ldst_val             (rob_uop_3_15_ldst_val),
  .rob_uop_3_14_ldst_val             (rob_uop_3_14_ldst_val),
  .rob_uop_3_13_ldst_val             (rob_uop_3_13_ldst_val),
  .rob_uop_3_12_ldst_val             (rob_uop_3_12_ldst_val),
  .rob_uop_3_11_ldst_val             (rob_uop_3_11_ldst_val),
  .rob_uop_3_10_ldst_val             (rob_uop_3_10_ldst_val),
  .rob_uop_3_9_ldst_val              (rob_uop_3_9_ldst_val),
  .rob_uop_3_8_ldst_val              (rob_uop_3_8_ldst_val),
  .rob_uop_3_7_ldst_val              (rob_uop_3_7_ldst_val),
  .rob_uop_3_6_ldst_val              (rob_uop_3_6_ldst_val),
  .rob_uop_3_5_ldst_val              (rob_uop_3_5_ldst_val),
  .rob_uop_3_4_ldst_val              (rob_uop_3_4_ldst_val),
  .rob_uop_3_3_ldst_val              (rob_uop_3_3_ldst_val),
  .rob_uop_3_2_ldst_val              (rob_uop_3_2_ldst_val),
  .rob_uop_3_1_ldst_val              (rob_uop_3_1_ldst_val),
  .rob_uop_3_0_ldst_val              (rob_uop_3_0_ldst_val),
  ._GEN_1835                         (_GEN_1920),
  ._GEN_1836                         (_GEN_1986),
  ._GEN_1837                         (_GEN_2052),
  ._GEN_1838                         (_GEN_2118),
  .flush_commit_mask_3               (flush_commit_mask_3),
  .flush_commit_mask_2               (flush_commit_mask_2),
  .flush_commit_mask_1               (flush_commit_mask_1),
  .flush_commit_mask_0               (flush_commit_mask_0),
  .rob_head_fflags_0                 (casez_tmp_29),
  ._rob_uop_com_idx_fp_val           (casez_tmp_27),
  ._fflags_val_0_T                   (_fflags_val_0_T),
  ._io_commit_uops_0_uses_ldq_output (casez_tmp_20),
  ._io_commit_uops_0_uses_stq_output (casez_tmp_21),
  .rob_head_fflags_1                 (casez_tmp_49),
  ._rob_uop_1_com_idx_fp_val         (casez_tmp_47),
  ._fflags_val_1_T                   (_fflags_val_1_T),
  ._io_commit_uops_1_uses_ldq_output (casez_tmp_40),
  ._io_commit_uops_1_uses_stq_output (casez_tmp_41),
  .rob_head_fflags_2                 (casez_tmp_69),
  ._rob_uop_2_com_idx_fp_val         (casez_tmp_67),
  ._fflags_val_2_T                   (_fflags_val_2_T),
  ._io_commit_uops_2_uses_ldq_output (casez_tmp_60),
  ._io_commit_uops_2_uses_stq_output (casez_tmp_61),
  .rob_head_fflags_3                 (casez_tmp_89),
  ._rob_uop_3_com_idx_fp_val         (casez_tmp_87),
  ._fflags_val_3_T                   (_fflags_val_3_T),
  ._io_commit_uops_3_uses_ldq_output (casez_tmp_80),
  ._io_commit_uops_3_uses_stq_output (casez_tmp_81),
  .exception_thrown                  (exception_thrown),
  ._io_ready_T_3                     (~r_xcpt_val),
  .empty                             (empty),
  .r_xcpt_val                        (r_xcpt_val),
  .rob_head                          (rob_head),
  .r_xcpt_uop_rob_idx                (r_xcpt_uop_rob_idx),
  .rob_tail_idx                      (rob_tail_idx),
  .reset                             (reset),
  .full                              (full),
  ._maybe_full_T                     (~rob_deq),
  ._io_ready_T                       (_io_ready_T),
  .rob_state                         (rob_state),
  ._GEN_1839                         (|_GEN_2284),
  .rob_exception_3_31                (rob_exception_3_31),
  .rob_exception_3_30                (rob_exception_3_30),
  .rob_exception_3_29                (rob_exception_3_29),
  .rob_exception_3_28                (rob_exception_3_28),
  .rob_exception_3_27                (rob_exception_3_27),
  .rob_exception_3_26                (rob_exception_3_26),
  .rob_exception_3_25                (rob_exception_3_25),
  .rob_exception_3_24                (rob_exception_3_24),
  .rob_exception_3_23                (rob_exception_3_23),
  .rob_exception_3_22                (rob_exception_3_22),
  .rob_exception_3_21                (rob_exception_3_21),
  .rob_exception_3_20                (rob_exception_3_20),
  .rob_exception_3_19                (rob_exception_3_19),
  .rob_exception_3_18                (rob_exception_3_18),
  .rob_exception_3_17                (rob_exception_3_17),
  .rob_exception_3_16                (rob_exception_3_16),
  .rob_exception_3_15                (rob_exception_3_15),
  .rob_exception_3_14                (rob_exception_3_14),
  .rob_exception_3_13                (rob_exception_3_13),
  .rob_exception_3_12                (rob_exception_3_12),
  .rob_exception_3_11                (rob_exception_3_11),
  .rob_exception_3_10                (rob_exception_3_10),
  .rob_exception_3_9                 (rob_exception_3_9),
  .rob_exception_3_8                 (rob_exception_3_8),
  .rob_exception_3_7                 (rob_exception_3_7),
  .rob_exception_3_6                 (rob_exception_3_6),
  .rob_exception_3_5                 (rob_exception_3_5),
  .rob_exception_3_4                 (rob_exception_3_4),
  .rob_exception_3_3                 (rob_exception_3_3),
  .rob_exception_3_2                 (rob_exception_3_2),
  .rob_exception_3_1                 (rob_exception_3_1),
  .rob_exception_3_0                 (rob_exception_3_0),
  .rob_exception_2_31                (rob_exception_2_31),
  .rob_exception_2_30                (rob_exception_2_30),
  .rob_exception_2_29                (rob_exception_2_29),
  .rob_exception_2_28                (rob_exception_2_28),
  .rob_exception_2_27                (rob_exception_2_27),
  .rob_exception_2_26                (rob_exception_2_26),
  .rob_exception_2_25                (rob_exception_2_25),
  .rob_exception_2_24                (rob_exception_2_24),
  .rob_exception_2_23                (rob_exception_2_23),
  .rob_exception_2_22                (rob_exception_2_22),
  .rob_exception_2_21                (rob_exception_2_21),
  .rob_exception_2_20                (rob_exception_2_20),
  .rob_exception_2_19                (rob_exception_2_19),
  .rob_exception_2_18                (rob_exception_2_18),
  .rob_exception_2_17                (rob_exception_2_17),
  .rob_exception_2_16                (rob_exception_2_16),
  .rob_exception_2_15                (rob_exception_2_15),
  .rob_exception_2_14                (rob_exception_2_14),
  .rob_exception_2_13                (rob_exception_2_13),
  .rob_exception_2_12                (rob_exception_2_12),
  .rob_exception_2_11                (rob_exception_2_11),
  .rob_exception_2_10                (rob_exception_2_10),
  .rob_exception_2_9                 (rob_exception_2_9),
  .rob_exception_2_8                 (rob_exception_2_8),
  .rob_exception_2_7                 (rob_exception_2_7),
  .rob_exception_2_6                 (rob_exception_2_6),
  .rob_exception_2_5                 (rob_exception_2_5),
  .rob_exception_2_4                 (rob_exception_2_4),
  .rob_exception_2_3                 (rob_exception_2_3),
  .rob_exception_2_2                 (rob_exception_2_2),
  .rob_exception_2_1                 (rob_exception_2_1),
  .rob_exception_2_0                 (rob_exception_2_0),
  .rob_exception_1_31                (rob_exception_1_31),
  .rob_exception_1_30                (rob_exception_1_30),
  .rob_exception_1_29                (rob_exception_1_29),
  .rob_exception_1_28                (rob_exception_1_28),
  .rob_exception_1_27                (rob_exception_1_27),
  .rob_exception_1_26                (rob_exception_1_26),
  .rob_exception_1_25                (rob_exception_1_25),
  .rob_exception_1_24                (rob_exception_1_24),
  .rob_exception_1_23                (rob_exception_1_23),
  .rob_exception_1_22                (rob_exception_1_22),
  .rob_exception_1_21                (rob_exception_1_21),
  .rob_exception_1_20                (rob_exception_1_20),
  .rob_exception_1_19                (rob_exception_1_19),
  .rob_exception_1_18                (rob_exception_1_18),
  .rob_exception_1_17                (rob_exception_1_17),
  .rob_exception_1_16                (rob_exception_1_16),
  .rob_exception_1_15                (rob_exception_1_15),
  .rob_exception_1_14                (rob_exception_1_14),
  .rob_exception_1_13                (rob_exception_1_13),
  .rob_exception_1_12                (rob_exception_1_12),
  .rob_exception_1_11                (rob_exception_1_11),
  .rob_exception_1_10                (rob_exception_1_10),
  .rob_exception_1_9                 (rob_exception_1_9),
  .rob_exception_1_8                 (rob_exception_1_8),
  .rob_exception_1_7                 (rob_exception_1_7),
  .rob_exception_1_6                 (rob_exception_1_6),
  .rob_exception_1_5                 (rob_exception_1_5),
  .rob_exception_1_4                 (rob_exception_1_4),
  .rob_exception_1_3                 (rob_exception_1_3),
  .rob_exception_1_2                 (rob_exception_1_2),
  .rob_exception_1_1                 (rob_exception_1_1),
  .rob_exception_1_0                 (rob_exception_1_0),
  .rob_exception__31                 (rob_exception__31),
  .rob_exception__30                 (rob_exception__30),
  .rob_exception__29                 (rob_exception__29),
  .rob_exception__28                 (rob_exception__28),
  .rob_exception__27                 (rob_exception__27),
  .rob_exception__26                 (rob_exception__26),
  .rob_exception__25                 (rob_exception__25),
  .rob_exception__24                 (rob_exception__24),
  .rob_exception__23                 (rob_exception__23),
  .rob_exception__22                 (rob_exception__22),
  .rob_exception__21                 (rob_exception__21),
  .rob_exception__20                 (rob_exception__20),
  .rob_exception__19                 (rob_exception__19),
  .rob_exception__18                 (rob_exception__18),
  .rob_exception__17                 (rob_exception__17),
  .rob_exception__16                 (rob_exception__16),
  .rob_exception__15                 (rob_exception__15),
  .rob_exception__14                 (rob_exception__14),
  .rob_exception__13                 (rob_exception__13),
  .rob_exception__12                 (rob_exception__12),
  .rob_exception__11                 (rob_exception__11),
  .rob_exception__10                 (rob_exception__10),
  .rob_exception__9                  (rob_exception__9),
  .rob_exception__8                  (rob_exception__8),
  .rob_exception__7                  (rob_exception__7),
  .rob_exception__6                  (rob_exception__6),
  .rob_exception__5                  (rob_exception__5),
  .rob_exception__4                  (rob_exception__4),
  .rob_exception__3                  (rob_exception__3),
  .rob_exception__2                  (rob_exception__2),
  .rob_exception__1                  (rob_exception__1),
  .rob_exception__0                  (rob_exception__0),
  ._io_ready_T_1                     (~full),
  .io_enq_valids_0                   (io_enq_valids_0),
  .io_enq_valids_1                   (io_enq_valids_1),
  .io_enq_valids_2                   (io_enq_valids_2),
  .rob_head_idx                      (rob_head_idx),
  ._GEN_1840                         (_GEN_705),
  ._GEN_1841                         (_GEN_833),
  ._GEN_1842                         (_GEN_897),
  .io_lxcpt_bits_cause               (io_lxcpt_bits_cause),
  ._GEN_1843                         (_GEN_1260),
  ._GEN_1844                         (_GEN_1326),
  ._GEN_1845                         (_GEN_1359),
  ._GEN_1846                         (_GEN_1722),
  ._GEN_1847                         (_GEN_1788),
  ._GEN_1848                         (_GEN_1821),
  .io_enq_valids_3                   (io_enq_valids_3),
  ._GEN_1849                         (_GEN_2184),
  ._GEN_1850                         (_GEN_2250),
  ._GEN_1851                         (_GEN_2283)
);
bind CSRFile CSRFile_assert CSRFile_assert (
  .io_exception      (io_exception),
  .insn_break        (insn_break),
  .insn_call         (insn_call),
  .insn_ret          (insn_ret),
  ._io_interrupt_T   (~_io_singleStep_output),
  .io_retire         (io_retire),
  .reg_singleStepped (reg_singleStepped),
  .reg_mstatus_fs    (reg_mstatus_fs),
  .reset             (reset),
  .clock             (clock),
  .set_fs_dirty      (set_fs_dirty)
);
bind BoomCore BoomCore_assert BoomCore_assert (
  .rob_io_commit_rollback                     (_rob_io_commit_rollback),
  ._dec_hazards_T_28                          (|_b1_mispredict_mask_T_10),
  .b2_mispredict                              (b2_mispredict),
  .rob_io_com_xcpt_valid                      (_rob_io_com_xcpt_valid),
  ._io_ifu_commit_valid_T                     (_io_ifu_commit_valid_T),
  .rob_io_commit_valids_2                     (_rob_io_commit_valids_2),
  .rob_io_commit_valids_3                     (_rob_io_commit_valids_3),
  ._GEN                                       (|_alu_exe_unit_io_iresp_bits_uop_dst_rtype),
  .alu_exe_unit_io_iresp_valid                (_alu_exe_unit_io_iresp_valid),
  ._rob_io_debug_wb_valids_2_T                (_rob_io_debug_wb_valids_2_T),
  ._GEN_0                                     (|_alu_exe_unit_1_io_iresp_bits_uop_dst_rtype),
  .alu_exe_unit_1_io_iresp_valid              (_alu_exe_unit_1_io_iresp_valid),
  ._rob_io_debug_wb_valids_3_T                (_rob_io_debug_wb_valids_3_T),
  ._GEN_1                                     (|_alu_exe_unit_2_io_iresp_bits_uop_dst_rtype),
  .alu_exe_unit_2_io_iresp_valid              (_alu_exe_unit_2_io_iresp_valid),
  ._rob_io_debug_wb_valids_4_T                (_rob_io_debug_wb_valids_4_T),
  ._GEN_2                                     (|_alu_exe_unit_3_io_iresp_bits_uop_dst_rtype),
  .alu_exe_unit_3_io_iresp_valid              (_alu_exe_unit_3_io_iresp_valid),
  ._rob_io_debug_wb_valids_5_T                (_rob_io_debug_wb_valids_5_T),
  .alu_exe_unit_io_iresp_bits_uop_dst_rtype   (_alu_exe_unit_io_iresp_bits_uop_dst_rtype),
  ._rob_io_debug_wb_valids_2_T_2              (~(|_alu_exe_unit_io_iresp_bits_uop_dst_rtype)),
  .alu_exe_unit_1_io_iresp_bits_uop_dst_rtype (_alu_exe_unit_1_io_iresp_bits_uop_dst_rtype),
  ._rob_io_debug_wb_valids_3_T_2              (~(|_alu_exe_unit_1_io_iresp_bits_uop_dst_rtype)),
  .alu_exe_unit_2_io_iresp_bits_uop_dst_rtype (_alu_exe_unit_2_io_iresp_bits_uop_dst_rtype),
  ._rob_io_debug_wb_valids_4_T_2              (~(|_alu_exe_unit_2_io_iresp_bits_uop_dst_rtype)),
  .alu_exe_unit_3_io_iresp_bits_uop_dst_rtype (_alu_exe_unit_3_io_iresp_bits_uop_dst_rtype),
  ._rob_io_debug_wb_valids_5_T_2              (~(|_alu_exe_unit_3_io_iresp_bits_uop_dst_rtype)),
  .FpPipeline_io_wakeups_0_valid              (_FpPipeline_io_wakeups_0_valid),
  .FpPipeline_io_wakeups_0_bits_uop_dst_rtype (_FpPipeline_io_wakeups_0_bits_uop_dst_rtype),
  .FpPipeline_io_wakeups_0_bits_uop_fp_val    (_FpPipeline_io_wakeups_0_bits_uop_fp_val),
  .FpPipeline_io_wakeups_1_valid              (_FpPipeline_io_wakeups_1_valid),
  .FpPipeline_io_wakeups_1_bits_uop_dst_rtype (_FpPipeline_io_wakeups_1_bits_uop_dst_rtype),
  .FpPipeline_io_wakeups_1_bits_uop_fp_val    (_FpPipeline_io_wakeups_1_bits_uop_fp_val),
  .FpPipeline_io_wakeups_2_valid              (_FpPipeline_io_wakeups_2_valid),
  .FpPipeline_io_wakeups_2_bits_uop_dst_rtype (_FpPipeline_io_wakeups_2_bits_uop_dst_rtype),
  .FpPipeline_io_wakeups_2_bits_uop_fp_val    (_FpPipeline_io_wakeups_2_bits_uop_fp_val),
  .FpPipeline_io_wakeups_3_valid              (_FpPipeline_io_wakeups_3_valid),
  .FpPipeline_io_wakeups_3_bits_uop_dst_rtype (_FpPipeline_io_wakeups_3_bits_uop_dst_rtype),
  .FpPipeline_io_wakeups_3_bits_uop_fp_val    (_FpPipeline_io_wakeups_3_bits_uop_fp_val),
  .csr_io_singleStep                          (_csr_io_singleStep),
  ._brinfos_3_valid_T                         (~_rob_io_flush_valid),
  .clock                                      (clock),
  .reset                                      (reset),
  .csr_io_csr_stall                           (_csr_io_csr_stall),
  .rob_io_commit_valids_1                     (_rob_io_commit_valids_1),
  .rob_io_commit_valids_0                     (_rob_io_commit_valids_0)
);
bind NBDTLB NBDTLB_assert NBDTLB_assert (
  .vpn_0               (io_req_0_bits_vaddr[38:12]),
  .io_sfence_bits_addr (io_sfence_bits_addr),
  .io_sfence_bits_rs1  (io_sfence_bits_rs1),
  .vpn_1               (io_req_1_bits_vaddr[38:12]),
  .io_sfence_valid     (io_sfence_valid),
  .reset               (reset),
  .clock               (clock)
);
bind LSU LSU_assert LSU_assert (
  .io_core_brupdate_b2_mispredict            (io_core_brupdate_b2_mispredict),
  ._stq_stq_execute_head_valid_1             (casez_tmp),
  .stq_tail                                  (stq_tail),
  .stq_execute_head                          (stq_execute_head),
  .stq_head                                  (stq_head),
  .ldq_tail                                  (ldq_tail),
  .io_core_dis_uops_0_bits_ldq_idx           (io_core_dis_uops_0_bits_ldq_idx),
  .ldq_31_valid                              (ldq_31_valid),
  .ldq_30_valid                              (ldq_30_valid),
  .ldq_29_valid                              (ldq_29_valid),
  .ldq_28_valid                              (ldq_28_valid),
  .ldq_27_valid                              (ldq_27_valid),
  .ldq_26_valid                              (ldq_26_valid),
  .ldq_25_valid                              (ldq_25_valid),
  .ldq_24_valid                              (ldq_24_valid),
  .ldq_23_valid                              (ldq_23_valid),
  .ldq_22_valid                              (ldq_22_valid),
  .ldq_21_valid                              (ldq_21_valid),
  .ldq_20_valid                              (ldq_20_valid),
  .ldq_19_valid                              (ldq_19_valid),
  .ldq_18_valid                              (ldq_18_valid),
  .ldq_17_valid                              (ldq_17_valid),
  .ldq_16_valid                              (ldq_16_valid),
  .ldq_15_valid                              (ldq_15_valid),
  .ldq_14_valid                              (ldq_14_valid),
  .ldq_13_valid                              (ldq_13_valid),
  .ldq_12_valid                              (ldq_12_valid),
  .ldq_11_valid                              (ldq_11_valid),
  .ldq_10_valid                              (ldq_10_valid),
  .ldq_9_valid                               (ldq_9_valid),
  .ldq_8_valid                               (ldq_8_valid),
  .ldq_7_valid                               (ldq_7_valid),
  .ldq_6_valid                               (ldq_6_valid),
  .ldq_5_valid                               (ldq_5_valid),
  .ldq_4_valid                               (ldq_4_valid),
  .ldq_3_valid                               (ldq_3_valid),
  .ldq_2_valid                               (ldq_2_valid),
  .ldq_1_valid                               (ldq_1_valid),
  .ldq_0_valid                               (ldq_0_valid),
  .io_core_dis_uops_0_bits_stq_idx           (io_core_dis_uops_0_bits_stq_idx),
  .stq_31_valid                              (stq_31_valid),
  .stq_30_valid                              (stq_30_valid),
  .stq_29_valid                              (stq_29_valid),
  .stq_28_valid                              (stq_28_valid),
  .stq_27_valid                              (stq_27_valid),
  .stq_26_valid                              (stq_26_valid),
  .stq_25_valid                              (stq_25_valid),
  .stq_24_valid                              (stq_24_valid),
  .stq_23_valid                              (stq_23_valid),
  .stq_22_valid                              (stq_22_valid),
  .stq_21_valid                              (stq_21_valid),
  .stq_20_valid                              (stq_20_valid),
  .stq_19_valid                              (stq_19_valid),
  .stq_18_valid                              (stq_18_valid),
  .stq_17_valid                              (stq_17_valid),
  .stq_16_valid                              (stq_16_valid),
  .stq_15_valid                              (stq_15_valid),
  .stq_14_valid                              (stq_14_valid),
  .stq_13_valid                              (stq_13_valid),
  .stq_12_valid                              (stq_12_valid),
  .stq_11_valid                              (stq_11_valid),
  .stq_10_valid                              (stq_10_valid),
  .stq_9_valid                               (stq_9_valid),
  .stq_8_valid                               (stq_8_valid),
  .stq_7_valid                               (stq_7_valid),
  .stq_6_valid                               (stq_6_valid),
  .stq_5_valid                               (stq_5_valid),
  .stq_4_valid                               (stq_4_valid),
  .stq_3_valid                               (stq_3_valid),
  .stq_2_valid                               (stq_2_valid),
  .stq_1_valid                               (stq_1_valid),
  .stq_0_valid                               (stq_0_valid),
  .dis_ld_val                                (dis_ld_val),
  .dis_st_val                                (dis_st_val),
  ._GEN                                      (_GEN_66),
  .io_core_dis_uops_1_bits_ldq_idx           (io_core_dis_uops_1_bits_ldq_idx),
  ._ldq_T_35_bits_youngest_stq_idx           (_ldq_T_35_bits_youngest_stq_idx),
  .io_core_dis_uops_1_bits_stq_idx           (io_core_dis_uops_1_bits_stq_idx),
  .dis_ld_val_1                              (dis_ld_val_1),
  .dis_st_val_1                              (dis_st_val_1),
  ._GEN_0                                    (_GEN_164),
  .io_core_dis_uops_2_bits_ldq_idx           (io_core_dis_uops_2_bits_ldq_idx),
  ._ldq_T_75_bits_youngest_stq_idx           (_ldq_T_75_bits_youngest_stq_idx),
  .io_core_dis_uops_2_bits_stq_idx           (io_core_dis_uops_2_bits_stq_idx),
  .dis_ld_val_2                              (dis_ld_val_2),
  .dis_st_val_2                              (dis_st_val_2),
  ._GEN_1                                    (_GEN_231),
  .io_core_dis_uops_3_bits_ldq_idx           (io_core_dis_uops_3_bits_ldq_idx),
  ._ldq_T_115_bits_youngest_stq_idx          (_ldq_T_115_bits_youngest_stq_idx),
  .io_core_dis_uops_3_bits_stq_idx           (io_core_dis_uops_3_bits_stq_idx),
  .dis_ld_val_3                              (dis_ld_val_3),
  .dis_st_val_3                              (dis_st_val_3),
  .exe_req_0_valid                           (exe_req_0_valid),
  .will_fire_std_incoming_0                  (will_fire_std_incoming_0),
  .will_fire_sfence_0                        (will_fire_sfence_0),
  ._exe_cmd_T                                (_exe_cmd_T),
  .will_fire_sta_incoming_0                  (will_fire_sta_incoming_0),
  .exe_req_1_valid                           (exe_req_1_valid),
  .will_fire_std_incoming_1                  (will_fire_std_incoming_1),
  .will_fire_sfence_1                        (will_fire_sfence_1),
  ._exe_cmd_T_7                              (_exe_cmd_T_7),
  .will_fire_sta_incoming_1                  (will_fire_sta_incoming_1),
  ._GEN_2                                    (|hella_state),
  .hella_req_cmd                             (hella_req_cmd),
  .exe_tlb_valid_0                           (~_will_fire_store_commit_0_T_2),
  ._exe_tlb_uop_T_2                          (_exe_tlb_uop_T_2),
  .io_core_exe_1_req_bits_sfence_valid       (io_core_exe_1_req_bits_sfence_valid),
  .io_core_exe_1_req_bits_uop_is_fence       (io_core_exe_1_req_bits_uop_is_fence),
  .io_core_exe_0_req_bits_uop_is_fence       (io_core_exe_0_req_bits_uop_is_fence),
  .exe_req_0_bits_mxcpt_valid                (exe_req_0_bits_mxcpt_valid),
  .mem_incoming_uop_out_ctrl_is_sta          (mem_incoming_uop_out_ctrl_is_sta),
  .mem_incoming_uop_out_ctrl_is_load         (mem_incoming_uop_out_ctrl_is_load),
  .can_fire_load_incoming_0                  (can_fire_load_incoming_0),
  .will_fire_stad_incoming_0                 (will_fire_stad_incoming_0),
  .exe_tlb_valid_1                           (~_will_fire_store_commit_1_T_2),
  ._exe_tlb_uop_T_9                          (_exe_tlb_uop_T_9),
  .will_fire_load_retry_1                    (will_fire_load_retry_1),
  .will_fire_sta_retry_1                     (will_fire_sta_retry_1),
  .stq_retry_idx                             (stq_retry_idx),
  .stq_31_bits_uop_is_fence                  (stq_31_bits_uop_is_fence),
  .stq_30_bits_uop_is_fence                  (stq_30_bits_uop_is_fence),
  .stq_29_bits_uop_is_fence                  (stq_29_bits_uop_is_fence),
  .stq_28_bits_uop_is_fence                  (stq_28_bits_uop_is_fence),
  .stq_27_bits_uop_is_fence                  (stq_27_bits_uop_is_fence),
  .stq_26_bits_uop_is_fence                  (stq_26_bits_uop_is_fence),
  .stq_25_bits_uop_is_fence                  (stq_25_bits_uop_is_fence),
  .stq_24_bits_uop_is_fence                  (stq_24_bits_uop_is_fence),
  .stq_23_bits_uop_is_fence                  (stq_23_bits_uop_is_fence),
  .stq_22_bits_uop_is_fence                  (stq_22_bits_uop_is_fence),
  .stq_21_bits_uop_is_fence                  (stq_21_bits_uop_is_fence),
  .stq_20_bits_uop_is_fence                  (stq_20_bits_uop_is_fence),
  .stq_19_bits_uop_is_fence                  (stq_19_bits_uop_is_fence),
  .stq_18_bits_uop_is_fence                  (stq_18_bits_uop_is_fence),
  .stq_17_bits_uop_is_fence                  (stq_17_bits_uop_is_fence),
  .stq_16_bits_uop_is_fence                  (stq_16_bits_uop_is_fence),
  .stq_15_bits_uop_is_fence                  (stq_15_bits_uop_is_fence),
  .stq_14_bits_uop_is_fence                  (stq_14_bits_uop_is_fence),
  .stq_13_bits_uop_is_fence                  (stq_13_bits_uop_is_fence),
  .stq_12_bits_uop_is_fence                  (stq_12_bits_uop_is_fence),
  .stq_11_bits_uop_is_fence                  (stq_11_bits_uop_is_fence),
  .stq_10_bits_uop_is_fence                  (stq_10_bits_uop_is_fence),
  .stq_9_bits_uop_is_fence                   (stq_9_bits_uop_is_fence),
  .stq_8_bits_uop_is_fence                   (stq_8_bits_uop_is_fence),
  .stq_7_bits_uop_is_fence                   (stq_7_bits_uop_is_fence),
  .stq_6_bits_uop_is_fence                   (stq_6_bits_uop_is_fence),
  .stq_5_bits_uop_is_fence                   (stq_5_bits_uop_is_fence),
  .stq_4_bits_uop_is_fence                   (stq_4_bits_uop_is_fence),
  .stq_3_bits_uop_is_fence                   (stq_3_bits_uop_is_fence),
  .stq_2_bits_uop_is_fence                   (stq_2_bits_uop_is_fence),
  .stq_1_bits_uop_is_fence                   (stq_1_bits_uop_is_fence),
  .stq_0_bits_uop_is_fence                   (stq_0_bits_uop_is_fence),
  .ldq_retry_idx                             (ldq_retry_idx),
  .clock                                     (clock),
  ._GEN_3                                    (_GEN_297),
  .io_core_dis_uops_3_bits_is_fence          (io_core_dis_uops_3_bits_is_fence),
  ._GEN_4                                    (_GEN_199),
  .io_core_dis_uops_2_bits_is_fence          (io_core_dis_uops_2_bits_is_fence),
  ._GEN_5                                    (_GEN_132),
  .io_core_dis_uops_1_bits_is_fence          (io_core_dis_uops_1_bits_is_fence),
  ._GEN_6                                    (_GEN_34),
  .io_core_dis_uops_0_bits_is_fence          (io_core_dis_uops_0_bits_is_fence),
  ._GEN_7                                    (_GEN_298),
  ._GEN_8                                    (_GEN_200),
  ._GEN_9                                    (_GEN_133),
  ._GEN_10                                   (_GEN_35),
  ._GEN_11                                   (_GEN_299),
  ._GEN_12                                   (_GEN_201),
  ._GEN_13                                   (_GEN_134),
  ._GEN_14                                   (_GEN_36),
  ._GEN_15                                   (_GEN_300),
  ._GEN_16                                   (_GEN_202),
  ._GEN_17                                   (_GEN_135),
  ._GEN_18                                   (_GEN_37),
  ._GEN_19                                   (_GEN_301),
  ._GEN_20                                   (_GEN_203),
  ._GEN_21                                   (_GEN_136),
  ._GEN_22                                   (_GEN_38),
  ._GEN_23                                   (_GEN_302),
  ._GEN_24                                   (_GEN_204),
  ._GEN_25                                   (_GEN_137),
  ._GEN_26                                   (_GEN_39),
  ._GEN_27                                   (_GEN_303),
  ._GEN_28                                   (_GEN_205),
  ._GEN_29                                   (_GEN_138),
  ._GEN_30                                   (_GEN_40),
  ._GEN_31                                   (_GEN_304),
  ._GEN_32                                   (_GEN_206),
  ._GEN_33                                   (_GEN_139),
  ._GEN_34                                   (_GEN_41),
  ._GEN_35                                   (_GEN_305),
  ._GEN_36                                   (_GEN_207),
  ._GEN_37                                   (_GEN_140),
  ._GEN_38                                   (_GEN_42),
  ._GEN_39                                   (_GEN_306),
  ._GEN_40                                   (_GEN_208),
  ._GEN_41                                   (_GEN_141),
  ._GEN_42                                   (_GEN_43),
  ._GEN_43                                   (_GEN_307),
  ._GEN_44                                   (_GEN_209),
  ._GEN_45                                   (_GEN_142),
  ._GEN_46                                   (_GEN_44),
  ._GEN_47                                   (_GEN_308),
  ._GEN_48                                   (_GEN_210),
  ._GEN_49                                   (_GEN_143),
  ._GEN_50                                   (_GEN_45),
  ._GEN_51                                   (_GEN_309),
  ._GEN_52                                   (_GEN_211),
  ._GEN_53                                   (_GEN_144),
  ._GEN_54                                   (_GEN_46),
  ._GEN_55                                   (_GEN_310),
  ._GEN_56                                   (_GEN_212),
  ._GEN_57                                   (_GEN_145),
  ._GEN_58                                   (_GEN_47),
  ._GEN_59                                   (_GEN_311),
  ._GEN_60                                   (_GEN_213),
  ._GEN_61                                   (_GEN_146),
  ._GEN_62                                   (_GEN_48),
  ._GEN_63                                   (_GEN_312),
  ._GEN_64                                   (_GEN_214),
  ._GEN_65                                   (_GEN_147),
  ._GEN_66                                   (_GEN_49),
  ._GEN_67                                   (_GEN_313),
  ._GEN_68                                   (_GEN_215),
  ._GEN_69                                   (_GEN_148),
  ._GEN_70                                   (_GEN_50),
  ._GEN_71                                   (_GEN_314),
  ._GEN_72                                   (_GEN_216),
  ._GEN_73                                   (_GEN_149),
  ._GEN_74                                   (_GEN_51),
  ._GEN_75                                   (_GEN_315),
  ._GEN_76                                   (_GEN_217),
  ._GEN_77                                   (_GEN_150),
  ._GEN_78                                   (_GEN_52),
  ._GEN_79                                   (_GEN_316),
  ._GEN_80                                   (_GEN_218),
  ._GEN_81                                   (_GEN_151),
  ._GEN_82                                   (_GEN_53),
  ._GEN_83                                   (_GEN_317),
  ._GEN_84                                   (_GEN_219),
  ._GEN_85                                   (_GEN_152),
  ._GEN_86                                   (_GEN_54),
  ._GEN_87                                   (_GEN_318),
  ._GEN_88                                   (_GEN_220),
  ._GEN_89                                   (_GEN_153),
  ._GEN_90                                   (_GEN_55),
  ._GEN_91                                   (_GEN_319),
  ._GEN_92                                   (_GEN_221),
  ._GEN_93                                   (_GEN_154),
  ._GEN_94                                   (_GEN_56),
  ._GEN_95                                   (_GEN_320),
  ._GEN_96                                   (_GEN_222),
  ._GEN_97                                   (_GEN_155),
  ._GEN_98                                   (_GEN_57),
  ._GEN_99                                   (_GEN_321),
  ._GEN_100                                  (_GEN_223),
  ._GEN_101                                  (_GEN_156),
  ._GEN_102                                  (_GEN_58),
  ._GEN_103                                  (_GEN_322),
  ._GEN_104                                  (_GEN_224),
  ._GEN_105                                  (_GEN_157),
  ._GEN_106                                  (_GEN_59),
  ._GEN_107                                  (_GEN_323),
  ._GEN_108                                  (_GEN_225),
  ._GEN_109                                  (_GEN_158),
  ._GEN_110                                  (_GEN_60),
  ._GEN_111                                  (_GEN_324),
  ._GEN_112                                  (_GEN_226),
  ._GEN_113                                  (_GEN_159),
  ._GEN_114                                  (_GEN_61),
  ._GEN_115                                  (_GEN_325),
  ._GEN_116                                  (_GEN_227),
  ._GEN_117                                  (_GEN_160),
  ._GEN_118                                  (_GEN_62),
  ._GEN_119                                  (_GEN_326),
  ._GEN_120                                  (_GEN_228),
  ._GEN_121                                  (_GEN_161),
  ._GEN_122                                  (_GEN_63),
  ._GEN_123                                  (_GEN_327),
  ._GEN_124                                  (_GEN_229),
  ._GEN_125                                  (_GEN_162),
  ._GEN_126                                  (_GEN_64),
  ._GEN_127                                  (_GEN_328),
  ._GEN_128                                  (_GEN_230),
  ._GEN_129                                  (_GEN_163),
  ._GEN_130                                  (_GEN_65),
  .io_core_exe_0_req_bits_sfence_valid       (io_core_exe_0_req_bits_sfence_valid),
  .exe_req_1_bits_mxcpt_valid                (exe_req_1_bits_mxcpt_valid),
  .exe_req_1_bits_uop_ctrl_is_sta            (exe_req_1_bits_uop_ctrl_is_sta),
  .io_core_dis_uops_3_bits_ctrl_is_sta       (io_core_dis_uops_3_bits_ctrl_is_sta),
  .io_core_dis_uops_2_bits_ctrl_is_sta       (io_core_dis_uops_2_bits_ctrl_is_sta),
  .io_core_dis_uops_1_bits_ctrl_is_sta       (io_core_dis_uops_1_bits_ctrl_is_sta),
  .io_core_dis_uops_0_bits_ctrl_is_sta       (io_core_dis_uops_0_bits_ctrl_is_sta),
  ._GEN_131                                  (_GEN_2),
  ._GEN_132                                  (_GEN_100),
  ._GEN_133                                  (_GEN_167),
  ._GEN_134                                  (_GEN_265),
  ._GEN_135                                  (_GEN_1235),
  ._GEN_136                                  (_GEN_3),
  ._GEN_137                                  (_GEN_101),
  ._GEN_138                                  (_GEN_168),
  ._GEN_139                                  (_GEN_266),
  ._GEN_140                                  (_GEN_4),
  ._GEN_141                                  (_GEN_102),
  ._GEN_142                                  (_GEN_169),
  ._GEN_143                                  (_GEN_267),
  ._GEN_144                                  (_GEN_5),
  ._GEN_145                                  (_GEN_103),
  ._GEN_146                                  (_GEN_170),
  ._GEN_147                                  (_GEN_268),
  ._GEN_148                                  (_GEN_6),
  ._GEN_149                                  (_GEN_104),
  ._GEN_150                                  (_GEN_171),
  ._GEN_151                                  (_GEN_269),
  ._GEN_152                                  (_GEN_7),
  ._GEN_153                                  (_GEN_105),
  ._GEN_154                                  (_GEN_172),
  ._GEN_155                                  (_GEN_270),
  ._GEN_156                                  (_GEN_8),
  ._GEN_157                                  (_GEN_106),
  ._GEN_158                                  (_GEN_173),
  ._GEN_159                                  (_GEN_271),
  ._GEN_160                                  (_GEN_9),
  ._GEN_161                                  (_GEN_107),
  ._GEN_162                                  (_GEN_174),
  ._GEN_163                                  (_GEN_272),
  ._GEN_164                                  (_GEN_10),
  ._GEN_165                                  (_GEN_108),
  ._GEN_166                                  (_GEN_175),
  ._GEN_167                                  (_GEN_273),
  ._GEN_168                                  (_GEN_11),
  ._GEN_169                                  (_GEN_109),
  ._GEN_170                                  (_GEN_176),
  ._GEN_171                                  (_GEN_274),
  ._GEN_172                                  (_GEN_12),
  ._GEN_173                                  (_GEN_110),
  ._GEN_174                                  (_GEN_177),
  ._GEN_175                                  (_GEN_275),
  ._GEN_176                                  (_GEN_13),
  ._GEN_177                                  (_GEN_111),
  ._GEN_178                                  (_GEN_178),
  ._GEN_179                                  (_GEN_276),
  ._GEN_180                                  (_GEN_14),
  ._GEN_181                                  (_GEN_112),
  ._GEN_182                                  (_GEN_179),
  ._GEN_183                                  (_GEN_277),
  ._GEN_184                                  (_GEN_15),
  ._GEN_185                                  (_GEN_113),
  ._GEN_186                                  (_GEN_180),
  ._GEN_187                                  (_GEN_278),
  ._GEN_188                                  (_GEN_16),
  ._GEN_189                                  (_GEN_114),
  ._GEN_190                                  (_GEN_181),
  ._GEN_191                                  (_GEN_279),
  ._GEN_192                                  (_GEN_17),
  ._GEN_193                                  (_GEN_115),
  ._GEN_194                                  (_GEN_182),
  ._GEN_195                                  (_GEN_280),
  ._GEN_196                                  (_GEN_18),
  ._GEN_197                                  (_GEN_116),
  ._GEN_198                                  (_GEN_183),
  ._GEN_199                                  (_GEN_281),
  ._GEN_200                                  (_GEN_19),
  ._GEN_201                                  (_GEN_117),
  ._GEN_202                                  (_GEN_184),
  ._GEN_203                                  (_GEN_282),
  ._GEN_204                                  (_GEN_20),
  ._GEN_205                                  (_GEN_118),
  ._GEN_206                                  (_GEN_185),
  ._GEN_207                                  (_GEN_283),
  ._GEN_208                                  (_GEN_21),
  ._GEN_209                                  (_GEN_119),
  ._GEN_210                                  (_GEN_186),
  ._GEN_211                                  (_GEN_284),
  ._GEN_212                                  (_GEN_22),
  ._GEN_213                                  (_GEN_120),
  ._GEN_214                                  (_GEN_187),
  ._GEN_215                                  (_GEN_285),
  ._GEN_216                                  (_GEN_23),
  ._GEN_217                                  (_GEN_121),
  ._GEN_218                                  (_GEN_188),
  ._GEN_219                                  (_GEN_286),
  ._GEN_220                                  (_GEN_24),
  ._GEN_221                                  (_GEN_122),
  ._GEN_222                                  (_GEN_189),
  ._GEN_223                                  (_GEN_287),
  ._GEN_224                                  (_GEN_25),
  ._GEN_225                                  (_GEN_123),
  ._GEN_226                                  (_GEN_190),
  ._GEN_227                                  (_GEN_288),
  ._GEN_228                                  (_GEN_26),
  ._GEN_229                                  (_GEN_124),
  ._GEN_230                                  (_GEN_191),
  ._GEN_231                                  (_GEN_289),
  ._GEN_232                                  (_GEN_27),
  ._GEN_233                                  (_GEN_125),
  ._GEN_234                                  (_GEN_192),
  ._GEN_235                                  (_GEN_290),
  ._GEN_236                                  (_GEN_28),
  ._GEN_237                                  (_GEN_126),
  ._GEN_238                                  (_GEN_193),
  ._GEN_239                                  (_GEN_291),
  ._GEN_240                                  (_GEN_29),
  ._GEN_241                                  (_GEN_127),
  ._GEN_242                                  (_GEN_194),
  ._GEN_243                                  (_GEN_292),
  ._GEN_244                                  (_GEN_30),
  ._GEN_245                                  (_GEN_128),
  ._GEN_246                                  (_GEN_195),
  ._GEN_247                                  (_GEN_293),
  ._GEN_248                                  (_GEN_31),
  ._GEN_249                                  (_GEN_129),
  ._GEN_250                                  (_GEN_196),
  ._GEN_251                                  (_GEN_294),
  ._GEN_252                                  (_GEN_32),
  ._GEN_253                                  (_GEN_130),
  ._GEN_254                                  (_GEN_197),
  ._GEN_255                                  (_GEN_295),
  ._GEN_256                                  (_GEN_33),
  ._GEN_257                                  (_GEN_131),
  ._GEN_258                                  (_GEN_198),
  ._GEN_259                                  (_GEN_296),
  .exe_req_1_bits_uop_ctrl_is_load           (exe_req_1_bits_uop_ctrl_is_load),
  .io_core_dis_uops_3_bits_ctrl_is_load      (io_core_dis_uops_3_bits_ctrl_is_load),
  .io_core_dis_uops_2_bits_ctrl_is_load      (io_core_dis_uops_2_bits_ctrl_is_load),
  .io_core_dis_uops_1_bits_ctrl_is_load      (io_core_dis_uops_1_bits_ctrl_is_load),
  .io_core_dis_uops_0_bits_ctrl_is_load      (io_core_dis_uops_0_bits_ctrl_is_load),
  .can_fire_load_incoming_1                  (can_fire_load_incoming_1),
  .will_fire_stad_incoming_1                 (will_fire_stad_incoming_1),
  .exe_req_0_bits_sfence_valid               (exe_req_0_bits_sfence_valid),
  .exe_tlb_paddr_0                           (exe_tlb_paddr_0),
  .dtlb_io_resp_0_paddr                      (_dtlb_io_resp_0_paddr),
  .mem_xcpt_uops_0_uses_ldq                  (mem_xcpt_uops_0_uses_ldq),
  .exe_tlb_uop_0_uses_stq                    (exe_tlb_uop_0_uses_stq),
  .exe_req_1_bits_sfence_valid               (exe_req_1_bits_sfence_valid),
  .exe_tlb_paddr_1                           (exe_tlb_paddr_1),
  .dtlb_io_resp_1_paddr                      (_dtlb_io_resp_1_paddr),
  .mem_xcpt_uops_1_uses_ldq                  (mem_xcpt_uops_1_uses_ldq),
  .exe_tlb_uop_1_uses_stq                    (exe_tlb_uop_1_uses_stq),
  .ldq_incoming_idx_0                        (ldq_incoming_idx_0),
  .ldq_31_bits_executed                      (ldq_31_bits_executed),
  .ldq_30_bits_executed                      (ldq_30_bits_executed),
  .ldq_29_bits_executed                      (ldq_29_bits_executed),
  .ldq_28_bits_executed                      (ldq_28_bits_executed),
  .ldq_27_bits_executed                      (ldq_27_bits_executed),
  .ldq_26_bits_executed                      (ldq_26_bits_executed),
  .ldq_25_bits_executed                      (ldq_25_bits_executed),
  .ldq_24_bits_executed                      (ldq_24_bits_executed),
  .ldq_23_bits_executed                      (ldq_23_bits_executed),
  .ldq_22_bits_executed                      (ldq_22_bits_executed),
  .ldq_21_bits_executed                      (ldq_21_bits_executed),
  .ldq_20_bits_executed                      (ldq_20_bits_executed),
  .ldq_19_bits_executed                      (ldq_19_bits_executed),
  .ldq_18_bits_executed                      (ldq_18_bits_executed),
  .ldq_17_bits_executed                      (ldq_17_bits_executed),
  .ldq_16_bits_executed                      (ldq_16_bits_executed),
  .ldq_15_bits_executed                      (ldq_15_bits_executed),
  .ldq_14_bits_executed                      (ldq_14_bits_executed),
  .ldq_13_bits_executed                      (ldq_13_bits_executed),
  .ldq_12_bits_executed                      (ldq_12_bits_executed),
  .ldq_11_bits_executed                      (ldq_11_bits_executed),
  .ldq_10_bits_executed                      (ldq_10_bits_executed),
  .ldq_9_bits_executed                       (ldq_9_bits_executed),
  .ldq_8_bits_executed                       (ldq_8_bits_executed),
  .ldq_7_bits_executed                       (ldq_7_bits_executed),
  .ldq_6_bits_executed                       (ldq_6_bits_executed),
  .ldq_5_bits_executed                       (ldq_5_bits_executed),
  .ldq_4_bits_executed                       (ldq_4_bits_executed),
  .ldq_3_bits_executed                       (ldq_3_bits_executed),
  .ldq_2_bits_executed                       (ldq_2_bits_executed),
  .ldq_1_bits_executed                       (ldq_1_bits_executed),
  .ldq_0_bits_executed                       (ldq_0_bits_executed),
  .ldq_31_bits_addr_valid                    (ldq_31_bits_addr_valid),
  .ldq_30_bits_addr_valid                    (ldq_30_bits_addr_valid),
  .ldq_29_bits_addr_valid                    (ldq_29_bits_addr_valid),
  .ldq_28_bits_addr_valid                    (ldq_28_bits_addr_valid),
  .ldq_27_bits_addr_valid                    (ldq_27_bits_addr_valid),
  .ldq_26_bits_addr_valid                    (ldq_26_bits_addr_valid),
  .ldq_25_bits_addr_valid                    (ldq_25_bits_addr_valid),
  .ldq_24_bits_addr_valid                    (ldq_24_bits_addr_valid),
  .ldq_23_bits_addr_valid                    (ldq_23_bits_addr_valid),
  .ldq_22_bits_addr_valid                    (ldq_22_bits_addr_valid),
  .ldq_21_bits_addr_valid                    (ldq_21_bits_addr_valid),
  .ldq_20_bits_addr_valid                    (ldq_20_bits_addr_valid),
  .ldq_19_bits_addr_valid                    (ldq_19_bits_addr_valid),
  .ldq_18_bits_addr_valid                    (ldq_18_bits_addr_valid),
  .ldq_17_bits_addr_valid                    (ldq_17_bits_addr_valid),
  .ldq_16_bits_addr_valid                    (ldq_16_bits_addr_valid),
  .ldq_15_bits_addr_valid                    (ldq_15_bits_addr_valid),
  .ldq_14_bits_addr_valid                    (ldq_14_bits_addr_valid),
  .ldq_13_bits_addr_valid                    (ldq_13_bits_addr_valid),
  .ldq_12_bits_addr_valid                    (ldq_12_bits_addr_valid),
  .ldq_11_bits_addr_valid                    (ldq_11_bits_addr_valid),
  .ldq_10_bits_addr_valid                    (ldq_10_bits_addr_valid),
  .ldq_9_bits_addr_valid                     (ldq_9_bits_addr_valid),
  .ldq_8_bits_addr_valid                     (ldq_8_bits_addr_valid),
  .ldq_7_bits_addr_valid                     (ldq_7_bits_addr_valid),
  .ldq_6_bits_addr_valid                     (ldq_6_bits_addr_valid),
  .ldq_5_bits_addr_valid                     (ldq_5_bits_addr_valid),
  .ldq_4_bits_addr_valid                     (ldq_4_bits_addr_valid),
  .ldq_3_bits_addr_valid                     (ldq_3_bits_addr_valid),
  .ldq_2_bits_addr_valid                     (ldq_2_bits_addr_valid),
  .ldq_1_bits_addr_valid                     (ldq_1_bits_addr_valid),
  .ldq_0_bits_addr_valid                     (ldq_0_bits_addr_valid),
  .stq_incoming_e_0_bits_addr_valid          (casez_tmp_18),
  .sidx                                      (sidx),
  .stq_31_bits_data_valid                    (stq_31_bits_data_valid),
  .stq_30_bits_data_valid                    (stq_30_bits_data_valid),
  .stq_29_bits_data_valid                    (stq_29_bits_data_valid),
  .stq_28_bits_data_valid                    (stq_28_bits_data_valid),
  .stq_27_bits_data_valid                    (stq_27_bits_data_valid),
  .stq_26_bits_data_valid                    (stq_26_bits_data_valid),
  .stq_25_bits_data_valid                    (stq_25_bits_data_valid),
  .stq_24_bits_data_valid                    (stq_24_bits_data_valid),
  .stq_23_bits_data_valid                    (stq_23_bits_data_valid),
  .stq_22_bits_data_valid                    (stq_22_bits_data_valid),
  .stq_21_bits_data_valid                    (stq_21_bits_data_valid),
  .stq_20_bits_data_valid                    (stq_20_bits_data_valid),
  .stq_19_bits_data_valid                    (stq_19_bits_data_valid),
  .stq_18_bits_data_valid                    (stq_18_bits_data_valid),
  .stq_17_bits_data_valid                    (stq_17_bits_data_valid),
  .stq_16_bits_data_valid                    (stq_16_bits_data_valid),
  .stq_15_bits_data_valid                    (stq_15_bits_data_valid),
  .stq_14_bits_data_valid                    (stq_14_bits_data_valid),
  .stq_13_bits_data_valid                    (stq_13_bits_data_valid),
  .stq_12_bits_data_valid                    (stq_12_bits_data_valid),
  .stq_11_bits_data_valid                    (stq_11_bits_data_valid),
  .stq_10_bits_data_valid                    (stq_10_bits_data_valid),
  .stq_9_bits_data_valid                     (stq_9_bits_data_valid),
  .stq_8_bits_data_valid                     (stq_8_bits_data_valid),
  .stq_7_bits_data_valid                     (stq_7_bits_data_valid),
  .stq_6_bits_data_valid                     (stq_6_bits_data_valid),
  .stq_5_bits_data_valid                     (stq_5_bits_data_valid),
  .stq_4_bits_data_valid                     (stq_4_bits_data_valid),
  .stq_3_bits_data_valid                     (stq_3_bits_data_valid),
  .stq_2_bits_data_valid                     (stq_2_bits_data_valid),
  .stq_1_bits_data_valid                     (stq_1_bits_data_valid),
  .stq_0_bits_data_valid                     (stq_0_bits_data_valid),
  .ldq_incoming_idx_1                        (ldq_incoming_idx_1),
  .mem_ldq_wakeup_e_out_bits_addr_is_virtual (casez_tmp_33),
  .mem_ldq_wakeup_e_out_bits_executed        (casez_tmp_34),
  ._GEN_140251                               (_GEN_140251),
  ._GEN_140205                               (_GEN_140205),
  .stq_incoming_e_1_bits_addr_valid          (casez_tmp_27),
  .sidx_1                                    (sidx_1),
  ._GEN_260                                  (_GEN_331),
  ._GEN_261                                  (_GEN_1177),
  .io_dmem_nack_0_bits_uop_ldq_idx           (io_dmem_nack_0_bits_uop_ldq_idx),
  .io_dmem_nack_0_bits_uop_uses_stq          (io_dmem_nack_0_bits_uop_uses_stq),
  .io_dmem_resp_0_bits_is_hella              (io_dmem_resp_0_bits_is_hella),
  .send_iresp                                (send_iresp),
  .send_fresp                                (send_fresp),
  .io_dmem_nack_1_bits_uop_ldq_idx           (io_dmem_nack_1_bits_uop_ldq_idx),
  .io_dmem_nack_1_bits_uop_uses_stq          (io_dmem_nack_1_bits_uop_uses_stq),
  .io_dmem_resp_1_bits_is_hella              (io_dmem_resp_1_bits_is_hella),
  .send_iresp_1                              (send_iresp_1),
  .send_fresp_1                              (send_fresp_1),
  .stq_0_bits_committed                      (stq_0_bits_committed),
  ._GEN_262                                  (_GEN_1186),
  .stq_1_bits_committed                      (stq_1_bits_committed),
  ._GEN_263                                  (_GEN_1187),
  .stq_2_bits_committed                      (stq_2_bits_committed),
  ._GEN_264                                  (_GEN_1188),
  .stq_3_bits_committed                      (stq_3_bits_committed),
  ._GEN_265                                  (_GEN_1189),
  .stq_4_bits_committed                      (stq_4_bits_committed),
  ._GEN_266                                  (_GEN_1190),
  .stq_5_bits_committed                      (stq_5_bits_committed),
  ._GEN_267                                  (_GEN_1191),
  .stq_6_bits_committed                      (stq_6_bits_committed),
  ._GEN_268                                  (_GEN_1192),
  .stq_7_bits_committed                      (stq_7_bits_committed),
  ._GEN_269                                  (_GEN_1193),
  .stq_8_bits_committed                      (stq_8_bits_committed),
  ._GEN_270                                  (_GEN_1194),
  .stq_9_bits_committed                      (stq_9_bits_committed),
  ._GEN_271                                  (_GEN_1195),
  .stq_10_bits_committed                     (stq_10_bits_committed),
  ._GEN_272                                  (_GEN_1196),
  .stq_11_bits_committed                     (stq_11_bits_committed),
  ._GEN_273                                  (_GEN_1197),
  .stq_12_bits_committed                     (stq_12_bits_committed),
  ._GEN_274                                  (_GEN_1198),
  .stq_13_bits_committed                     (stq_13_bits_committed),
  ._GEN_275                                  (_GEN_1199),
  .stq_14_bits_committed                     (stq_14_bits_committed),
  ._GEN_276                                  (_GEN_1200),
  .stq_15_bits_committed                     (stq_15_bits_committed),
  ._GEN_277                                  (_GEN_1201),
  .stq_16_bits_committed                     (stq_16_bits_committed),
  ._GEN_278                                  (_GEN_1202),
  .stq_17_bits_committed                     (stq_17_bits_committed),
  ._GEN_279                                  (_GEN_1203),
  .stq_18_bits_committed                     (stq_18_bits_committed),
  ._GEN_280                                  (_GEN_1204),
  .stq_19_bits_committed                     (stq_19_bits_committed),
  ._GEN_281                                  (_GEN_1205),
  .stq_20_bits_committed                     (stq_20_bits_committed),
  ._GEN_282                                  (_GEN_1206),
  .stq_21_bits_committed                     (stq_21_bits_committed),
  ._GEN_283                                  (_GEN_1207),
  .stq_22_bits_committed                     (stq_22_bits_committed),
  ._GEN_284                                  (_GEN_1208),
  .stq_23_bits_committed                     (stq_23_bits_committed),
  ._GEN_285                                  (_GEN_1209),
  .stq_24_bits_committed                     (stq_24_bits_committed),
  ._GEN_286                                  (_GEN_1210),
  .stq_25_bits_committed                     (stq_25_bits_committed),
  ._GEN_287                                  (_GEN_1211),
  .stq_26_bits_committed                     (stq_26_bits_committed),
  ._GEN_288                                  (_GEN_1212),
  .stq_27_bits_committed                     (stq_27_bits_committed),
  ._GEN_289                                  (_GEN_1213),
  .stq_28_bits_committed                     (stq_28_bits_committed),
  ._GEN_290                                  (_GEN_1214),
  .stq_29_bits_committed                     (stq_29_bits_committed),
  ._GEN_291                                  (_GEN_1215),
  .stq_30_bits_committed                     (stq_30_bits_committed),
  ._GEN_292                                  (_GEN_1216),
  .stq_31_bits_committed                     (stq_31_bits_committed),
  ._GEN_293                                  (_GEN_1217),
  .idx                                       (idx),
  .ldq_31_bits_succeeded                     (ldq_31_bits_succeeded),
  .ldq_30_bits_succeeded                     (ldq_30_bits_succeeded),
  .ldq_29_bits_succeeded                     (ldq_29_bits_succeeded),
  .ldq_28_bits_succeeded                     (ldq_28_bits_succeeded),
  .ldq_27_bits_succeeded                     (ldq_27_bits_succeeded),
  .ldq_26_bits_succeeded                     (ldq_26_bits_succeeded),
  .ldq_25_bits_succeeded                     (ldq_25_bits_succeeded),
  .ldq_24_bits_succeeded                     (ldq_24_bits_succeeded),
  .ldq_23_bits_succeeded                     (ldq_23_bits_succeeded),
  .ldq_22_bits_succeeded                     (ldq_22_bits_succeeded),
  .ldq_21_bits_succeeded                     (ldq_21_bits_succeeded),
  .ldq_20_bits_succeeded                     (ldq_20_bits_succeeded),
  .ldq_19_bits_succeeded                     (ldq_19_bits_succeeded),
  .ldq_18_bits_succeeded                     (ldq_18_bits_succeeded),
  .ldq_17_bits_succeeded                     (ldq_17_bits_succeeded),
  .ldq_16_bits_succeeded                     (ldq_16_bits_succeeded),
  .ldq_15_bits_succeeded                     (ldq_15_bits_succeeded),
  .ldq_14_bits_succeeded                     (ldq_14_bits_succeeded),
  .ldq_13_bits_succeeded                     (ldq_13_bits_succeeded),
  .ldq_12_bits_succeeded                     (ldq_12_bits_succeeded),
  .ldq_11_bits_succeeded                     (ldq_11_bits_succeeded),
  .ldq_10_bits_succeeded                     (ldq_10_bits_succeeded),
  .ldq_9_bits_succeeded                      (ldq_9_bits_succeeded),
  .ldq_8_bits_succeeded                      (ldq_8_bits_succeeded),
  .ldq_7_bits_succeeded                      (ldq_7_bits_succeeded),
  .ldq_6_bits_succeeded                      (ldq_6_bits_succeeded),
  .ldq_5_bits_succeeded                      (ldq_5_bits_succeeded),
  .ldq_4_bits_succeeded                      (ldq_4_bits_succeeded),
  .ldq_3_bits_succeeded                      (ldq_3_bits_succeeded),
  .ldq_2_bits_succeeded                      (ldq_2_bits_succeeded),
  .ldq_1_bits_succeeded                      (ldq_1_bits_succeeded),
  .ldq_0_bits_succeeded                      (ldq_0_bits_succeeded),
  .ldq_31_bits_forward_std_val               (ldq_31_bits_forward_std_val),
  .ldq_30_bits_forward_std_val               (ldq_30_bits_forward_std_val),
  .ldq_29_bits_forward_std_val               (ldq_29_bits_forward_std_val),
  .ldq_28_bits_forward_std_val               (ldq_28_bits_forward_std_val),
  .ldq_27_bits_forward_std_val               (ldq_27_bits_forward_std_val),
  .ldq_26_bits_forward_std_val               (ldq_26_bits_forward_std_val),
  .ldq_25_bits_forward_std_val               (ldq_25_bits_forward_std_val),
  .ldq_24_bits_forward_std_val               (ldq_24_bits_forward_std_val),
  .ldq_23_bits_forward_std_val               (ldq_23_bits_forward_std_val),
  .ldq_22_bits_forward_std_val               (ldq_22_bits_forward_std_val),
  .ldq_21_bits_forward_std_val               (ldq_21_bits_forward_std_val),
  .ldq_20_bits_forward_std_val               (ldq_20_bits_forward_std_val),
  .ldq_19_bits_forward_std_val               (ldq_19_bits_forward_std_val),
  .ldq_18_bits_forward_std_val               (ldq_18_bits_forward_std_val),
  .ldq_17_bits_forward_std_val               (ldq_17_bits_forward_std_val),
  .ldq_16_bits_forward_std_val               (ldq_16_bits_forward_std_val),
  .ldq_15_bits_forward_std_val               (ldq_15_bits_forward_std_val),
  .ldq_14_bits_forward_std_val               (ldq_14_bits_forward_std_val),
  .ldq_13_bits_forward_std_val               (ldq_13_bits_forward_std_val),
  .ldq_12_bits_forward_std_val               (ldq_12_bits_forward_std_val),
  .ldq_11_bits_forward_std_val               (ldq_11_bits_forward_std_val),
  .ldq_10_bits_forward_std_val               (ldq_10_bits_forward_std_val),
  .ldq_9_bits_forward_std_val                (ldq_9_bits_forward_std_val),
  .ldq_8_bits_forward_std_val                (ldq_8_bits_forward_std_val),
  .ldq_7_bits_forward_std_val                (ldq_7_bits_forward_std_val),
  .ldq_6_bits_forward_std_val                (ldq_6_bits_forward_std_val),
  .ldq_5_bits_forward_std_val                (ldq_5_bits_forward_std_val),
  .ldq_4_bits_forward_std_val                (ldq_4_bits_forward_std_val),
  .ldq_3_bits_forward_std_val                (ldq_3_bits_forward_std_val),
  .ldq_2_bits_forward_std_val                (ldq_2_bits_forward_std_val),
  .ldq_1_bits_forward_std_val                (ldq_1_bits_forward_std_val),
  .ldq_0_bits_forward_std_val                (ldq_0_bits_forward_std_val),
  .idx_1                                     (idx_1),
  .idx_2                                     (idx_2),
  .idx_3                                     (idx_3),
  .reset                                     (reset),
  .mem_xcpt_valids_0                         (mem_xcpt_valids_0),
  .mem_xcpt_valids_1                         (mem_xcpt_valids_1),
  ._stq_idx_T                                (_stq_idx_T),
  ._GEN_294                                  (_GEN_335),
  .will_fire_load_wakeup_1                   (will_fire_load_wakeup_1),
  .will_fire_hella_incoming_1                (will_fire_hella_incoming_1),
  .will_fire_hella_wakeup_1                  (will_fire_hella_wakeup_1),
  ._GEN_295                                  (_GEN_341),
  ._GEN_296                                  (_GEN_342),
  ._stq_bits_data_bits_T_2                   (_stq_bits_data_bits_T_2),
  ._GEN_297                                  (_GEN_1230),
  .io_dmem_nack_0_bits_uop_uses_ldq          (io_dmem_nack_0_bits_uop_uses_ldq),
  .io_dmem_nack_0_valid                      (io_dmem_nack_0_valid),
  .io_dmem_nack_0_bits_is_hella              (io_dmem_nack_0_bits_is_hella),
  ._GEN_298                                  (_GEN_1178),
  .io_dmem_resp_0_valid                      (io_dmem_resp_0_valid),
  .io_dmem_resp_0_bits_uop_uses_stq          (io_dmem_resp_0_bits_uop_uses_stq),
  .io_dmem_resp_0_bits_uop_uses_ldq          (io_dmem_resp_0_bits_uop_uses_ldq),
  ._GEN_299                                  (_GEN_1232),
  .io_dmem_nack_1_bits_uop_uses_ldq          (io_dmem_nack_1_bits_uop_uses_ldq),
  .io_dmem_nack_1_valid                      (io_dmem_nack_1_valid),
  .io_dmem_nack_1_bits_is_hella              (io_dmem_nack_1_bits_is_hella),
  ._GEN_300                                  (_GEN_1182),
  .io_dmem_resp_1_valid                      (io_dmem_resp_1_valid),
  .io_dmem_resp_1_bits_uop_uses_stq          (io_dmem_resp_1_bits_uop_uses_stq),
  .io_dmem_resp_1_bits_uop_uses_ldq          (io_dmem_resp_1_bits_uop_uses_ldq),
  .commit_load                               (commit_load),
  .commit_store                              (commit_store),
  .commit_load_1                             (commit_load_1),
  .commit_store_1                            (commit_store_1),
  .commit_load_2                             (commit_load_2),
  .commit_store_2                            (commit_store_2),
  .commit_load_3                             (commit_load_3),
  .commit_store_3                            (commit_store_3)
);
bind PTW PTW_assert PTW_assert (
  .l2_hit                      (l2_hit),
  ._r_pte_T_2                  (_r_pte_T_2),
  .clock                       (clock),
  ._GEN                        (|state),
  ._GEN_0                      (_GEN_17),
  .pte_cache_hit               (pte_cache_hit),
  ._GEN_1                      (_GEN_19),
  ._resp_ae_ptw_T              (~(count[1])),
  ._GEN_2                      (_GEN_22),
  .s2_hit_vec_0                (s2_hit_vec_0),
  .l2_error                    (l2_error),
  ._s0_suitable_T_1            (~_arb_io_out_bits_bits_need_gpa),
  .arb_io_out_bits_bits_stage2 (_arb_io_out_bits_bits_stage2),
  ._GEN_3                      (_GEN_18),
  .state                       (state),
  .reset                       (reset),
  ._GEN_4                      (_GEN_21),
  ._GEN_5                      (_GEN_26),
  .mem_resp_valid              (mem_resp_valid),
  .io_mem_s2_nack              (io_mem_s2_nack)
);
bind TLBuffer_15 TLMonitor_42_assert TLMonitor_42_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_b_bits_opcode  (_nodeIn_b_q_io_deq_bits_opcode),
  .io_in_b_bits_address (_nodeIn_b_q_io_deq_bits_address),
  .io_in_b_bits_size    (_nodeIn_b_q_io_deq_bits_size),
  .io_in_b_bits_source  (_nodeIn_b_q_io_deq_bits_source),
  .io_in_b_bits_param   (_nodeIn_b_q_io_deq_bits_param),
  .io_in_b_bits_mask    (_nodeIn_b_q_io_deq_bits_mask),
  .io_in_b_bits_corrupt (_nodeIn_b_q_io_deq_bits_corrupt),
  .io_in_c_bits_address (auto_in_c_bits_address),
  .io_in_c_bits_source  (auto_in_c_bits_source),
  .io_in_c_bits_size    (auto_in_c_bits_size),
  .io_in_c_bits_param   (auto_in_c_bits_param),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink),
  .io_in_b_ready        (auto_in_b_ready),
  .io_in_b_valid        (_nodeIn_b_q_io_deq_valid),
  .io_in_c_bits_opcode  (auto_in_c_bits_opcode),
  .io_in_c_ready        (_nodeOut_c_q_io_enq_ready),
  .io_in_c_valid        (auto_in_c_valid),
  .io_in_e_bits_sink    (auto_in_e_bits_sink),
  .io_in_e_ready        (_nodeOut_e_q_io_enq_ready),
  .io_in_e_valid        (auto_in_e_valid)
);
bind TLPLIC TLMonitor_43_assert TLMonitor_43_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN_1),
  .io_in_d_bits_source  (_out_back_q_io_deq_bits_extra_tlrr_extra_source),
  .io_in_d_bits_size    (_out_back_q_io_deq_bits_extra_tlrr_extra_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_out_back_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_out_back_q_io_deq_valid)
);
bind TLPLIC TLPLIC_assert TLPLIC_assert (
  .claimer_1                   (claimer_1),
  .claimer_0                   (claimer_0),
  .completer_1                 (completer_1),
  .completer_0                 (completer_0),
  .completerDev                (_out_back_q_io_deq_bits_data[32]),
  .out_back_q_io_deq_bits_data (_out_back_q_io_deq_bits_data),
  .reset                       (reset),
  .clock                       (clock)
);
bind CLINT TLMonitor_44_assert TLMonitor_44_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN),
  .io_in_d_bits_source  (auto_in_a_bits_source),
  .io_in_d_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_in_d_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_in_a_valid)
);
bind TLXbar_10 TLMonitor_45_assert TLMonitor_45_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_d_bits_opcode  ((muxState_0 ? auto_out_0_d_bits_opcode : 3'h0) | (muxState_1 ? auto_out_1_d_bits_opcode : 3'h0)),
  .io_in_d_bits_size    ((muxState_0 ? auto_out_0_d_bits_size : 2'h0) | {muxState_1, 1'h0}),
  .io_in_d_bits_param   (muxState_0 ? auto_out_0_d_bits_param : 2'h0),
  .io_in_d_bits_corrupt (_in_0_d_bits_T),
  .io_in_d_bits_denied  (_in_0_d_bits_T_6),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (muxState_0 & auto_out_0_d_bits_sink)
);
bind TLXbar_10 TLXbar_10_assert TLXbar_10_assert (
  .winner_1        (winner_1),
  .winner_0        (winner_0),
  ._in_0_d_valid_T (_in_0_d_valid_T),
  .reset           (reset),
  .clock           (clock)
);
bind TLDebugModuleOuter TLMonitor_46_assert TLMonitor_46_assert (
  .io_in_a_bits_address (auto_dmi_in_a_bits_address),
  .io_in_d_bits_opcode  (_GEN),
  .io_in_a_bits_opcode  (auto_dmi_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_dmi_in_d_ready),
  .io_in_a_valid        (auto_dmi_in_a_valid),
  .io_in_d_ready        (auto_dmi_in_d_ready),
  .io_in_d_valid        (auto_dmi_in_a_valid)
);
bind TLBusBypassBar TLMonitor_47_assert TLMonitor_47_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_source  (~bypass & auto_out_1_d_bits_source),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_d_bits_param   (nodeIn_d_bits_param),
  .io_in_d_bits_corrupt (nodeIn_d_bits_corrupt),
  .io_in_d_bits_denied  (nodeIn_d_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid),
  .io_in_d_bits_sink    (nodeIn_d_bits_sink)
);
bind TLError_1 TLMonitor_48_assert TLMonitor_48_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_d_bits_param   (nodeIn_d_bits_param),
  .io_in_d_bits_corrupt (nodeIn_d_bits_corrupt),
  .io_in_d_bits_denied  (muxState_1),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLError_1 TLError_1_assert TLError_1_assert (
  .idle  (idle),
  .clock (clock),
  .reset (reset),
  .done  (done)
);
bind TLAsyncCrossingSource TLMonitor_49_assert TLMonitor_49_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_d_bits_opcode  (_nodeIn_d_sink_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_sink_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_sink_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_sink_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_sink_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_sink_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_source_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_sink_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_sink_io_deq_bits_sink)
);
bind TLDebugModuleInner TLMonitor_50_assert TLMonitor_50_assert (
  .io_in_a_bits_source  (auto_dmi_in_a_bits_source),
  .io_in_a_bits_size    (auto_dmi_in_a_bits_size),
  .io_in_a_bits_address (auto_dmi_in_a_bits_address),
  .io_in_a_bits_param   (auto_dmi_in_a_bits_param),
  .io_in_a_bits_mask    (auto_dmi_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_dmi_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN_3),
  .io_in_d_bits_source  (auto_dmi_in_a_bits_source),
  .io_in_d_bits_size    (auto_dmi_in_a_bits_size),
  .io_in_a_bits_opcode  (auto_dmi_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_dmi_in_d_ready),
  .io_in_a_valid        (auto_dmi_in_a_valid),
  .io_in_d_ready        (auto_dmi_in_d_ready),
  .io_in_d_valid        (auto_dmi_in_a_valid)
);
bind TLDebugModuleInner TLMonitor_51_assert TLMonitor_51_assert (
  .io_in_a_bits_source  (auto_tl_in_a_bits_source),
  .io_in_a_bits_size    (auto_tl_in_a_bits_size),
  .io_in_a_bits_address (auto_tl_in_a_bits_address),
  .io_in_a_bits_param   (auto_tl_in_a_bits_param),
  .io_in_a_bits_mask    (auto_tl_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_tl_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN_4),
  .io_in_d_bits_source  (auto_tl_in_a_bits_source),
  .io_in_d_bits_size    (auto_tl_in_a_bits_size),
  .io_in_a_bits_opcode  (auto_tl_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_tl_in_d_ready),
  .io_in_a_valid        (auto_tl_in_a_valid),
  .io_in_d_ready        (auto_tl_in_d_ready),
  .io_in_d_valid        (auto_tl_in_a_valid)
);
bind TLDebugModuleInner TLDebugModuleInner_assert TLDebugModuleInner_assert (
  .auto_tl_in_a_bits_data (auto_tl_in_a_bits_data),
  ._GEN                   (~io_dmactive),
  ._GEN_0                 (_GEN_2),
  .hartExceptionWrEn      (hartExceptionWrEn),
  .io_dmactive            (io_dmactive),
  .hartGoingWrEn          (hartGoingWrEn),
  .reset                  (reset),
  .goAbstract             (goAbstract),
  .clock                  (clock),
  ._errorBusy_T_14        (|ctrlStateReg),
  ._GEN_1                 (_GEN_0),
  .ctrlStateReg           (ctrlStateReg)
);
bind TLROM TLMonitor_52_assert TLMonitor_52_assert (
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_in_d_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (auto_in_a_valid),
  .io_in_d_bits_size    (auto_in_a_bits_size)
);
bind TLUART TLMonitor_53_assert TLMonitor_53_assert (
  .io_in_a_bits_source  (_buffer_auto_out_a_bits_source),
  .io_in_a_bits_size    (_buffer_auto_out_a_bits_size),
  .io_in_a_bits_address (_buffer_auto_out_a_bits_address),
  .io_in_a_bits_param   (_buffer_auto_out_a_bits_param),
  .io_in_a_bits_mask    (_buffer_auto_out_a_bits_mask),
  .io_in_a_bits_corrupt (_buffer_auto_out_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN),
  .io_in_d_bits_source  (_buffer_auto_out_a_bits_source),
  .io_in_d_bits_size    (_buffer_auto_out_a_bits_size),
  .io_in_a_bits_opcode  (_buffer_auto_out_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_buffer_auto_out_d_ready),
  .io_in_a_valid        (_buffer_auto_out_a_valid),
  .io_in_d_ready        (_buffer_auto_out_d_ready),
  .io_in_d_valid        (_buffer_auto_out_a_valid)
);
bind UARTTx UARTTx_assert UARTTx_assert (
  .io_in_bits (io_in_bits),
  ._GEN       (_GEN),
  .reset      (reset),
  .clock      (clock)
);
bind TLXbar_11 TLMonitor_54_assert TLMonitor_54_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (nodeIn_d_bits_opcode),
  .io_in_d_bits_source  (nodeIn_d_bits_source),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (nodeIn_a_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLXbar_11 TLXbar_11_assert TLXbar_11_assert (
  .winner_1        (winner_1),
  .winner_0        (winner_0),
  ._in_0_d_valid_T (_in_0_d_valid_T),
  .reset           (reset),
  .clock           (clock)
);
bind TileClockGater TLMonitor_55_assert TLMonitor_55_assert (
  .io_in_a_bits_source  (auto_clock_gater_in_1_a_bits_source),
  .io_in_a_bits_size    (auto_clock_gater_in_1_a_bits_size),
  .io_in_a_bits_address (auto_clock_gater_in_1_a_bits_address),
  .io_in_a_bits_param   (auto_clock_gater_in_1_a_bits_param),
  .io_in_a_bits_mask    (auto_clock_gater_in_1_a_bits_mask),
  .io_in_a_bits_corrupt (auto_clock_gater_in_1_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN),
  .io_in_d_bits_source  (auto_clock_gater_in_1_a_bits_source),
  .io_in_d_bits_size    (auto_clock_gater_in_1_a_bits_size),
  .io_in_a_bits_opcode  (auto_clock_gater_in_1_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_clock_gater_in_1_d_ready),
  .io_in_a_valid        (auto_clock_gater_in_1_a_valid),
  .io_in_d_ready        (auto_clock_gater_in_1_d_ready),
  .io_in_d_valid        (auto_clock_gater_in_1_a_valid)
);
bind TLFragmenter_7 TLMonitor_56_assert TLMonitor_56_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLFragmenter_7 TLFragmenter_7_assert TLFragmenter_7_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind TileResetSetter TLMonitor_57_assert TLMonitor_57_assert (
  .io_in_a_bits_source  (auto_tl_in_a_bits_source),
  .io_in_a_bits_size    (auto_tl_in_a_bits_size),
  .io_in_a_bits_address (auto_tl_in_a_bits_address),
  .io_in_a_bits_param   (auto_tl_in_a_bits_param),
  .io_in_a_bits_mask    (auto_tl_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_tl_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_GEN),
  .io_in_d_bits_source  (auto_tl_in_a_bits_source),
  .io_in_d_bits_size    (auto_tl_in_a_bits_size),
  .io_in_a_bits_opcode  (auto_tl_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (auto_tl_in_d_ready),
  .io_in_a_valid        (auto_tl_in_a_valid),
  .io_in_d_ready        (auto_tl_in_d_ready),
  .io_in_d_valid        (auto_tl_in_a_valid)
);
bind TLFragmenter_8 TLMonitor_58_assert TLMonitor_58_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_source  (auto_in_a_bits_source),
  .io_in_a_bits_param   (auto_in_a_bits_param),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (auto_out_d_bits_opcode),
  .io_in_d_bits_source  (auto_out_d_bits_source[10:4]),
  .io_in_d_bits_size    (nodeIn_d_bits_size),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_repeater_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (nodeIn_d_valid)
);
bind TLFragmenter_8 TLFragmenter_8_assert TLFragmenter_8_assert (
  ._repeater_io_repeat_T     (_repeater_io_deq_bits_opcode[2]),
  .repeater_io_full          (_repeater_io_full),
  .repeater_io_deq_bits_mask (_repeater_io_deq_bits_mask),
  .reset                     (reset),
  .clock                     (clock)
);
bind CaptureUpdateChain CaptureUpdateChain_assert CaptureUpdateChain_assert (
  .io_chainIn_update  (io_chainIn_update),
  .io_chainIn_shift   (io_chainIn_shift),
  .io_chainIn_capture (io_chainIn_capture),
  .reset              (reset),
  .clock              (clock)
);
bind CaptureUpdateChain_1 CaptureUpdateChain_1_assert CaptureUpdateChain_1_assert (
  .io_chainIn_update  (io_chainIn_update),
  .io_chainIn_shift   (io_chainIn_shift),
  .io_chainIn_capture (io_chainIn_capture),
  .reset              (reset),
  .clock              (clock)
);
bind CaptureChain CaptureChain_assert CaptureChain_assert (
  .io_chainIn_update  (io_chainIn_update),
  .io_chainIn_shift   (io_chainIn_shift),
  .io_chainIn_capture (io_chainIn_capture),
  .reset              (reset),
  .clock              (clock)
);
bind CaptureUpdateChain_2 CaptureUpdateChain_2_assert CaptureUpdateChain_2_assert (
  .io_chainIn_update  (io_chainIn_update),
  .io_chainIn_shift   (io_chainIn_shift),
  .io_chainIn_capture (io_chainIn_capture),
  .reset              (reset),
  .clock              (clock)
);
bind JtagBypassChain JtagBypassChain_assert JtagBypassChain_assert (
  .io_chainIn_update  (io_chainIn_update),
  .io_chainIn_shift   (io_chainIn_shift),
  .io_chainIn_capture (io_chainIn_capture),
  .reset              (reset),
  .clock              (clock)
);
bind DebugTransportModuleJTAG DebugTransportModuleJTAG_assert DebugTransportModuleJTAG_assert (
  .dmiAccessChain_io_update_valid (_dmiAccessChain_io_update_valid),
  ._GEN                           (_GEN_0),
  ._GEN_0                         (_GEN_1),
  .stickyBusyReg                  (stickyBusyReg),
  .io_jtag_reset                  (io_jtag_reset),
  .io_jtag_clock                  (io_jtag_clock)
);
bind TSIToTileLink TSIToTileLink_assert TSIToTileLink_assert (
  ._GEN   (_GEN_3),
  ._GEN_0 (|cmd),
  .reset  (reset),
  ._GEN_1 (_GEN_2),
  .clock  (clock)
);
bind TLSerdesser_1 TLMonitor_59_assert TLMonitor_59_assert (
  .io_in_a_bits_address (auto_manager_in_a_bits_address),
  .io_in_a_bits_size    (auto_manager_in_a_bits_size),
  .io_in_a_bits_source  (auto_manager_in_a_bits_source),
  .io_in_a_bits_param   (auto_manager_in_a_bits_param),
  .io_in_a_bits_mask    (auto_manager_in_a_bits_mask),
  .io_in_a_bits_corrupt (auto_manager_in_a_bits_corrupt),
  .io_in_d_bits_opcode  (_inDes_io_out_bits_opcode),
  .io_in_d_bits_source  (_inDes_io_out_bits_source[0]),
  .io_in_d_bits_size    (_inDes_io_out_bits_size[3:0]),
  .io_in_d_bits_param   (_inDes_io_out_bits_param[1:0]),
  .io_in_d_bits_corrupt (_inDes_io_out_bits_corrupt),
  .io_in_d_bits_denied  (_inDes_io_out_bits_union[0]),
  .io_in_a_bits_opcode  (auto_manager_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_outArb_io_in_4_ready),
  .io_in_a_valid        (auto_manager_in_a_valid),
  .io_in_d_ready        (auto_manager_in_d_ready),
  .io_in_d_valid        (managerNodeIn_d_valid),
  .io_in_d_bits_sink    (_inDes_io_out_bits_union[4:1])
);
bind TLBuffer_18 TLMonitor_60_assert TLMonitor_60_assert (
  .io_in_a_bits_address (auto_in_a_bits_address),
  .io_in_a_bits_size    (auto_in_a_bits_size),
  .io_in_a_bits_mask    (auto_in_a_bits_mask),
  .io_in_d_bits_opcode  (_nodeIn_d_q_io_deq_bits_opcode),
  .io_in_d_bits_source  (_nodeIn_d_q_io_deq_bits_source),
  .io_in_d_bits_size    (_nodeIn_d_q_io_deq_bits_size),
  .io_in_d_bits_param   (_nodeIn_d_q_io_deq_bits_param),
  .io_in_d_bits_corrupt (_nodeIn_d_q_io_deq_bits_corrupt),
  .io_in_d_bits_denied  (_nodeIn_d_q_io_deq_bits_denied),
  .io_in_a_bits_opcode  (auto_in_a_bits_opcode),
  .clock                (clock),
  .reset                (reset),
  .io_in_a_ready        (_nodeOut_a_q_io_enq_ready),
  .io_in_a_valid        (auto_in_a_valid),
  .io_in_d_ready        (auto_in_d_ready),
  .io_in_d_valid        (_nodeIn_d_q_io_deq_valid),
  .io_in_d_bits_sink    (_nodeIn_d_q_io_deq_bits_sink)
);
bind UARTAdapter UARTAdapter_assert UARTAdapter_assert (
  .txq_io_enq_ready (_txq_io_enq_ready),
  .txm_io_out_valid (_txm_io_out_valid),
  .reset            (reset),
  .clock            (clock)
);
bind TestHarness TestHarness_assert TestHarness_assert (
  .jtag_exit                                (_jtag_exit),
  .success_exit_sim_exit                    (_success_exit_sim_exit),
  ._GEN                                     (~_harnessBinderReset_catcher_io_sync_reset),
  .source_1_clk                             (_source_1_clk),
  .harnessBinderReset_catcher_io_sync_reset (_harnessBinderReset_catcher_io_sync_reset)
);
