// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

module Rob(
  input         clock,
                reset,
                io_enq_valids_0,
                io_enq_valids_1,
                io_enq_valids_2,
                io_enq_valids_3,
  input  [6:0]  io_enq_uops_0_uopc,
  input         io_enq_uops_0_is_rvc,
                io_enq_uops_0_is_br,
                io_enq_uops_0_is_jalr,
  input  [19:0] io_enq_uops_0_br_mask,
  input  [5:0]  io_enq_uops_0_ftq_idx,
  input         io_enq_uops_0_edge_inst,
  input  [5:0]  io_enq_uops_0_pc_lob,
  input  [6:0]  io_enq_uops_0_rob_idx,
                io_enq_uops_0_pdst,
                io_enq_uops_0_stale_pdst,
  input         io_enq_uops_0_exception,
  input  [63:0] io_enq_uops_0_exc_cause,
  input         io_enq_uops_0_is_fence,
                io_enq_uops_0_is_fencei,
                io_enq_uops_0_uses_ldq,
                io_enq_uops_0_uses_stq,
                io_enq_uops_0_is_sys_pc2epc,
                io_enq_uops_0_is_unique,
                io_enq_uops_0_flush_on_commit,
  input  [5:0]  io_enq_uops_0_ldst,
  input         io_enq_uops_0_ldst_val,
  input  [1:0]  io_enq_uops_0_dst_rtype,
  input         io_enq_uops_0_fp_val,
  input  [6:0]  io_enq_uops_1_uopc,
  input         io_enq_uops_1_is_rvc,
                io_enq_uops_1_is_br,
                io_enq_uops_1_is_jalr,
  input  [19:0] io_enq_uops_1_br_mask,
  input  [5:0]  io_enq_uops_1_ftq_idx,
  input         io_enq_uops_1_edge_inst,
  input  [5:0]  io_enq_uops_1_pc_lob,
  input  [6:0]  io_enq_uops_1_rob_idx,
                io_enq_uops_1_pdst,
                io_enq_uops_1_stale_pdst,
  input         io_enq_uops_1_exception,
  input  [63:0] io_enq_uops_1_exc_cause,
  input         io_enq_uops_1_is_fence,
                io_enq_uops_1_is_fencei,
                io_enq_uops_1_uses_ldq,
                io_enq_uops_1_uses_stq,
                io_enq_uops_1_is_sys_pc2epc,
                io_enq_uops_1_is_unique,
                io_enq_uops_1_flush_on_commit,
  input  [5:0]  io_enq_uops_1_ldst,
  input         io_enq_uops_1_ldst_val,
  input  [1:0]  io_enq_uops_1_dst_rtype,
  input         io_enq_uops_1_fp_val,
  input  [6:0]  io_enq_uops_2_uopc,
  input         io_enq_uops_2_is_rvc,
                io_enq_uops_2_is_br,
                io_enq_uops_2_is_jalr,
  input  [19:0] io_enq_uops_2_br_mask,
  input  [5:0]  io_enq_uops_2_ftq_idx,
  input         io_enq_uops_2_edge_inst,
  input  [5:0]  io_enq_uops_2_pc_lob,
  input  [6:0]  io_enq_uops_2_rob_idx,
                io_enq_uops_2_pdst,
                io_enq_uops_2_stale_pdst,
  input         io_enq_uops_2_exception,
  input  [63:0] io_enq_uops_2_exc_cause,
  input         io_enq_uops_2_is_fence,
                io_enq_uops_2_is_fencei,
                io_enq_uops_2_uses_ldq,
                io_enq_uops_2_uses_stq,
                io_enq_uops_2_is_sys_pc2epc,
                io_enq_uops_2_is_unique,
                io_enq_uops_2_flush_on_commit,
  input  [5:0]  io_enq_uops_2_ldst,
  input         io_enq_uops_2_ldst_val,
  input  [1:0]  io_enq_uops_2_dst_rtype,
  input         io_enq_uops_2_fp_val,
  input  [6:0]  io_enq_uops_3_uopc,
  input         io_enq_uops_3_is_rvc,
                io_enq_uops_3_is_br,
                io_enq_uops_3_is_jalr,
  input  [19:0] io_enq_uops_3_br_mask,
  input  [5:0]  io_enq_uops_3_ftq_idx,
  input         io_enq_uops_3_edge_inst,
  input  [5:0]  io_enq_uops_3_pc_lob,
  input  [6:0]  io_enq_uops_3_rob_idx,
                io_enq_uops_3_pdst,
                io_enq_uops_3_stale_pdst,
  input         io_enq_uops_3_exception,
  input  [63:0] io_enq_uops_3_exc_cause,
  input         io_enq_uops_3_is_fence,
                io_enq_uops_3_is_fencei,
                io_enq_uops_3_uses_ldq,
                io_enq_uops_3_uses_stq,
                io_enq_uops_3_is_sys_pc2epc,
                io_enq_uops_3_is_unique,
                io_enq_uops_3_flush_on_commit,
  input  [5:0]  io_enq_uops_3_ldst,
  input         io_enq_uops_3_ldst_val,
  input  [1:0]  io_enq_uops_3_dst_rtype,
  input         io_enq_uops_3_fp_val,
                io_enq_partial_stall,
  input  [39:0] io_xcpt_fetch_pc,
  input  [19:0] io_brupdate_b1_resolve_mask,
                io_brupdate_b1_mispredict_mask,
  input  [6:0]  io_brupdate_b2_uop_rob_idx,
  input         io_brupdate_b2_mispredict,
                io_wb_resps_0_valid,
  input  [6:0]  io_wb_resps_0_bits_uop_rob_idx,
                io_wb_resps_0_bits_uop_pdst,
  input         io_wb_resps_0_bits_predicated,
                io_wb_resps_1_valid,
  input  [6:0]  io_wb_resps_1_bits_uop_rob_idx,
                io_wb_resps_1_bits_uop_pdst,
  input         io_wb_resps_2_valid,
  input  [6:0]  io_wb_resps_2_bits_uop_rob_idx,
                io_wb_resps_2_bits_uop_pdst,
  input         io_wb_resps_3_valid,
  input  [6:0]  io_wb_resps_3_bits_uop_rob_idx,
                io_wb_resps_3_bits_uop_pdst,
  input         io_wb_resps_4_valid,
  input  [6:0]  io_wb_resps_4_bits_uop_rob_idx,
                io_wb_resps_4_bits_uop_pdst,
  input         io_wb_resps_5_valid,
  input  [6:0]  io_wb_resps_5_bits_uop_rob_idx,
                io_wb_resps_5_bits_uop_pdst,
  input         io_wb_resps_6_valid,
  input  [6:0]  io_wb_resps_6_bits_uop_rob_idx,
                io_wb_resps_6_bits_uop_pdst,
  input         io_wb_resps_6_bits_predicated,
                io_wb_resps_7_valid,
  input  [6:0]  io_wb_resps_7_bits_uop_rob_idx,
                io_wb_resps_7_bits_uop_pdst,
  input         io_wb_resps_8_valid,
  input  [6:0]  io_wb_resps_8_bits_uop_rob_idx,
                io_wb_resps_8_bits_uop_pdst,
  input         io_wb_resps_9_valid,
  input  [6:0]  io_wb_resps_9_bits_uop_rob_idx,
                io_wb_resps_9_bits_uop_pdst,
  input         io_lsu_clr_bsy_0_valid,
  input  [6:0]  io_lsu_clr_bsy_0_bits,
  input         io_lsu_clr_bsy_1_valid,
  input  [6:0]  io_lsu_clr_bsy_1_bits,
  input         io_lsu_clr_bsy_2_valid,
  input  [6:0]  io_lsu_clr_bsy_2_bits,
  input         io_fflags_0_valid,
  input  [6:0]  io_fflags_0_bits_uop_rob_idx,
  input  [4:0]  io_fflags_0_bits_flags,
  input         io_fflags_2_valid,
  input  [6:0]  io_fflags_2_bits_uop_rob_idx,
  input  [4:0]  io_fflags_2_bits_flags,
  input         io_fflags_3_valid,
  input  [6:0]  io_fflags_3_bits_uop_rob_idx,
  input  [4:0]  io_fflags_3_bits_flags,
  input         io_lxcpt_valid,
  input  [19:0] io_lxcpt_bits_uop_br_mask,
  input  [6:0]  io_lxcpt_bits_uop_rob_idx,
  input  [4:0]  io_lxcpt_bits_cause,
  input  [39:0] io_lxcpt_bits_badvaddr,
  input         io_csr_stall,
  output [6:0]  io_rob_tail_idx,
                io_rob_head_idx,
  output        io_commit_valids_0,
                io_commit_valids_1,
                io_commit_valids_2,
                io_commit_valids_3,
                io_commit_arch_valids_0,
                io_commit_arch_valids_1,
                io_commit_arch_valids_2,
                io_commit_arch_valids_3,
  output [5:0]  io_commit_uops_0_ftq_idx,
  output [6:0]  io_commit_uops_0_pdst,
                io_commit_uops_0_stale_pdst,
  output        io_commit_uops_0_is_fencei,
                io_commit_uops_0_uses_ldq,
                io_commit_uops_0_uses_stq,
  output [5:0]  io_commit_uops_0_ldst,
  output        io_commit_uops_0_ldst_val,
  output [1:0]  io_commit_uops_0_dst_rtype,
  output [5:0]  io_commit_uops_1_ftq_idx,
  output [6:0]  io_commit_uops_1_pdst,
                io_commit_uops_1_stale_pdst,
  output        io_commit_uops_1_is_fencei,
                io_commit_uops_1_uses_ldq,
                io_commit_uops_1_uses_stq,
  output [5:0]  io_commit_uops_1_ldst,
  output        io_commit_uops_1_ldst_val,
  output [1:0]  io_commit_uops_1_dst_rtype,
  output [5:0]  io_commit_uops_2_ftq_idx,
  output [6:0]  io_commit_uops_2_pdst,
                io_commit_uops_2_stale_pdst,
  output        io_commit_uops_2_is_fencei,
                io_commit_uops_2_uses_ldq,
                io_commit_uops_2_uses_stq,
  output [5:0]  io_commit_uops_2_ldst,
  output        io_commit_uops_2_ldst_val,
  output [1:0]  io_commit_uops_2_dst_rtype,
  output [5:0]  io_commit_uops_3_ftq_idx,
  output [6:0]  io_commit_uops_3_pdst,
                io_commit_uops_3_stale_pdst,
  output        io_commit_uops_3_is_fencei,
                io_commit_uops_3_uses_ldq,
                io_commit_uops_3_uses_stq,
  output [5:0]  io_commit_uops_3_ldst,
  output        io_commit_uops_3_ldst_val,
  output [1:0]  io_commit_uops_3_dst_rtype,
  output        io_commit_fflags_valid,
  output [4:0]  io_commit_fflags_bits,
  output        io_commit_rbk_valids_0,
                io_commit_rbk_valids_1,
                io_commit_rbk_valids_2,
                io_commit_rbk_valids_3,
                io_commit_rollback,
                io_com_load_is_at_rob_head,
                io_com_xcpt_valid,
  output [5:0]  io_com_xcpt_bits_ftq_idx,
  output        io_com_xcpt_bits_edge_inst,
  output [5:0]  io_com_xcpt_bits_pc_lob,
  output [63:0] io_com_xcpt_bits_cause,
                io_com_xcpt_bits_badvaddr,
  output        io_flush_valid,
  output [5:0]  io_flush_bits_ftq_idx,
  output        io_flush_bits_edge_inst,
                io_flush_bits_is_rvc,
  output [5:0]  io_flush_bits_pc_lob,
  output [2:0]  io_flush_bits_flush_typ,
  output        io_empty,
                io_ready,
                io_flush_frontend
);

  reg         casez_tmp;
  reg         casez_tmp_0;
  reg         casez_tmp_1;
  reg         casez_tmp_2;
  reg         casez_tmp_3;
  reg         casez_tmp_4;
  reg         casez_tmp_5;
  reg         casez_tmp_6;
  reg         casez_tmp_7;
  reg         casez_tmp_8;
  reg         casez_tmp_9;
  reg         casez_tmp_10;
  reg         casez_tmp_11;
  reg  [6:0]  casez_tmp_12;
  reg         casez_tmp_13;
  reg  [5:0]  casez_tmp_14;
  reg         casez_tmp_15;
  reg  [5:0]  casez_tmp_16;
  reg  [6:0]  casez_tmp_17;
  reg  [6:0]  casez_tmp_18;
  reg         casez_tmp_19;
  reg         casez_tmp_20;
  reg         casez_tmp_21;
  reg         casez_tmp_22;
  reg         casez_tmp_23;
  reg  [5:0]  casez_tmp_24;
  reg         casez_tmp_25;
  reg  [1:0]  casez_tmp_26;
  reg         casez_tmp_27;
  reg         casez_tmp_28;
  reg  [4:0]  casez_tmp_29;
  reg         casez_tmp_30;
  reg         casez_tmp_31;
  reg  [6:0]  casez_tmp_32;
  reg         casez_tmp_33;
  reg  [5:0]  casez_tmp_34;
  reg         casez_tmp_35;
  reg  [5:0]  casez_tmp_36;
  reg  [6:0]  casez_tmp_37;
  reg  [6:0]  casez_tmp_38;
  reg         casez_tmp_39;
  reg         casez_tmp_40;
  reg         casez_tmp_41;
  reg         casez_tmp_42;
  reg         casez_tmp_43;
  reg  [5:0]  casez_tmp_44;
  reg         casez_tmp_45;
  reg  [1:0]  casez_tmp_46;
  reg         casez_tmp_47;
  reg         casez_tmp_48;
  reg  [4:0]  casez_tmp_49;
  reg         casez_tmp_50;
  reg         casez_tmp_51;
  reg  [6:0]  casez_tmp_52;
  reg         casez_tmp_53;
  reg  [5:0]  casez_tmp_54;
  reg         casez_tmp_55;
  reg  [5:0]  casez_tmp_56;
  reg  [6:0]  casez_tmp_57;
  reg  [6:0]  casez_tmp_58;
  reg         casez_tmp_59;
  reg         casez_tmp_60;
  reg         casez_tmp_61;
  reg         casez_tmp_62;
  reg         casez_tmp_63;
  reg  [5:0]  casez_tmp_64;
  reg         casez_tmp_65;
  reg  [1:0]  casez_tmp_66;
  reg         casez_tmp_67;
  reg         casez_tmp_68;
  reg  [4:0]  casez_tmp_69;
  reg         casez_tmp_70;
  reg         casez_tmp_71;
  reg  [6:0]  casez_tmp_72;
  reg         casez_tmp_73;
  reg  [5:0]  casez_tmp_74;
  reg         casez_tmp_75;
  reg  [5:0]  casez_tmp_76;
  reg  [6:0]  casez_tmp_77;
  reg  [6:0]  casez_tmp_78;
  reg         casez_tmp_79;
  reg         casez_tmp_80;
  reg         casez_tmp_81;
  reg         casez_tmp_82;
  reg         casez_tmp_83;
  reg  [5:0]  casez_tmp_84;
  reg         casez_tmp_85;
  reg  [1:0]  casez_tmp_86;
  reg         casez_tmp_87;
  reg         casez_tmp_88;
  reg  [4:0]  casez_tmp_89;
  reg         casez_tmp_90;
  reg  [19:0] casez_tmp_91;
  reg  [5:0]  casez_tmp_92;
  reg  [6:0]  casez_tmp_93;
  reg  [63:0] casez_tmp_94;
  reg  [1:0]  casez_tmp_95;
  reg         casez_tmp_96;
  reg  [1:0]  rob_state;
  reg  [4:0]  rob_head;
  reg  [1:0]  rob_head_lsb;
  wire [6:0]  rob_head_idx = {rob_head, rob_head_lsb};
  reg  [4:0]  rob_tail;
  reg  [1:0]  rob_tail_lsb;
  wire [6:0]  rob_tail_idx = {rob_tail, rob_tail_lsb};
  wire        _io_commit_rollback_T_3 = rob_state == 2'h2;
  wire [4:0]  com_idx = _io_commit_rollback_T_3 ? rob_tail : rob_head;
  reg         maybe_full;
  reg         r_xcpt_val;
  reg  [19:0] r_xcpt_uop_br_mask;
  reg  [6:0]  r_xcpt_uop_rob_idx;
  reg  [63:0] r_xcpt_uop_exc_cause;
  reg  [39:0] r_xcpt_badvaddr;
  reg         rob_val__31;
  reg         rob_val__30;
  reg         rob_val__29;
  reg         rob_val__28;
  reg         rob_val__27;
  reg         rob_val__26;
  reg         rob_val__25;
  reg         rob_val__24;
  reg         rob_val__23;
  reg         rob_val__22;
  reg         rob_val__21;
  reg         rob_val__20;
  reg         rob_val__19;
  reg         rob_val__18;
  reg         rob_val__17;
  reg         rob_val__16;
  reg         rob_val__15;
  reg         rob_val__14;
  reg         rob_val__13;
  reg         rob_val__12;
  reg         rob_val__11;
  reg         rob_val__10;
  reg         rob_val__9;
  reg         rob_val__8;
  reg         rob_val__7;
  reg         rob_val__6;
  reg         rob_val__5;
  reg         rob_val__4;
  reg         rob_val__3;
  reg         rob_val__2;
  reg         rob_val__1;
  reg         rob_val__0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp = rob_val__0;
      5'b00001:
        casez_tmp = rob_val__1;
      5'b00010:
        casez_tmp = rob_val__2;
      5'b00011:
        casez_tmp = rob_val__3;
      5'b00100:
        casez_tmp = rob_val__4;
      5'b00101:
        casez_tmp = rob_val__5;
      5'b00110:
        casez_tmp = rob_val__6;
      5'b00111:
        casez_tmp = rob_val__7;
      5'b01000:
        casez_tmp = rob_val__8;
      5'b01001:
        casez_tmp = rob_val__9;
      5'b01010:
        casez_tmp = rob_val__10;
      5'b01011:
        casez_tmp = rob_val__11;
      5'b01100:
        casez_tmp = rob_val__12;
      5'b01101:
        casez_tmp = rob_val__13;
      5'b01110:
        casez_tmp = rob_val__14;
      5'b01111:
        casez_tmp = rob_val__15;
      5'b10000:
        casez_tmp = rob_val__16;
      5'b10001:
        casez_tmp = rob_val__17;
      5'b10010:
        casez_tmp = rob_val__18;
      5'b10011:
        casez_tmp = rob_val__19;
      5'b10100:
        casez_tmp = rob_val__20;
      5'b10101:
        casez_tmp = rob_val__21;
      5'b10110:
        casez_tmp = rob_val__22;
      5'b10111:
        casez_tmp = rob_val__23;
      5'b11000:
        casez_tmp = rob_val__24;
      5'b11001:
        casez_tmp = rob_val__25;
      5'b11010:
        casez_tmp = rob_val__26;
      5'b11011:
        casez_tmp = rob_val__27;
      5'b11100:
        casez_tmp = rob_val__28;
      5'b11101:
        casez_tmp = rob_val__29;
      5'b11110:
        casez_tmp = rob_val__30;
      default:
        casez_tmp = rob_val__31;
    endcase
  end // always @(*)
  reg         rob_bsy__31;
  reg         rob_bsy__30;
  reg         rob_bsy__29;
  reg         rob_bsy__28;
  reg         rob_bsy__27;
  reg         rob_bsy__26;
  reg         rob_bsy__25;
  reg         rob_bsy__24;
  reg         rob_bsy__23;
  reg         rob_bsy__22;
  reg         rob_bsy__21;
  reg         rob_bsy__20;
  reg         rob_bsy__19;
  reg         rob_bsy__18;
  reg         rob_bsy__17;
  reg         rob_bsy__16;
  reg         rob_bsy__15;
  reg         rob_bsy__14;
  reg         rob_bsy__13;
  reg         rob_bsy__12;
  reg         rob_bsy__11;
  reg         rob_bsy__10;
  reg         rob_bsy__9;
  reg         rob_bsy__8;
  reg         rob_bsy__7;
  reg         rob_bsy__6;
  reg         rob_bsy__5;
  reg         rob_bsy__4;
  reg         rob_bsy__3;
  reg         rob_bsy__2;
  reg         rob_bsy__1;
  reg         rob_bsy__0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_0 = rob_bsy__0;
      5'b00001:
        casez_tmp_0 = rob_bsy__1;
      5'b00010:
        casez_tmp_0 = rob_bsy__2;
      5'b00011:
        casez_tmp_0 = rob_bsy__3;
      5'b00100:
        casez_tmp_0 = rob_bsy__4;
      5'b00101:
        casez_tmp_0 = rob_bsy__5;
      5'b00110:
        casez_tmp_0 = rob_bsy__6;
      5'b00111:
        casez_tmp_0 = rob_bsy__7;
      5'b01000:
        casez_tmp_0 = rob_bsy__8;
      5'b01001:
        casez_tmp_0 = rob_bsy__9;
      5'b01010:
        casez_tmp_0 = rob_bsy__10;
      5'b01011:
        casez_tmp_0 = rob_bsy__11;
      5'b01100:
        casez_tmp_0 = rob_bsy__12;
      5'b01101:
        casez_tmp_0 = rob_bsy__13;
      5'b01110:
        casez_tmp_0 = rob_bsy__14;
      5'b01111:
        casez_tmp_0 = rob_bsy__15;
      5'b10000:
        casez_tmp_0 = rob_bsy__16;
      5'b10001:
        casez_tmp_0 = rob_bsy__17;
      5'b10010:
        casez_tmp_0 = rob_bsy__18;
      5'b10011:
        casez_tmp_0 = rob_bsy__19;
      5'b10100:
        casez_tmp_0 = rob_bsy__20;
      5'b10101:
        casez_tmp_0 = rob_bsy__21;
      5'b10110:
        casez_tmp_0 = rob_bsy__22;
      5'b10111:
        casez_tmp_0 = rob_bsy__23;
      5'b11000:
        casez_tmp_0 = rob_bsy__24;
      5'b11001:
        casez_tmp_0 = rob_bsy__25;
      5'b11010:
        casez_tmp_0 = rob_bsy__26;
      5'b11011:
        casez_tmp_0 = rob_bsy__27;
      5'b11100:
        casez_tmp_0 = rob_bsy__28;
      5'b11101:
        casez_tmp_0 = rob_bsy__29;
      5'b11110:
        casez_tmp_0 = rob_bsy__30;
      default:
        casez_tmp_0 = rob_bsy__31;
    endcase
  end // always @(*)
  wire        can_commit_0 = casez_tmp & ~casez_tmp_0 & ~io_csr_stall;
  reg         rob_exception__31;
  reg         rob_exception__30;
  reg         rob_exception__29;
  reg         rob_exception__28;
  reg         rob_exception__27;
  reg         rob_exception__26;
  reg         rob_exception__25;
  reg         rob_exception__24;
  reg         rob_exception__23;
  reg         rob_exception__22;
  reg         rob_exception__21;
  reg         rob_exception__20;
  reg         rob_exception__19;
  reg         rob_exception__18;
  reg         rob_exception__17;
  reg         rob_exception__16;
  reg         rob_exception__15;
  reg         rob_exception__14;
  reg         rob_exception__13;
  reg         rob_exception__12;
  reg         rob_exception__11;
  reg         rob_exception__10;
  reg         rob_exception__9;
  reg         rob_exception__8;
  reg         rob_exception__7;
  reg         rob_exception__6;
  reg         rob_exception__5;
  reg         rob_exception__4;
  reg         rob_exception__3;
  reg         rob_exception__2;
  reg         rob_exception__1;
  reg         rob_exception__0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_1 = rob_exception__0;
      5'b00001:
        casez_tmp_1 = rob_exception__1;
      5'b00010:
        casez_tmp_1 = rob_exception__2;
      5'b00011:
        casez_tmp_1 = rob_exception__3;
      5'b00100:
        casez_tmp_1 = rob_exception__4;
      5'b00101:
        casez_tmp_1 = rob_exception__5;
      5'b00110:
        casez_tmp_1 = rob_exception__6;
      5'b00111:
        casez_tmp_1 = rob_exception__7;
      5'b01000:
        casez_tmp_1 = rob_exception__8;
      5'b01001:
        casez_tmp_1 = rob_exception__9;
      5'b01010:
        casez_tmp_1 = rob_exception__10;
      5'b01011:
        casez_tmp_1 = rob_exception__11;
      5'b01100:
        casez_tmp_1 = rob_exception__12;
      5'b01101:
        casez_tmp_1 = rob_exception__13;
      5'b01110:
        casez_tmp_1 = rob_exception__14;
      5'b01111:
        casez_tmp_1 = rob_exception__15;
      5'b10000:
        casez_tmp_1 = rob_exception__16;
      5'b10001:
        casez_tmp_1 = rob_exception__17;
      5'b10010:
        casez_tmp_1 = rob_exception__18;
      5'b10011:
        casez_tmp_1 = rob_exception__19;
      5'b10100:
        casez_tmp_1 = rob_exception__20;
      5'b10101:
        casez_tmp_1 = rob_exception__21;
      5'b10110:
        casez_tmp_1 = rob_exception__22;
      5'b10111:
        casez_tmp_1 = rob_exception__23;
      5'b11000:
        casez_tmp_1 = rob_exception__24;
      5'b11001:
        casez_tmp_1 = rob_exception__25;
      5'b11010:
        casez_tmp_1 = rob_exception__26;
      5'b11011:
        casez_tmp_1 = rob_exception__27;
      5'b11100:
        casez_tmp_1 = rob_exception__28;
      5'b11101:
        casez_tmp_1 = rob_exception__29;
      5'b11110:
        casez_tmp_1 = rob_exception__30;
      default:
        casez_tmp_1 = rob_exception__31;
    endcase
  end // always @(*)
  wire        can_throw_exception_0 = casez_tmp & casez_tmp_1;
  reg         block_commit_REG;
  reg         block_commit_REG_2;
  wire        block_commit = rob_state != 2'h1 & rob_state != 2'h3 | block_commit_REG | block_commit_REG_2;
  wire        _io_commit_valids_0_output = can_commit_0 & ~can_throw_exception_0 & ~block_commit;
  reg         rob_val_1_31;
  reg         rob_val_1_30;
  reg         rob_val_1_29;
  reg         rob_val_1_28;
  reg         rob_val_1_27;
  reg         rob_val_1_26;
  reg         rob_val_1_25;
  reg         rob_val_1_24;
  reg         rob_val_1_23;
  reg         rob_val_1_22;
  reg         rob_val_1_21;
  reg         rob_val_1_20;
  reg         rob_val_1_19;
  reg         rob_val_1_18;
  reg         rob_val_1_17;
  reg         rob_val_1_16;
  reg         rob_val_1_15;
  reg         rob_val_1_14;
  reg         rob_val_1_13;
  reg         rob_val_1_12;
  reg         rob_val_1_11;
  reg         rob_val_1_10;
  reg         rob_val_1_9;
  reg         rob_val_1_8;
  reg         rob_val_1_7;
  reg         rob_val_1_6;
  reg         rob_val_1_5;
  reg         rob_val_1_4;
  reg         rob_val_1_3;
  reg         rob_val_1_2;
  reg         rob_val_1_1;
  reg         rob_val_1_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_2 = rob_val_1_0;
      5'b00001:
        casez_tmp_2 = rob_val_1_1;
      5'b00010:
        casez_tmp_2 = rob_val_1_2;
      5'b00011:
        casez_tmp_2 = rob_val_1_3;
      5'b00100:
        casez_tmp_2 = rob_val_1_4;
      5'b00101:
        casez_tmp_2 = rob_val_1_5;
      5'b00110:
        casez_tmp_2 = rob_val_1_6;
      5'b00111:
        casez_tmp_2 = rob_val_1_7;
      5'b01000:
        casez_tmp_2 = rob_val_1_8;
      5'b01001:
        casez_tmp_2 = rob_val_1_9;
      5'b01010:
        casez_tmp_2 = rob_val_1_10;
      5'b01011:
        casez_tmp_2 = rob_val_1_11;
      5'b01100:
        casez_tmp_2 = rob_val_1_12;
      5'b01101:
        casez_tmp_2 = rob_val_1_13;
      5'b01110:
        casez_tmp_2 = rob_val_1_14;
      5'b01111:
        casez_tmp_2 = rob_val_1_15;
      5'b10000:
        casez_tmp_2 = rob_val_1_16;
      5'b10001:
        casez_tmp_2 = rob_val_1_17;
      5'b10010:
        casez_tmp_2 = rob_val_1_18;
      5'b10011:
        casez_tmp_2 = rob_val_1_19;
      5'b10100:
        casez_tmp_2 = rob_val_1_20;
      5'b10101:
        casez_tmp_2 = rob_val_1_21;
      5'b10110:
        casez_tmp_2 = rob_val_1_22;
      5'b10111:
        casez_tmp_2 = rob_val_1_23;
      5'b11000:
        casez_tmp_2 = rob_val_1_24;
      5'b11001:
        casez_tmp_2 = rob_val_1_25;
      5'b11010:
        casez_tmp_2 = rob_val_1_26;
      5'b11011:
        casez_tmp_2 = rob_val_1_27;
      5'b11100:
        casez_tmp_2 = rob_val_1_28;
      5'b11101:
        casez_tmp_2 = rob_val_1_29;
      5'b11110:
        casez_tmp_2 = rob_val_1_30;
      default:
        casez_tmp_2 = rob_val_1_31;
    endcase
  end // always @(*)
  reg         rob_bsy_1_31;
  reg         rob_bsy_1_30;
  reg         rob_bsy_1_29;
  reg         rob_bsy_1_28;
  reg         rob_bsy_1_27;
  reg         rob_bsy_1_26;
  reg         rob_bsy_1_25;
  reg         rob_bsy_1_24;
  reg         rob_bsy_1_23;
  reg         rob_bsy_1_22;
  reg         rob_bsy_1_21;
  reg         rob_bsy_1_20;
  reg         rob_bsy_1_19;
  reg         rob_bsy_1_18;
  reg         rob_bsy_1_17;
  reg         rob_bsy_1_16;
  reg         rob_bsy_1_15;
  reg         rob_bsy_1_14;
  reg         rob_bsy_1_13;
  reg         rob_bsy_1_12;
  reg         rob_bsy_1_11;
  reg         rob_bsy_1_10;
  reg         rob_bsy_1_9;
  reg         rob_bsy_1_8;
  reg         rob_bsy_1_7;
  reg         rob_bsy_1_6;
  reg         rob_bsy_1_5;
  reg         rob_bsy_1_4;
  reg         rob_bsy_1_3;
  reg         rob_bsy_1_2;
  reg         rob_bsy_1_1;
  reg         rob_bsy_1_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_3 = rob_bsy_1_0;
      5'b00001:
        casez_tmp_3 = rob_bsy_1_1;
      5'b00010:
        casez_tmp_3 = rob_bsy_1_2;
      5'b00011:
        casez_tmp_3 = rob_bsy_1_3;
      5'b00100:
        casez_tmp_3 = rob_bsy_1_4;
      5'b00101:
        casez_tmp_3 = rob_bsy_1_5;
      5'b00110:
        casez_tmp_3 = rob_bsy_1_6;
      5'b00111:
        casez_tmp_3 = rob_bsy_1_7;
      5'b01000:
        casez_tmp_3 = rob_bsy_1_8;
      5'b01001:
        casez_tmp_3 = rob_bsy_1_9;
      5'b01010:
        casez_tmp_3 = rob_bsy_1_10;
      5'b01011:
        casez_tmp_3 = rob_bsy_1_11;
      5'b01100:
        casez_tmp_3 = rob_bsy_1_12;
      5'b01101:
        casez_tmp_3 = rob_bsy_1_13;
      5'b01110:
        casez_tmp_3 = rob_bsy_1_14;
      5'b01111:
        casez_tmp_3 = rob_bsy_1_15;
      5'b10000:
        casez_tmp_3 = rob_bsy_1_16;
      5'b10001:
        casez_tmp_3 = rob_bsy_1_17;
      5'b10010:
        casez_tmp_3 = rob_bsy_1_18;
      5'b10011:
        casez_tmp_3 = rob_bsy_1_19;
      5'b10100:
        casez_tmp_3 = rob_bsy_1_20;
      5'b10101:
        casez_tmp_3 = rob_bsy_1_21;
      5'b10110:
        casez_tmp_3 = rob_bsy_1_22;
      5'b10111:
        casez_tmp_3 = rob_bsy_1_23;
      5'b11000:
        casez_tmp_3 = rob_bsy_1_24;
      5'b11001:
        casez_tmp_3 = rob_bsy_1_25;
      5'b11010:
        casez_tmp_3 = rob_bsy_1_26;
      5'b11011:
        casez_tmp_3 = rob_bsy_1_27;
      5'b11100:
        casez_tmp_3 = rob_bsy_1_28;
      5'b11101:
        casez_tmp_3 = rob_bsy_1_29;
      5'b11110:
        casez_tmp_3 = rob_bsy_1_30;
      default:
        casez_tmp_3 = rob_bsy_1_31;
    endcase
  end // always @(*)
  wire        can_commit_1 = casez_tmp_2 & ~casez_tmp_3 & ~io_csr_stall;
  reg         rob_exception_1_31;
  reg         rob_exception_1_30;
  reg         rob_exception_1_29;
  reg         rob_exception_1_28;
  reg         rob_exception_1_27;
  reg         rob_exception_1_26;
  reg         rob_exception_1_25;
  reg         rob_exception_1_24;
  reg         rob_exception_1_23;
  reg         rob_exception_1_22;
  reg         rob_exception_1_21;
  reg         rob_exception_1_20;
  reg         rob_exception_1_19;
  reg         rob_exception_1_18;
  reg         rob_exception_1_17;
  reg         rob_exception_1_16;
  reg         rob_exception_1_15;
  reg         rob_exception_1_14;
  reg         rob_exception_1_13;
  reg         rob_exception_1_12;
  reg         rob_exception_1_11;
  reg         rob_exception_1_10;
  reg         rob_exception_1_9;
  reg         rob_exception_1_8;
  reg         rob_exception_1_7;
  reg         rob_exception_1_6;
  reg         rob_exception_1_5;
  reg         rob_exception_1_4;
  reg         rob_exception_1_3;
  reg         rob_exception_1_2;
  reg         rob_exception_1_1;
  reg         rob_exception_1_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_4 = rob_exception_1_0;
      5'b00001:
        casez_tmp_4 = rob_exception_1_1;
      5'b00010:
        casez_tmp_4 = rob_exception_1_2;
      5'b00011:
        casez_tmp_4 = rob_exception_1_3;
      5'b00100:
        casez_tmp_4 = rob_exception_1_4;
      5'b00101:
        casez_tmp_4 = rob_exception_1_5;
      5'b00110:
        casez_tmp_4 = rob_exception_1_6;
      5'b00111:
        casez_tmp_4 = rob_exception_1_7;
      5'b01000:
        casez_tmp_4 = rob_exception_1_8;
      5'b01001:
        casez_tmp_4 = rob_exception_1_9;
      5'b01010:
        casez_tmp_4 = rob_exception_1_10;
      5'b01011:
        casez_tmp_4 = rob_exception_1_11;
      5'b01100:
        casez_tmp_4 = rob_exception_1_12;
      5'b01101:
        casez_tmp_4 = rob_exception_1_13;
      5'b01110:
        casez_tmp_4 = rob_exception_1_14;
      5'b01111:
        casez_tmp_4 = rob_exception_1_15;
      5'b10000:
        casez_tmp_4 = rob_exception_1_16;
      5'b10001:
        casez_tmp_4 = rob_exception_1_17;
      5'b10010:
        casez_tmp_4 = rob_exception_1_18;
      5'b10011:
        casez_tmp_4 = rob_exception_1_19;
      5'b10100:
        casez_tmp_4 = rob_exception_1_20;
      5'b10101:
        casez_tmp_4 = rob_exception_1_21;
      5'b10110:
        casez_tmp_4 = rob_exception_1_22;
      5'b10111:
        casez_tmp_4 = rob_exception_1_23;
      5'b11000:
        casez_tmp_4 = rob_exception_1_24;
      5'b11001:
        casez_tmp_4 = rob_exception_1_25;
      5'b11010:
        casez_tmp_4 = rob_exception_1_26;
      5'b11011:
        casez_tmp_4 = rob_exception_1_27;
      5'b11100:
        casez_tmp_4 = rob_exception_1_28;
      5'b11101:
        casez_tmp_4 = rob_exception_1_29;
      5'b11110:
        casez_tmp_4 = rob_exception_1_30;
      default:
        casez_tmp_4 = rob_exception_1_31;
    endcase
  end // always @(*)
  wire        can_throw_exception_1 = casez_tmp_2 & casez_tmp_4;
  wire        _GEN = casez_tmp & (~can_commit_0 | can_throw_exception_0) | block_commit;
  wire        _io_commit_valids_1_output = can_commit_1 & ~can_throw_exception_1 & ~_GEN;
  reg         rob_val_2_31;
  reg         rob_val_2_30;
  reg         rob_val_2_29;
  reg         rob_val_2_28;
  reg         rob_val_2_27;
  reg         rob_val_2_26;
  reg         rob_val_2_25;
  reg         rob_val_2_24;
  reg         rob_val_2_23;
  reg         rob_val_2_22;
  reg         rob_val_2_21;
  reg         rob_val_2_20;
  reg         rob_val_2_19;
  reg         rob_val_2_18;
  reg         rob_val_2_17;
  reg         rob_val_2_16;
  reg         rob_val_2_15;
  reg         rob_val_2_14;
  reg         rob_val_2_13;
  reg         rob_val_2_12;
  reg         rob_val_2_11;
  reg         rob_val_2_10;
  reg         rob_val_2_9;
  reg         rob_val_2_8;
  reg         rob_val_2_7;
  reg         rob_val_2_6;
  reg         rob_val_2_5;
  reg         rob_val_2_4;
  reg         rob_val_2_3;
  reg         rob_val_2_2;
  reg         rob_val_2_1;
  reg         rob_val_2_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_5 = rob_val_2_0;
      5'b00001:
        casez_tmp_5 = rob_val_2_1;
      5'b00010:
        casez_tmp_5 = rob_val_2_2;
      5'b00011:
        casez_tmp_5 = rob_val_2_3;
      5'b00100:
        casez_tmp_5 = rob_val_2_4;
      5'b00101:
        casez_tmp_5 = rob_val_2_5;
      5'b00110:
        casez_tmp_5 = rob_val_2_6;
      5'b00111:
        casez_tmp_5 = rob_val_2_7;
      5'b01000:
        casez_tmp_5 = rob_val_2_8;
      5'b01001:
        casez_tmp_5 = rob_val_2_9;
      5'b01010:
        casez_tmp_5 = rob_val_2_10;
      5'b01011:
        casez_tmp_5 = rob_val_2_11;
      5'b01100:
        casez_tmp_5 = rob_val_2_12;
      5'b01101:
        casez_tmp_5 = rob_val_2_13;
      5'b01110:
        casez_tmp_5 = rob_val_2_14;
      5'b01111:
        casez_tmp_5 = rob_val_2_15;
      5'b10000:
        casez_tmp_5 = rob_val_2_16;
      5'b10001:
        casez_tmp_5 = rob_val_2_17;
      5'b10010:
        casez_tmp_5 = rob_val_2_18;
      5'b10011:
        casez_tmp_5 = rob_val_2_19;
      5'b10100:
        casez_tmp_5 = rob_val_2_20;
      5'b10101:
        casez_tmp_5 = rob_val_2_21;
      5'b10110:
        casez_tmp_5 = rob_val_2_22;
      5'b10111:
        casez_tmp_5 = rob_val_2_23;
      5'b11000:
        casez_tmp_5 = rob_val_2_24;
      5'b11001:
        casez_tmp_5 = rob_val_2_25;
      5'b11010:
        casez_tmp_5 = rob_val_2_26;
      5'b11011:
        casez_tmp_5 = rob_val_2_27;
      5'b11100:
        casez_tmp_5 = rob_val_2_28;
      5'b11101:
        casez_tmp_5 = rob_val_2_29;
      5'b11110:
        casez_tmp_5 = rob_val_2_30;
      default:
        casez_tmp_5 = rob_val_2_31;
    endcase
  end // always @(*)
  reg         rob_bsy_2_31;
  reg         rob_bsy_2_30;
  reg         rob_bsy_2_29;
  reg         rob_bsy_2_28;
  reg         rob_bsy_2_27;
  reg         rob_bsy_2_26;
  reg         rob_bsy_2_25;
  reg         rob_bsy_2_24;
  reg         rob_bsy_2_23;
  reg         rob_bsy_2_22;
  reg         rob_bsy_2_21;
  reg         rob_bsy_2_20;
  reg         rob_bsy_2_19;
  reg         rob_bsy_2_18;
  reg         rob_bsy_2_17;
  reg         rob_bsy_2_16;
  reg         rob_bsy_2_15;
  reg         rob_bsy_2_14;
  reg         rob_bsy_2_13;
  reg         rob_bsy_2_12;
  reg         rob_bsy_2_11;
  reg         rob_bsy_2_10;
  reg         rob_bsy_2_9;
  reg         rob_bsy_2_8;
  reg         rob_bsy_2_7;
  reg         rob_bsy_2_6;
  reg         rob_bsy_2_5;
  reg         rob_bsy_2_4;
  reg         rob_bsy_2_3;
  reg         rob_bsy_2_2;
  reg         rob_bsy_2_1;
  reg         rob_bsy_2_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_6 = rob_bsy_2_0;
      5'b00001:
        casez_tmp_6 = rob_bsy_2_1;
      5'b00010:
        casez_tmp_6 = rob_bsy_2_2;
      5'b00011:
        casez_tmp_6 = rob_bsy_2_3;
      5'b00100:
        casez_tmp_6 = rob_bsy_2_4;
      5'b00101:
        casez_tmp_6 = rob_bsy_2_5;
      5'b00110:
        casez_tmp_6 = rob_bsy_2_6;
      5'b00111:
        casez_tmp_6 = rob_bsy_2_7;
      5'b01000:
        casez_tmp_6 = rob_bsy_2_8;
      5'b01001:
        casez_tmp_6 = rob_bsy_2_9;
      5'b01010:
        casez_tmp_6 = rob_bsy_2_10;
      5'b01011:
        casez_tmp_6 = rob_bsy_2_11;
      5'b01100:
        casez_tmp_6 = rob_bsy_2_12;
      5'b01101:
        casez_tmp_6 = rob_bsy_2_13;
      5'b01110:
        casez_tmp_6 = rob_bsy_2_14;
      5'b01111:
        casez_tmp_6 = rob_bsy_2_15;
      5'b10000:
        casez_tmp_6 = rob_bsy_2_16;
      5'b10001:
        casez_tmp_6 = rob_bsy_2_17;
      5'b10010:
        casez_tmp_6 = rob_bsy_2_18;
      5'b10011:
        casez_tmp_6 = rob_bsy_2_19;
      5'b10100:
        casez_tmp_6 = rob_bsy_2_20;
      5'b10101:
        casez_tmp_6 = rob_bsy_2_21;
      5'b10110:
        casez_tmp_6 = rob_bsy_2_22;
      5'b10111:
        casez_tmp_6 = rob_bsy_2_23;
      5'b11000:
        casez_tmp_6 = rob_bsy_2_24;
      5'b11001:
        casez_tmp_6 = rob_bsy_2_25;
      5'b11010:
        casez_tmp_6 = rob_bsy_2_26;
      5'b11011:
        casez_tmp_6 = rob_bsy_2_27;
      5'b11100:
        casez_tmp_6 = rob_bsy_2_28;
      5'b11101:
        casez_tmp_6 = rob_bsy_2_29;
      5'b11110:
        casez_tmp_6 = rob_bsy_2_30;
      default:
        casez_tmp_6 = rob_bsy_2_31;
    endcase
  end // always @(*)
  wire        can_commit_2 = casez_tmp_5 & ~casez_tmp_6 & ~io_csr_stall;
  reg         rob_exception_2_31;
  reg         rob_exception_2_30;
  reg         rob_exception_2_29;
  reg         rob_exception_2_28;
  reg         rob_exception_2_27;
  reg         rob_exception_2_26;
  reg         rob_exception_2_25;
  reg         rob_exception_2_24;
  reg         rob_exception_2_23;
  reg         rob_exception_2_22;
  reg         rob_exception_2_21;
  reg         rob_exception_2_20;
  reg         rob_exception_2_19;
  reg         rob_exception_2_18;
  reg         rob_exception_2_17;
  reg         rob_exception_2_16;
  reg         rob_exception_2_15;
  reg         rob_exception_2_14;
  reg         rob_exception_2_13;
  reg         rob_exception_2_12;
  reg         rob_exception_2_11;
  reg         rob_exception_2_10;
  reg         rob_exception_2_9;
  reg         rob_exception_2_8;
  reg         rob_exception_2_7;
  reg         rob_exception_2_6;
  reg         rob_exception_2_5;
  reg         rob_exception_2_4;
  reg         rob_exception_2_3;
  reg         rob_exception_2_2;
  reg         rob_exception_2_1;
  reg         rob_exception_2_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_7 = rob_exception_2_0;
      5'b00001:
        casez_tmp_7 = rob_exception_2_1;
      5'b00010:
        casez_tmp_7 = rob_exception_2_2;
      5'b00011:
        casez_tmp_7 = rob_exception_2_3;
      5'b00100:
        casez_tmp_7 = rob_exception_2_4;
      5'b00101:
        casez_tmp_7 = rob_exception_2_5;
      5'b00110:
        casez_tmp_7 = rob_exception_2_6;
      5'b00111:
        casez_tmp_7 = rob_exception_2_7;
      5'b01000:
        casez_tmp_7 = rob_exception_2_8;
      5'b01001:
        casez_tmp_7 = rob_exception_2_9;
      5'b01010:
        casez_tmp_7 = rob_exception_2_10;
      5'b01011:
        casez_tmp_7 = rob_exception_2_11;
      5'b01100:
        casez_tmp_7 = rob_exception_2_12;
      5'b01101:
        casez_tmp_7 = rob_exception_2_13;
      5'b01110:
        casez_tmp_7 = rob_exception_2_14;
      5'b01111:
        casez_tmp_7 = rob_exception_2_15;
      5'b10000:
        casez_tmp_7 = rob_exception_2_16;
      5'b10001:
        casez_tmp_7 = rob_exception_2_17;
      5'b10010:
        casez_tmp_7 = rob_exception_2_18;
      5'b10011:
        casez_tmp_7 = rob_exception_2_19;
      5'b10100:
        casez_tmp_7 = rob_exception_2_20;
      5'b10101:
        casez_tmp_7 = rob_exception_2_21;
      5'b10110:
        casez_tmp_7 = rob_exception_2_22;
      5'b10111:
        casez_tmp_7 = rob_exception_2_23;
      5'b11000:
        casez_tmp_7 = rob_exception_2_24;
      5'b11001:
        casez_tmp_7 = rob_exception_2_25;
      5'b11010:
        casez_tmp_7 = rob_exception_2_26;
      5'b11011:
        casez_tmp_7 = rob_exception_2_27;
      5'b11100:
        casez_tmp_7 = rob_exception_2_28;
      5'b11101:
        casez_tmp_7 = rob_exception_2_29;
      5'b11110:
        casez_tmp_7 = rob_exception_2_30;
      default:
        casez_tmp_7 = rob_exception_2_31;
    endcase
  end // always @(*)
  wire        can_throw_exception_2 = casez_tmp_5 & casez_tmp_7;
  wire        _GEN_0 = casez_tmp_2 & (~can_commit_1 | can_throw_exception_1) | _GEN;
  wire        _io_commit_valids_2_output = can_commit_2 & ~can_throw_exception_2 & ~_GEN_0;
  reg         rob_val_3_31;
  reg         rob_val_3_30;
  reg         rob_val_3_29;
  reg         rob_val_3_28;
  reg         rob_val_3_27;
  reg         rob_val_3_26;
  reg         rob_val_3_25;
  reg         rob_val_3_24;
  reg         rob_val_3_23;
  reg         rob_val_3_22;
  reg         rob_val_3_21;
  reg         rob_val_3_20;
  reg         rob_val_3_19;
  reg         rob_val_3_18;
  reg         rob_val_3_17;
  reg         rob_val_3_16;
  reg         rob_val_3_15;
  reg         rob_val_3_14;
  reg         rob_val_3_13;
  reg         rob_val_3_12;
  reg         rob_val_3_11;
  reg         rob_val_3_10;
  reg         rob_val_3_9;
  reg         rob_val_3_8;
  reg         rob_val_3_7;
  reg         rob_val_3_6;
  reg         rob_val_3_5;
  reg         rob_val_3_4;
  reg         rob_val_3_3;
  reg         rob_val_3_2;
  reg         rob_val_3_1;
  reg         rob_val_3_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_8 = rob_val_3_0;
      5'b00001:
        casez_tmp_8 = rob_val_3_1;
      5'b00010:
        casez_tmp_8 = rob_val_3_2;
      5'b00011:
        casez_tmp_8 = rob_val_3_3;
      5'b00100:
        casez_tmp_8 = rob_val_3_4;
      5'b00101:
        casez_tmp_8 = rob_val_3_5;
      5'b00110:
        casez_tmp_8 = rob_val_3_6;
      5'b00111:
        casez_tmp_8 = rob_val_3_7;
      5'b01000:
        casez_tmp_8 = rob_val_3_8;
      5'b01001:
        casez_tmp_8 = rob_val_3_9;
      5'b01010:
        casez_tmp_8 = rob_val_3_10;
      5'b01011:
        casez_tmp_8 = rob_val_3_11;
      5'b01100:
        casez_tmp_8 = rob_val_3_12;
      5'b01101:
        casez_tmp_8 = rob_val_3_13;
      5'b01110:
        casez_tmp_8 = rob_val_3_14;
      5'b01111:
        casez_tmp_8 = rob_val_3_15;
      5'b10000:
        casez_tmp_8 = rob_val_3_16;
      5'b10001:
        casez_tmp_8 = rob_val_3_17;
      5'b10010:
        casez_tmp_8 = rob_val_3_18;
      5'b10011:
        casez_tmp_8 = rob_val_3_19;
      5'b10100:
        casez_tmp_8 = rob_val_3_20;
      5'b10101:
        casez_tmp_8 = rob_val_3_21;
      5'b10110:
        casez_tmp_8 = rob_val_3_22;
      5'b10111:
        casez_tmp_8 = rob_val_3_23;
      5'b11000:
        casez_tmp_8 = rob_val_3_24;
      5'b11001:
        casez_tmp_8 = rob_val_3_25;
      5'b11010:
        casez_tmp_8 = rob_val_3_26;
      5'b11011:
        casez_tmp_8 = rob_val_3_27;
      5'b11100:
        casez_tmp_8 = rob_val_3_28;
      5'b11101:
        casez_tmp_8 = rob_val_3_29;
      5'b11110:
        casez_tmp_8 = rob_val_3_30;
      default:
        casez_tmp_8 = rob_val_3_31;
    endcase
  end // always @(*)
  reg         rob_bsy_3_31;
  reg         rob_bsy_3_30;
  reg         rob_bsy_3_29;
  reg         rob_bsy_3_28;
  reg         rob_bsy_3_27;
  reg         rob_bsy_3_26;
  reg         rob_bsy_3_25;
  reg         rob_bsy_3_24;
  reg         rob_bsy_3_23;
  reg         rob_bsy_3_22;
  reg         rob_bsy_3_21;
  reg         rob_bsy_3_20;
  reg         rob_bsy_3_19;
  reg         rob_bsy_3_18;
  reg         rob_bsy_3_17;
  reg         rob_bsy_3_16;
  reg         rob_bsy_3_15;
  reg         rob_bsy_3_14;
  reg         rob_bsy_3_13;
  reg         rob_bsy_3_12;
  reg         rob_bsy_3_11;
  reg         rob_bsy_3_10;
  reg         rob_bsy_3_9;
  reg         rob_bsy_3_8;
  reg         rob_bsy_3_7;
  reg         rob_bsy_3_6;
  reg         rob_bsy_3_5;
  reg         rob_bsy_3_4;
  reg         rob_bsy_3_3;
  reg         rob_bsy_3_2;
  reg         rob_bsy_3_1;
  reg         rob_bsy_3_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_9 = rob_bsy_3_0;
      5'b00001:
        casez_tmp_9 = rob_bsy_3_1;
      5'b00010:
        casez_tmp_9 = rob_bsy_3_2;
      5'b00011:
        casez_tmp_9 = rob_bsy_3_3;
      5'b00100:
        casez_tmp_9 = rob_bsy_3_4;
      5'b00101:
        casez_tmp_9 = rob_bsy_3_5;
      5'b00110:
        casez_tmp_9 = rob_bsy_3_6;
      5'b00111:
        casez_tmp_9 = rob_bsy_3_7;
      5'b01000:
        casez_tmp_9 = rob_bsy_3_8;
      5'b01001:
        casez_tmp_9 = rob_bsy_3_9;
      5'b01010:
        casez_tmp_9 = rob_bsy_3_10;
      5'b01011:
        casez_tmp_9 = rob_bsy_3_11;
      5'b01100:
        casez_tmp_9 = rob_bsy_3_12;
      5'b01101:
        casez_tmp_9 = rob_bsy_3_13;
      5'b01110:
        casez_tmp_9 = rob_bsy_3_14;
      5'b01111:
        casez_tmp_9 = rob_bsy_3_15;
      5'b10000:
        casez_tmp_9 = rob_bsy_3_16;
      5'b10001:
        casez_tmp_9 = rob_bsy_3_17;
      5'b10010:
        casez_tmp_9 = rob_bsy_3_18;
      5'b10011:
        casez_tmp_9 = rob_bsy_3_19;
      5'b10100:
        casez_tmp_9 = rob_bsy_3_20;
      5'b10101:
        casez_tmp_9 = rob_bsy_3_21;
      5'b10110:
        casez_tmp_9 = rob_bsy_3_22;
      5'b10111:
        casez_tmp_9 = rob_bsy_3_23;
      5'b11000:
        casez_tmp_9 = rob_bsy_3_24;
      5'b11001:
        casez_tmp_9 = rob_bsy_3_25;
      5'b11010:
        casez_tmp_9 = rob_bsy_3_26;
      5'b11011:
        casez_tmp_9 = rob_bsy_3_27;
      5'b11100:
        casez_tmp_9 = rob_bsy_3_28;
      5'b11101:
        casez_tmp_9 = rob_bsy_3_29;
      5'b11110:
        casez_tmp_9 = rob_bsy_3_30;
      default:
        casez_tmp_9 = rob_bsy_3_31;
    endcase
  end // always @(*)
  reg         rob_exception_3_31;
  reg         rob_exception_3_30;
  reg         rob_exception_3_29;
  reg         rob_exception_3_28;
  reg         rob_exception_3_27;
  reg         rob_exception_3_26;
  reg         rob_exception_3_25;
  reg         rob_exception_3_24;
  reg         rob_exception_3_23;
  reg         rob_exception_3_22;
  reg         rob_exception_3_21;
  reg         rob_exception_3_20;
  reg         rob_exception_3_19;
  reg         rob_exception_3_18;
  reg         rob_exception_3_17;
  reg         rob_exception_3_16;
  reg         rob_exception_3_15;
  reg         rob_exception_3_14;
  reg         rob_exception_3_13;
  reg         rob_exception_3_12;
  reg         rob_exception_3_11;
  reg         rob_exception_3_10;
  reg         rob_exception_3_9;
  reg         rob_exception_3_8;
  reg         rob_exception_3_7;
  reg         rob_exception_3_6;
  reg         rob_exception_3_5;
  reg         rob_exception_3_4;
  reg         rob_exception_3_3;
  reg         rob_exception_3_2;
  reg         rob_exception_3_1;
  reg         rob_exception_3_0;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_10 = rob_exception_3_0;
      5'b00001:
        casez_tmp_10 = rob_exception_3_1;
      5'b00010:
        casez_tmp_10 = rob_exception_3_2;
      5'b00011:
        casez_tmp_10 = rob_exception_3_3;
      5'b00100:
        casez_tmp_10 = rob_exception_3_4;
      5'b00101:
        casez_tmp_10 = rob_exception_3_5;
      5'b00110:
        casez_tmp_10 = rob_exception_3_6;
      5'b00111:
        casez_tmp_10 = rob_exception_3_7;
      5'b01000:
        casez_tmp_10 = rob_exception_3_8;
      5'b01001:
        casez_tmp_10 = rob_exception_3_9;
      5'b01010:
        casez_tmp_10 = rob_exception_3_10;
      5'b01011:
        casez_tmp_10 = rob_exception_3_11;
      5'b01100:
        casez_tmp_10 = rob_exception_3_12;
      5'b01101:
        casez_tmp_10 = rob_exception_3_13;
      5'b01110:
        casez_tmp_10 = rob_exception_3_14;
      5'b01111:
        casez_tmp_10 = rob_exception_3_15;
      5'b10000:
        casez_tmp_10 = rob_exception_3_16;
      5'b10001:
        casez_tmp_10 = rob_exception_3_17;
      5'b10010:
        casez_tmp_10 = rob_exception_3_18;
      5'b10011:
        casez_tmp_10 = rob_exception_3_19;
      5'b10100:
        casez_tmp_10 = rob_exception_3_20;
      5'b10101:
        casez_tmp_10 = rob_exception_3_21;
      5'b10110:
        casez_tmp_10 = rob_exception_3_22;
      5'b10111:
        casez_tmp_10 = rob_exception_3_23;
      5'b11000:
        casez_tmp_10 = rob_exception_3_24;
      5'b11001:
        casez_tmp_10 = rob_exception_3_25;
      5'b11010:
        casez_tmp_10 = rob_exception_3_26;
      5'b11011:
        casez_tmp_10 = rob_exception_3_27;
      5'b11100:
        casez_tmp_10 = rob_exception_3_28;
      5'b11101:
        casez_tmp_10 = rob_exception_3_29;
      5'b11110:
        casez_tmp_10 = rob_exception_3_30;
      default:
        casez_tmp_10 = rob_exception_3_31;
    endcase
  end // always @(*)
  wire        can_throw_exception_3 = casez_tmp_8 & casez_tmp_10;
  wire        _GEN_1 = casez_tmp_5 & (~can_commit_2 | can_throw_exception_2) | _GEN_0;
  wire        _io_commit_valids_3_output = casez_tmp_8 & ~casez_tmp_9 & ~io_csr_stall & ~can_throw_exception_3 & ~_GEN_1;
  reg  [4:0]  rob_fflags_0_0;
  reg  [4:0]  rob_fflags_0_1;
  reg  [4:0]  rob_fflags_0_2;
  reg  [4:0]  rob_fflags_0_3;
  reg  [4:0]  rob_fflags_0_4;
  reg  [4:0]  rob_fflags_0_5;
  reg  [4:0]  rob_fflags_0_6;
  reg  [4:0]  rob_fflags_0_7;
  reg  [4:0]  rob_fflags_0_8;
  reg  [4:0]  rob_fflags_0_9;
  reg  [4:0]  rob_fflags_0_10;
  reg  [4:0]  rob_fflags_0_11;
  reg  [4:0]  rob_fflags_0_12;
  reg  [4:0]  rob_fflags_0_13;
  reg  [4:0]  rob_fflags_0_14;
  reg  [4:0]  rob_fflags_0_15;
  reg  [4:0]  rob_fflags_0_16;
  reg  [4:0]  rob_fflags_0_17;
  reg  [4:0]  rob_fflags_0_18;
  reg  [4:0]  rob_fflags_0_19;
  reg  [4:0]  rob_fflags_0_20;
  reg  [4:0]  rob_fflags_0_21;
  reg  [4:0]  rob_fflags_0_22;
  reg  [4:0]  rob_fflags_0_23;
  reg  [4:0]  rob_fflags_0_24;
  reg  [4:0]  rob_fflags_0_25;
  reg  [4:0]  rob_fflags_0_26;
  reg  [4:0]  rob_fflags_0_27;
  reg  [4:0]  rob_fflags_0_28;
  reg  [4:0]  rob_fflags_0_29;
  reg  [4:0]  rob_fflags_0_30;
  reg  [4:0]  rob_fflags_0_31;
  reg  [4:0]  rob_fflags_1_0;
  reg  [4:0]  rob_fflags_1_1;
  reg  [4:0]  rob_fflags_1_2;
  reg  [4:0]  rob_fflags_1_3;
  reg  [4:0]  rob_fflags_1_4;
  reg  [4:0]  rob_fflags_1_5;
  reg  [4:0]  rob_fflags_1_6;
  reg  [4:0]  rob_fflags_1_7;
  reg  [4:0]  rob_fflags_1_8;
  reg  [4:0]  rob_fflags_1_9;
  reg  [4:0]  rob_fflags_1_10;
  reg  [4:0]  rob_fflags_1_11;
  reg  [4:0]  rob_fflags_1_12;
  reg  [4:0]  rob_fflags_1_13;
  reg  [4:0]  rob_fflags_1_14;
  reg  [4:0]  rob_fflags_1_15;
  reg  [4:0]  rob_fflags_1_16;
  reg  [4:0]  rob_fflags_1_17;
  reg  [4:0]  rob_fflags_1_18;
  reg  [4:0]  rob_fflags_1_19;
  reg  [4:0]  rob_fflags_1_20;
  reg  [4:0]  rob_fflags_1_21;
  reg  [4:0]  rob_fflags_1_22;
  reg  [4:0]  rob_fflags_1_23;
  reg  [4:0]  rob_fflags_1_24;
  reg  [4:0]  rob_fflags_1_25;
  reg  [4:0]  rob_fflags_1_26;
  reg  [4:0]  rob_fflags_1_27;
  reg  [4:0]  rob_fflags_1_28;
  reg  [4:0]  rob_fflags_1_29;
  reg  [4:0]  rob_fflags_1_30;
  reg  [4:0]  rob_fflags_1_31;
  reg  [4:0]  rob_fflags_2_0;
  reg  [4:0]  rob_fflags_2_1;
  reg  [4:0]  rob_fflags_2_2;
  reg  [4:0]  rob_fflags_2_3;
  reg  [4:0]  rob_fflags_2_4;
  reg  [4:0]  rob_fflags_2_5;
  reg  [4:0]  rob_fflags_2_6;
  reg  [4:0]  rob_fflags_2_7;
  reg  [4:0]  rob_fflags_2_8;
  reg  [4:0]  rob_fflags_2_9;
  reg  [4:0]  rob_fflags_2_10;
  reg  [4:0]  rob_fflags_2_11;
  reg  [4:0]  rob_fflags_2_12;
  reg  [4:0]  rob_fflags_2_13;
  reg  [4:0]  rob_fflags_2_14;
  reg  [4:0]  rob_fflags_2_15;
  reg  [4:0]  rob_fflags_2_16;
  reg  [4:0]  rob_fflags_2_17;
  reg  [4:0]  rob_fflags_2_18;
  reg  [4:0]  rob_fflags_2_19;
  reg  [4:0]  rob_fflags_2_20;
  reg  [4:0]  rob_fflags_2_21;
  reg  [4:0]  rob_fflags_2_22;
  reg  [4:0]  rob_fflags_2_23;
  reg  [4:0]  rob_fflags_2_24;
  reg  [4:0]  rob_fflags_2_25;
  reg  [4:0]  rob_fflags_2_26;
  reg  [4:0]  rob_fflags_2_27;
  reg  [4:0]  rob_fflags_2_28;
  reg  [4:0]  rob_fflags_2_29;
  reg  [4:0]  rob_fflags_2_30;
  reg  [4:0]  rob_fflags_2_31;
  reg  [4:0]  rob_fflags_3_0;
  reg  [4:0]  rob_fflags_3_1;
  reg  [4:0]  rob_fflags_3_2;
  reg  [4:0]  rob_fflags_3_3;
  reg  [4:0]  rob_fflags_3_4;
  reg  [4:0]  rob_fflags_3_5;
  reg  [4:0]  rob_fflags_3_6;
  reg  [4:0]  rob_fflags_3_7;
  reg  [4:0]  rob_fflags_3_8;
  reg  [4:0]  rob_fflags_3_9;
  reg  [4:0]  rob_fflags_3_10;
  reg  [4:0]  rob_fflags_3_11;
  reg  [4:0]  rob_fflags_3_12;
  reg  [4:0]  rob_fflags_3_13;
  reg  [4:0]  rob_fflags_3_14;
  reg  [4:0]  rob_fflags_3_15;
  reg  [4:0]  rob_fflags_3_16;
  reg  [4:0]  rob_fflags_3_17;
  reg  [4:0]  rob_fflags_3_18;
  reg  [4:0]  rob_fflags_3_19;
  reg  [4:0]  rob_fflags_3_20;
  reg  [4:0]  rob_fflags_3_21;
  reg  [4:0]  rob_fflags_3_22;
  reg  [4:0]  rob_fflags_3_23;
  reg  [4:0]  rob_fflags_3_24;
  reg  [4:0]  rob_fflags_3_25;
  reg  [4:0]  rob_fflags_3_26;
  reg  [4:0]  rob_fflags_3_27;
  reg  [4:0]  rob_fflags_3_28;
  reg  [4:0]  rob_fflags_3_29;
  reg  [4:0]  rob_fflags_3_30;
  reg  [4:0]  rob_fflags_3_31;
  reg  [6:0]  rob_uop__0_uopc;
  reg         rob_uop__0_is_rvc;
  reg  [19:0] rob_uop__0_br_mask;
  reg  [5:0]  rob_uop__0_ftq_idx;
  reg         rob_uop__0_edge_inst;
  reg  [5:0]  rob_uop__0_pc_lob;
  reg  [6:0]  rob_uop__0_pdst;
  reg  [6:0]  rob_uop__0_stale_pdst;
  reg         rob_uop__0_is_fencei;
  reg         rob_uop__0_uses_ldq;
  reg         rob_uop__0_uses_stq;
  reg         rob_uop__0_is_sys_pc2epc;
  reg         rob_uop__0_flush_on_commit;
  reg  [5:0]  rob_uop__0_ldst;
  reg         rob_uop__0_ldst_val;
  reg  [1:0]  rob_uop__0_dst_rtype;
  reg         rob_uop__0_fp_val;
  reg  [6:0]  rob_uop__1_uopc;
  reg         rob_uop__1_is_rvc;
  reg  [19:0] rob_uop__1_br_mask;
  reg  [5:0]  rob_uop__1_ftq_idx;
  reg         rob_uop__1_edge_inst;
  reg  [5:0]  rob_uop__1_pc_lob;
  reg  [6:0]  rob_uop__1_pdst;
  reg  [6:0]  rob_uop__1_stale_pdst;
  reg         rob_uop__1_is_fencei;
  reg         rob_uop__1_uses_ldq;
  reg         rob_uop__1_uses_stq;
  reg         rob_uop__1_is_sys_pc2epc;
  reg         rob_uop__1_flush_on_commit;
  reg  [5:0]  rob_uop__1_ldst;
  reg         rob_uop__1_ldst_val;
  reg  [1:0]  rob_uop__1_dst_rtype;
  reg         rob_uop__1_fp_val;
  reg  [6:0]  rob_uop__2_uopc;
  reg         rob_uop__2_is_rvc;
  reg  [19:0] rob_uop__2_br_mask;
  reg  [5:0]  rob_uop__2_ftq_idx;
  reg         rob_uop__2_edge_inst;
  reg  [5:0]  rob_uop__2_pc_lob;
  reg  [6:0]  rob_uop__2_pdst;
  reg  [6:0]  rob_uop__2_stale_pdst;
  reg         rob_uop__2_is_fencei;
  reg         rob_uop__2_uses_ldq;
  reg         rob_uop__2_uses_stq;
  reg         rob_uop__2_is_sys_pc2epc;
  reg         rob_uop__2_flush_on_commit;
  reg  [5:0]  rob_uop__2_ldst;
  reg         rob_uop__2_ldst_val;
  reg  [1:0]  rob_uop__2_dst_rtype;
  reg         rob_uop__2_fp_val;
  reg  [6:0]  rob_uop__3_uopc;
  reg         rob_uop__3_is_rvc;
  reg  [19:0] rob_uop__3_br_mask;
  reg  [5:0]  rob_uop__3_ftq_idx;
  reg         rob_uop__3_edge_inst;
  reg  [5:0]  rob_uop__3_pc_lob;
  reg  [6:0]  rob_uop__3_pdst;
  reg  [6:0]  rob_uop__3_stale_pdst;
  reg         rob_uop__3_is_fencei;
  reg         rob_uop__3_uses_ldq;
  reg         rob_uop__3_uses_stq;
  reg         rob_uop__3_is_sys_pc2epc;
  reg         rob_uop__3_flush_on_commit;
  reg  [5:0]  rob_uop__3_ldst;
  reg         rob_uop__3_ldst_val;
  reg  [1:0]  rob_uop__3_dst_rtype;
  reg         rob_uop__3_fp_val;
  reg  [6:0]  rob_uop__4_uopc;
  reg         rob_uop__4_is_rvc;
  reg  [19:0] rob_uop__4_br_mask;
  reg  [5:0]  rob_uop__4_ftq_idx;
  reg         rob_uop__4_edge_inst;
  reg  [5:0]  rob_uop__4_pc_lob;
  reg  [6:0]  rob_uop__4_pdst;
  reg  [6:0]  rob_uop__4_stale_pdst;
  reg         rob_uop__4_is_fencei;
  reg         rob_uop__4_uses_ldq;
  reg         rob_uop__4_uses_stq;
  reg         rob_uop__4_is_sys_pc2epc;
  reg         rob_uop__4_flush_on_commit;
  reg  [5:0]  rob_uop__4_ldst;
  reg         rob_uop__4_ldst_val;
  reg  [1:0]  rob_uop__4_dst_rtype;
  reg         rob_uop__4_fp_val;
  reg  [6:0]  rob_uop__5_uopc;
  reg         rob_uop__5_is_rvc;
  reg  [19:0] rob_uop__5_br_mask;
  reg  [5:0]  rob_uop__5_ftq_idx;
  reg         rob_uop__5_edge_inst;
  reg  [5:0]  rob_uop__5_pc_lob;
  reg  [6:0]  rob_uop__5_pdst;
  reg  [6:0]  rob_uop__5_stale_pdst;
  reg         rob_uop__5_is_fencei;
  reg         rob_uop__5_uses_ldq;
  reg         rob_uop__5_uses_stq;
  reg         rob_uop__5_is_sys_pc2epc;
  reg         rob_uop__5_flush_on_commit;
  reg  [5:0]  rob_uop__5_ldst;
  reg         rob_uop__5_ldst_val;
  reg  [1:0]  rob_uop__5_dst_rtype;
  reg         rob_uop__5_fp_val;
  reg  [6:0]  rob_uop__6_uopc;
  reg         rob_uop__6_is_rvc;
  reg  [19:0] rob_uop__6_br_mask;
  reg  [5:0]  rob_uop__6_ftq_idx;
  reg         rob_uop__6_edge_inst;
  reg  [5:0]  rob_uop__6_pc_lob;
  reg  [6:0]  rob_uop__6_pdst;
  reg  [6:0]  rob_uop__6_stale_pdst;
  reg         rob_uop__6_is_fencei;
  reg         rob_uop__6_uses_ldq;
  reg         rob_uop__6_uses_stq;
  reg         rob_uop__6_is_sys_pc2epc;
  reg         rob_uop__6_flush_on_commit;
  reg  [5:0]  rob_uop__6_ldst;
  reg         rob_uop__6_ldst_val;
  reg  [1:0]  rob_uop__6_dst_rtype;
  reg         rob_uop__6_fp_val;
  reg  [6:0]  rob_uop__7_uopc;
  reg         rob_uop__7_is_rvc;
  reg  [19:0] rob_uop__7_br_mask;
  reg  [5:0]  rob_uop__7_ftq_idx;
  reg         rob_uop__7_edge_inst;
  reg  [5:0]  rob_uop__7_pc_lob;
  reg  [6:0]  rob_uop__7_pdst;
  reg  [6:0]  rob_uop__7_stale_pdst;
  reg         rob_uop__7_is_fencei;
  reg         rob_uop__7_uses_ldq;
  reg         rob_uop__7_uses_stq;
  reg         rob_uop__7_is_sys_pc2epc;
  reg         rob_uop__7_flush_on_commit;
  reg  [5:0]  rob_uop__7_ldst;
  reg         rob_uop__7_ldst_val;
  reg  [1:0]  rob_uop__7_dst_rtype;
  reg         rob_uop__7_fp_val;
  reg  [6:0]  rob_uop__8_uopc;
  reg         rob_uop__8_is_rvc;
  reg  [19:0] rob_uop__8_br_mask;
  reg  [5:0]  rob_uop__8_ftq_idx;
  reg         rob_uop__8_edge_inst;
  reg  [5:0]  rob_uop__8_pc_lob;
  reg  [6:0]  rob_uop__8_pdst;
  reg  [6:0]  rob_uop__8_stale_pdst;
  reg         rob_uop__8_is_fencei;
  reg         rob_uop__8_uses_ldq;
  reg         rob_uop__8_uses_stq;
  reg         rob_uop__8_is_sys_pc2epc;
  reg         rob_uop__8_flush_on_commit;
  reg  [5:0]  rob_uop__8_ldst;
  reg         rob_uop__8_ldst_val;
  reg  [1:0]  rob_uop__8_dst_rtype;
  reg         rob_uop__8_fp_val;
  reg  [6:0]  rob_uop__9_uopc;
  reg         rob_uop__9_is_rvc;
  reg  [19:0] rob_uop__9_br_mask;
  reg  [5:0]  rob_uop__9_ftq_idx;
  reg         rob_uop__9_edge_inst;
  reg  [5:0]  rob_uop__9_pc_lob;
  reg  [6:0]  rob_uop__9_pdst;
  reg  [6:0]  rob_uop__9_stale_pdst;
  reg         rob_uop__9_is_fencei;
  reg         rob_uop__9_uses_ldq;
  reg         rob_uop__9_uses_stq;
  reg         rob_uop__9_is_sys_pc2epc;
  reg         rob_uop__9_flush_on_commit;
  reg  [5:0]  rob_uop__9_ldst;
  reg         rob_uop__9_ldst_val;
  reg  [1:0]  rob_uop__9_dst_rtype;
  reg         rob_uop__9_fp_val;
  reg  [6:0]  rob_uop__10_uopc;
  reg         rob_uop__10_is_rvc;
  reg  [19:0] rob_uop__10_br_mask;
  reg  [5:0]  rob_uop__10_ftq_idx;
  reg         rob_uop__10_edge_inst;
  reg  [5:0]  rob_uop__10_pc_lob;
  reg  [6:0]  rob_uop__10_pdst;
  reg  [6:0]  rob_uop__10_stale_pdst;
  reg         rob_uop__10_is_fencei;
  reg         rob_uop__10_uses_ldq;
  reg         rob_uop__10_uses_stq;
  reg         rob_uop__10_is_sys_pc2epc;
  reg         rob_uop__10_flush_on_commit;
  reg  [5:0]  rob_uop__10_ldst;
  reg         rob_uop__10_ldst_val;
  reg  [1:0]  rob_uop__10_dst_rtype;
  reg         rob_uop__10_fp_val;
  reg  [6:0]  rob_uop__11_uopc;
  reg         rob_uop__11_is_rvc;
  reg  [19:0] rob_uop__11_br_mask;
  reg  [5:0]  rob_uop__11_ftq_idx;
  reg         rob_uop__11_edge_inst;
  reg  [5:0]  rob_uop__11_pc_lob;
  reg  [6:0]  rob_uop__11_pdst;
  reg  [6:0]  rob_uop__11_stale_pdst;
  reg         rob_uop__11_is_fencei;
  reg         rob_uop__11_uses_ldq;
  reg         rob_uop__11_uses_stq;
  reg         rob_uop__11_is_sys_pc2epc;
  reg         rob_uop__11_flush_on_commit;
  reg  [5:0]  rob_uop__11_ldst;
  reg         rob_uop__11_ldst_val;
  reg  [1:0]  rob_uop__11_dst_rtype;
  reg         rob_uop__11_fp_val;
  reg  [6:0]  rob_uop__12_uopc;
  reg         rob_uop__12_is_rvc;
  reg  [19:0] rob_uop__12_br_mask;
  reg  [5:0]  rob_uop__12_ftq_idx;
  reg         rob_uop__12_edge_inst;
  reg  [5:0]  rob_uop__12_pc_lob;
  reg  [6:0]  rob_uop__12_pdst;
  reg  [6:0]  rob_uop__12_stale_pdst;
  reg         rob_uop__12_is_fencei;
  reg         rob_uop__12_uses_ldq;
  reg         rob_uop__12_uses_stq;
  reg         rob_uop__12_is_sys_pc2epc;
  reg         rob_uop__12_flush_on_commit;
  reg  [5:0]  rob_uop__12_ldst;
  reg         rob_uop__12_ldst_val;
  reg  [1:0]  rob_uop__12_dst_rtype;
  reg         rob_uop__12_fp_val;
  reg  [6:0]  rob_uop__13_uopc;
  reg         rob_uop__13_is_rvc;
  reg  [19:0] rob_uop__13_br_mask;
  reg  [5:0]  rob_uop__13_ftq_idx;
  reg         rob_uop__13_edge_inst;
  reg  [5:0]  rob_uop__13_pc_lob;
  reg  [6:0]  rob_uop__13_pdst;
  reg  [6:0]  rob_uop__13_stale_pdst;
  reg         rob_uop__13_is_fencei;
  reg         rob_uop__13_uses_ldq;
  reg         rob_uop__13_uses_stq;
  reg         rob_uop__13_is_sys_pc2epc;
  reg         rob_uop__13_flush_on_commit;
  reg  [5:0]  rob_uop__13_ldst;
  reg         rob_uop__13_ldst_val;
  reg  [1:0]  rob_uop__13_dst_rtype;
  reg         rob_uop__13_fp_val;
  reg  [6:0]  rob_uop__14_uopc;
  reg         rob_uop__14_is_rvc;
  reg  [19:0] rob_uop__14_br_mask;
  reg  [5:0]  rob_uop__14_ftq_idx;
  reg         rob_uop__14_edge_inst;
  reg  [5:0]  rob_uop__14_pc_lob;
  reg  [6:0]  rob_uop__14_pdst;
  reg  [6:0]  rob_uop__14_stale_pdst;
  reg         rob_uop__14_is_fencei;
  reg         rob_uop__14_uses_ldq;
  reg         rob_uop__14_uses_stq;
  reg         rob_uop__14_is_sys_pc2epc;
  reg         rob_uop__14_flush_on_commit;
  reg  [5:0]  rob_uop__14_ldst;
  reg         rob_uop__14_ldst_val;
  reg  [1:0]  rob_uop__14_dst_rtype;
  reg         rob_uop__14_fp_val;
  reg  [6:0]  rob_uop__15_uopc;
  reg         rob_uop__15_is_rvc;
  reg  [19:0] rob_uop__15_br_mask;
  reg  [5:0]  rob_uop__15_ftq_idx;
  reg         rob_uop__15_edge_inst;
  reg  [5:0]  rob_uop__15_pc_lob;
  reg  [6:0]  rob_uop__15_pdst;
  reg  [6:0]  rob_uop__15_stale_pdst;
  reg         rob_uop__15_is_fencei;
  reg         rob_uop__15_uses_ldq;
  reg         rob_uop__15_uses_stq;
  reg         rob_uop__15_is_sys_pc2epc;
  reg         rob_uop__15_flush_on_commit;
  reg  [5:0]  rob_uop__15_ldst;
  reg         rob_uop__15_ldst_val;
  reg  [1:0]  rob_uop__15_dst_rtype;
  reg         rob_uop__15_fp_val;
  reg  [6:0]  rob_uop__16_uopc;
  reg         rob_uop__16_is_rvc;
  reg  [19:0] rob_uop__16_br_mask;
  reg  [5:0]  rob_uop__16_ftq_idx;
  reg         rob_uop__16_edge_inst;
  reg  [5:0]  rob_uop__16_pc_lob;
  reg  [6:0]  rob_uop__16_pdst;
  reg  [6:0]  rob_uop__16_stale_pdst;
  reg         rob_uop__16_is_fencei;
  reg         rob_uop__16_uses_ldq;
  reg         rob_uop__16_uses_stq;
  reg         rob_uop__16_is_sys_pc2epc;
  reg         rob_uop__16_flush_on_commit;
  reg  [5:0]  rob_uop__16_ldst;
  reg         rob_uop__16_ldst_val;
  reg  [1:0]  rob_uop__16_dst_rtype;
  reg         rob_uop__16_fp_val;
  reg  [6:0]  rob_uop__17_uopc;
  reg         rob_uop__17_is_rvc;
  reg  [19:0] rob_uop__17_br_mask;
  reg  [5:0]  rob_uop__17_ftq_idx;
  reg         rob_uop__17_edge_inst;
  reg  [5:0]  rob_uop__17_pc_lob;
  reg  [6:0]  rob_uop__17_pdst;
  reg  [6:0]  rob_uop__17_stale_pdst;
  reg         rob_uop__17_is_fencei;
  reg         rob_uop__17_uses_ldq;
  reg         rob_uop__17_uses_stq;
  reg         rob_uop__17_is_sys_pc2epc;
  reg         rob_uop__17_flush_on_commit;
  reg  [5:0]  rob_uop__17_ldst;
  reg         rob_uop__17_ldst_val;
  reg  [1:0]  rob_uop__17_dst_rtype;
  reg         rob_uop__17_fp_val;
  reg  [6:0]  rob_uop__18_uopc;
  reg         rob_uop__18_is_rvc;
  reg  [19:0] rob_uop__18_br_mask;
  reg  [5:0]  rob_uop__18_ftq_idx;
  reg         rob_uop__18_edge_inst;
  reg  [5:0]  rob_uop__18_pc_lob;
  reg  [6:0]  rob_uop__18_pdst;
  reg  [6:0]  rob_uop__18_stale_pdst;
  reg         rob_uop__18_is_fencei;
  reg         rob_uop__18_uses_ldq;
  reg         rob_uop__18_uses_stq;
  reg         rob_uop__18_is_sys_pc2epc;
  reg         rob_uop__18_flush_on_commit;
  reg  [5:0]  rob_uop__18_ldst;
  reg         rob_uop__18_ldst_val;
  reg  [1:0]  rob_uop__18_dst_rtype;
  reg         rob_uop__18_fp_val;
  reg  [6:0]  rob_uop__19_uopc;
  reg         rob_uop__19_is_rvc;
  reg  [19:0] rob_uop__19_br_mask;
  reg  [5:0]  rob_uop__19_ftq_idx;
  reg         rob_uop__19_edge_inst;
  reg  [5:0]  rob_uop__19_pc_lob;
  reg  [6:0]  rob_uop__19_pdst;
  reg  [6:0]  rob_uop__19_stale_pdst;
  reg         rob_uop__19_is_fencei;
  reg         rob_uop__19_uses_ldq;
  reg         rob_uop__19_uses_stq;
  reg         rob_uop__19_is_sys_pc2epc;
  reg         rob_uop__19_flush_on_commit;
  reg  [5:0]  rob_uop__19_ldst;
  reg         rob_uop__19_ldst_val;
  reg  [1:0]  rob_uop__19_dst_rtype;
  reg         rob_uop__19_fp_val;
  reg  [6:0]  rob_uop__20_uopc;
  reg         rob_uop__20_is_rvc;
  reg  [19:0] rob_uop__20_br_mask;
  reg  [5:0]  rob_uop__20_ftq_idx;
  reg         rob_uop__20_edge_inst;
  reg  [5:0]  rob_uop__20_pc_lob;
  reg  [6:0]  rob_uop__20_pdst;
  reg  [6:0]  rob_uop__20_stale_pdst;
  reg         rob_uop__20_is_fencei;
  reg         rob_uop__20_uses_ldq;
  reg         rob_uop__20_uses_stq;
  reg         rob_uop__20_is_sys_pc2epc;
  reg         rob_uop__20_flush_on_commit;
  reg  [5:0]  rob_uop__20_ldst;
  reg         rob_uop__20_ldst_val;
  reg  [1:0]  rob_uop__20_dst_rtype;
  reg         rob_uop__20_fp_val;
  reg  [6:0]  rob_uop__21_uopc;
  reg         rob_uop__21_is_rvc;
  reg  [19:0] rob_uop__21_br_mask;
  reg  [5:0]  rob_uop__21_ftq_idx;
  reg         rob_uop__21_edge_inst;
  reg  [5:0]  rob_uop__21_pc_lob;
  reg  [6:0]  rob_uop__21_pdst;
  reg  [6:0]  rob_uop__21_stale_pdst;
  reg         rob_uop__21_is_fencei;
  reg         rob_uop__21_uses_ldq;
  reg         rob_uop__21_uses_stq;
  reg         rob_uop__21_is_sys_pc2epc;
  reg         rob_uop__21_flush_on_commit;
  reg  [5:0]  rob_uop__21_ldst;
  reg         rob_uop__21_ldst_val;
  reg  [1:0]  rob_uop__21_dst_rtype;
  reg         rob_uop__21_fp_val;
  reg  [6:0]  rob_uop__22_uopc;
  reg         rob_uop__22_is_rvc;
  reg  [19:0] rob_uop__22_br_mask;
  reg  [5:0]  rob_uop__22_ftq_idx;
  reg         rob_uop__22_edge_inst;
  reg  [5:0]  rob_uop__22_pc_lob;
  reg  [6:0]  rob_uop__22_pdst;
  reg  [6:0]  rob_uop__22_stale_pdst;
  reg         rob_uop__22_is_fencei;
  reg         rob_uop__22_uses_ldq;
  reg         rob_uop__22_uses_stq;
  reg         rob_uop__22_is_sys_pc2epc;
  reg         rob_uop__22_flush_on_commit;
  reg  [5:0]  rob_uop__22_ldst;
  reg         rob_uop__22_ldst_val;
  reg  [1:0]  rob_uop__22_dst_rtype;
  reg         rob_uop__22_fp_val;
  reg  [6:0]  rob_uop__23_uopc;
  reg         rob_uop__23_is_rvc;
  reg  [19:0] rob_uop__23_br_mask;
  reg  [5:0]  rob_uop__23_ftq_idx;
  reg         rob_uop__23_edge_inst;
  reg  [5:0]  rob_uop__23_pc_lob;
  reg  [6:0]  rob_uop__23_pdst;
  reg  [6:0]  rob_uop__23_stale_pdst;
  reg         rob_uop__23_is_fencei;
  reg         rob_uop__23_uses_ldq;
  reg         rob_uop__23_uses_stq;
  reg         rob_uop__23_is_sys_pc2epc;
  reg         rob_uop__23_flush_on_commit;
  reg  [5:0]  rob_uop__23_ldst;
  reg         rob_uop__23_ldst_val;
  reg  [1:0]  rob_uop__23_dst_rtype;
  reg         rob_uop__23_fp_val;
  reg  [6:0]  rob_uop__24_uopc;
  reg         rob_uop__24_is_rvc;
  reg  [19:0] rob_uop__24_br_mask;
  reg  [5:0]  rob_uop__24_ftq_idx;
  reg         rob_uop__24_edge_inst;
  reg  [5:0]  rob_uop__24_pc_lob;
  reg  [6:0]  rob_uop__24_pdst;
  reg  [6:0]  rob_uop__24_stale_pdst;
  reg         rob_uop__24_is_fencei;
  reg         rob_uop__24_uses_ldq;
  reg         rob_uop__24_uses_stq;
  reg         rob_uop__24_is_sys_pc2epc;
  reg         rob_uop__24_flush_on_commit;
  reg  [5:0]  rob_uop__24_ldst;
  reg         rob_uop__24_ldst_val;
  reg  [1:0]  rob_uop__24_dst_rtype;
  reg         rob_uop__24_fp_val;
  reg  [6:0]  rob_uop__25_uopc;
  reg         rob_uop__25_is_rvc;
  reg  [19:0] rob_uop__25_br_mask;
  reg  [5:0]  rob_uop__25_ftq_idx;
  reg         rob_uop__25_edge_inst;
  reg  [5:0]  rob_uop__25_pc_lob;
  reg  [6:0]  rob_uop__25_pdst;
  reg  [6:0]  rob_uop__25_stale_pdst;
  reg         rob_uop__25_is_fencei;
  reg         rob_uop__25_uses_ldq;
  reg         rob_uop__25_uses_stq;
  reg         rob_uop__25_is_sys_pc2epc;
  reg         rob_uop__25_flush_on_commit;
  reg  [5:0]  rob_uop__25_ldst;
  reg         rob_uop__25_ldst_val;
  reg  [1:0]  rob_uop__25_dst_rtype;
  reg         rob_uop__25_fp_val;
  reg  [6:0]  rob_uop__26_uopc;
  reg         rob_uop__26_is_rvc;
  reg  [19:0] rob_uop__26_br_mask;
  reg  [5:0]  rob_uop__26_ftq_idx;
  reg         rob_uop__26_edge_inst;
  reg  [5:0]  rob_uop__26_pc_lob;
  reg  [6:0]  rob_uop__26_pdst;
  reg  [6:0]  rob_uop__26_stale_pdst;
  reg         rob_uop__26_is_fencei;
  reg         rob_uop__26_uses_ldq;
  reg         rob_uop__26_uses_stq;
  reg         rob_uop__26_is_sys_pc2epc;
  reg         rob_uop__26_flush_on_commit;
  reg  [5:0]  rob_uop__26_ldst;
  reg         rob_uop__26_ldst_val;
  reg  [1:0]  rob_uop__26_dst_rtype;
  reg         rob_uop__26_fp_val;
  reg  [6:0]  rob_uop__27_uopc;
  reg         rob_uop__27_is_rvc;
  reg  [19:0] rob_uop__27_br_mask;
  reg  [5:0]  rob_uop__27_ftq_idx;
  reg         rob_uop__27_edge_inst;
  reg  [5:0]  rob_uop__27_pc_lob;
  reg  [6:0]  rob_uop__27_pdst;
  reg  [6:0]  rob_uop__27_stale_pdst;
  reg         rob_uop__27_is_fencei;
  reg         rob_uop__27_uses_ldq;
  reg         rob_uop__27_uses_stq;
  reg         rob_uop__27_is_sys_pc2epc;
  reg         rob_uop__27_flush_on_commit;
  reg  [5:0]  rob_uop__27_ldst;
  reg         rob_uop__27_ldst_val;
  reg  [1:0]  rob_uop__27_dst_rtype;
  reg         rob_uop__27_fp_val;
  reg  [6:0]  rob_uop__28_uopc;
  reg         rob_uop__28_is_rvc;
  reg  [19:0] rob_uop__28_br_mask;
  reg  [5:0]  rob_uop__28_ftq_idx;
  reg         rob_uop__28_edge_inst;
  reg  [5:0]  rob_uop__28_pc_lob;
  reg  [6:0]  rob_uop__28_pdst;
  reg  [6:0]  rob_uop__28_stale_pdst;
  reg         rob_uop__28_is_fencei;
  reg         rob_uop__28_uses_ldq;
  reg         rob_uop__28_uses_stq;
  reg         rob_uop__28_is_sys_pc2epc;
  reg         rob_uop__28_flush_on_commit;
  reg  [5:0]  rob_uop__28_ldst;
  reg         rob_uop__28_ldst_val;
  reg  [1:0]  rob_uop__28_dst_rtype;
  reg         rob_uop__28_fp_val;
  reg  [6:0]  rob_uop__29_uopc;
  reg         rob_uop__29_is_rvc;
  reg  [19:0] rob_uop__29_br_mask;
  reg  [5:0]  rob_uop__29_ftq_idx;
  reg         rob_uop__29_edge_inst;
  reg  [5:0]  rob_uop__29_pc_lob;
  reg  [6:0]  rob_uop__29_pdst;
  reg  [6:0]  rob_uop__29_stale_pdst;
  reg         rob_uop__29_is_fencei;
  reg         rob_uop__29_uses_ldq;
  reg         rob_uop__29_uses_stq;
  reg         rob_uop__29_is_sys_pc2epc;
  reg         rob_uop__29_flush_on_commit;
  reg  [5:0]  rob_uop__29_ldst;
  reg         rob_uop__29_ldst_val;
  reg  [1:0]  rob_uop__29_dst_rtype;
  reg         rob_uop__29_fp_val;
  reg  [6:0]  rob_uop__30_uopc;
  reg         rob_uop__30_is_rvc;
  reg  [19:0] rob_uop__30_br_mask;
  reg  [5:0]  rob_uop__30_ftq_idx;
  reg         rob_uop__30_edge_inst;
  reg  [5:0]  rob_uop__30_pc_lob;
  reg  [6:0]  rob_uop__30_pdst;
  reg  [6:0]  rob_uop__30_stale_pdst;
  reg         rob_uop__30_is_fencei;
  reg         rob_uop__30_uses_ldq;
  reg         rob_uop__30_uses_stq;
  reg         rob_uop__30_is_sys_pc2epc;
  reg         rob_uop__30_flush_on_commit;
  reg  [5:0]  rob_uop__30_ldst;
  reg         rob_uop__30_ldst_val;
  reg  [1:0]  rob_uop__30_dst_rtype;
  reg         rob_uop__30_fp_val;
  reg  [6:0]  rob_uop__31_uopc;
  reg         rob_uop__31_is_rvc;
  reg  [19:0] rob_uop__31_br_mask;
  reg  [5:0]  rob_uop__31_ftq_idx;
  reg         rob_uop__31_edge_inst;
  reg  [5:0]  rob_uop__31_pc_lob;
  reg  [6:0]  rob_uop__31_pdst;
  reg  [6:0]  rob_uop__31_stale_pdst;
  reg         rob_uop__31_is_fencei;
  reg         rob_uop__31_uses_ldq;
  reg         rob_uop__31_uses_stq;
  reg         rob_uop__31_is_sys_pc2epc;
  reg         rob_uop__31_flush_on_commit;
  reg  [5:0]  rob_uop__31_ldst;
  reg         rob_uop__31_ldst_val;
  reg  [1:0]  rob_uop__31_dst_rtype;
  reg         rob_uop__31_fp_val;
  reg         rob_predicated__0;
  reg         rob_predicated__1;
  reg         rob_predicated__2;
  reg         rob_predicated__3;
  reg         rob_predicated__4;
  reg         rob_predicated__5;
  reg         rob_predicated__6;
  reg         rob_predicated__7;
  reg         rob_predicated__8;
  reg         rob_predicated__9;
  reg         rob_predicated__10;
  reg         rob_predicated__11;
  reg         rob_predicated__12;
  reg         rob_predicated__13;
  reg         rob_predicated__14;
  reg         rob_predicated__15;
  reg         rob_predicated__16;
  reg         rob_predicated__17;
  reg         rob_predicated__18;
  reg         rob_predicated__19;
  reg         rob_predicated__20;
  reg         rob_predicated__21;
  reg         rob_predicated__22;
  reg         rob_predicated__23;
  reg         rob_predicated__24;
  reg         rob_predicated__25;
  reg         rob_predicated__26;
  reg         rob_predicated__27;
  reg         rob_predicated__28;
  reg         rob_predicated__29;
  reg         rob_predicated__30;
  reg         rob_predicated__31;
  wire        _GEN_2 = rob_tail == 5'h0;
  wire        _GEN_3 = rob_tail == 5'h1;
  wire        _GEN_4 = rob_tail == 5'h2;
  wire        _GEN_5 = rob_tail == 5'h3;
  wire        _GEN_6 = rob_tail == 5'h4;
  wire        _GEN_7 = rob_tail == 5'h5;
  wire        _GEN_8 = rob_tail == 5'h6;
  wire        _GEN_9 = rob_tail == 5'h7;
  wire        _GEN_10 = rob_tail == 5'h8;
  wire        _GEN_11 = rob_tail == 5'h9;
  wire        _GEN_12 = rob_tail == 5'hA;
  wire        _GEN_13 = rob_tail == 5'hB;
  wire        _GEN_14 = rob_tail == 5'hC;
  wire        _GEN_15 = rob_tail == 5'hD;
  wire        _GEN_16 = rob_tail == 5'hE;
  wire        _GEN_17 = rob_tail == 5'hF;
  wire        _GEN_18 = rob_tail == 5'h10;
  wire        _GEN_19 = rob_tail == 5'h11;
  wire        _GEN_20 = rob_tail == 5'h12;
  wire        _GEN_21 = rob_tail == 5'h13;
  wire        _GEN_22 = rob_tail == 5'h14;
  wire        _GEN_23 = rob_tail == 5'h15;
  wire        _GEN_24 = rob_tail == 5'h16;
  wire        _GEN_25 = rob_tail == 5'h17;
  wire        _GEN_26 = rob_tail == 5'h18;
  wire        _GEN_27 = rob_tail == 5'h19;
  wire        _GEN_28 = rob_tail == 5'h1A;
  wire        _GEN_29 = rob_tail == 5'h1B;
  wire        _GEN_30 = rob_tail == 5'h1C;
  wire        _GEN_31 = rob_tail == 5'h1D;
  wire        _GEN_32 = rob_tail == 5'h1E;
  wire        _GEN_33 = io_enq_valids_0 & _GEN_2;
  wire        _GEN_34 = io_enq_valids_0 & _GEN_3;
  wire        _GEN_35 = io_enq_valids_0 & _GEN_4;
  wire        _GEN_36 = io_enq_valids_0 & _GEN_5;
  wire        _GEN_37 = io_enq_valids_0 & _GEN_6;
  wire        _GEN_38 = io_enq_valids_0 & _GEN_7;
  wire        _GEN_39 = io_enq_valids_0 & _GEN_8;
  wire        _GEN_40 = io_enq_valids_0 & _GEN_9;
  wire        _GEN_41 = io_enq_valids_0 & _GEN_10;
  wire        _GEN_42 = io_enq_valids_0 & _GEN_11;
  wire        _GEN_43 = io_enq_valids_0 & _GEN_12;
  wire        _GEN_44 = io_enq_valids_0 & _GEN_13;
  wire        _GEN_45 = io_enq_valids_0 & _GEN_14;
  wire        _GEN_46 = io_enq_valids_0 & _GEN_15;
  wire        _GEN_47 = io_enq_valids_0 & _GEN_16;
  wire        _GEN_48 = io_enq_valids_0 & _GEN_17;
  wire        _GEN_49 = io_enq_valids_0 & _GEN_18;
  wire        _GEN_50 = io_enq_valids_0 & _GEN_19;
  wire        _GEN_51 = io_enq_valids_0 & _GEN_20;
  wire        _GEN_52 = io_enq_valids_0 & _GEN_21;
  wire        _GEN_53 = io_enq_valids_0 & _GEN_22;
  wire        _GEN_54 = io_enq_valids_0 & _GEN_23;
  wire        _GEN_55 = io_enq_valids_0 & _GEN_24;
  wire        _GEN_56 = io_enq_valids_0 & _GEN_25;
  wire        _GEN_57 = io_enq_valids_0 & _GEN_26;
  wire        _GEN_58 = io_enq_valids_0 & _GEN_27;
  wire        _GEN_59 = io_enq_valids_0 & _GEN_28;
  wire        _GEN_60 = io_enq_valids_0 & _GEN_29;
  wire        _GEN_61 = io_enq_valids_0 & _GEN_30;
  wire        _GEN_62 = io_enq_valids_0 & _GEN_31;
  wire        _GEN_63 = io_enq_valids_0 & _GEN_32;
  wire        _GEN_64 = io_enq_valids_0 & (&rob_tail);
  wire        _GEN_65 = io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_66 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_67 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_68 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_69 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_70 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_71 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_72 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_73 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_74 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_75 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_76 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_77 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_78 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_79 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_80 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_81 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_82 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_83 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_84 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_85 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_86 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_87 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_88 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_89 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_90 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_91 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_92 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_93 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_94 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_95 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_96 = io_wb_resps_0_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_97 = _GEN_65 & _GEN_66;
  wire        _GEN_98 = _GEN_65 & _GEN_67;
  wire        _GEN_99 = _GEN_65 & _GEN_68;
  wire        _GEN_100 = _GEN_65 & _GEN_69;
  wire        _GEN_101 = _GEN_65 & _GEN_70;
  wire        _GEN_102 = _GEN_65 & _GEN_71;
  wire        _GEN_103 = _GEN_65 & _GEN_72;
  wire        _GEN_104 = _GEN_65 & _GEN_73;
  wire        _GEN_105 = _GEN_65 & _GEN_74;
  wire        _GEN_106 = _GEN_65 & _GEN_75;
  wire        _GEN_107 = _GEN_65 & _GEN_76;
  wire        _GEN_108 = _GEN_65 & _GEN_77;
  wire        _GEN_109 = _GEN_65 & _GEN_78;
  wire        _GEN_110 = _GEN_65 & _GEN_79;
  wire        _GEN_111 = _GEN_65 & _GEN_80;
  wire        _GEN_112 = _GEN_65 & _GEN_81;
  wire        _GEN_113 = _GEN_65 & _GEN_82;
  wire        _GEN_114 = _GEN_65 & _GEN_83;
  wire        _GEN_115 = _GEN_65 & _GEN_84;
  wire        _GEN_116 = _GEN_65 & _GEN_85;
  wire        _GEN_117 = _GEN_65 & _GEN_86;
  wire        _GEN_118 = _GEN_65 & _GEN_87;
  wire        _GEN_119 = _GEN_65 & _GEN_88;
  wire        _GEN_120 = _GEN_65 & _GEN_89;
  wire        _GEN_121 = _GEN_65 & _GEN_90;
  wire        _GEN_122 = _GEN_65 & _GEN_91;
  wire        _GEN_123 = _GEN_65 & _GEN_92;
  wire        _GEN_124 = _GEN_65 & _GEN_93;
  wire        _GEN_125 = _GEN_65 & _GEN_94;
  wire        _GEN_126 = _GEN_65 & _GEN_95;
  wire        _GEN_127 = _GEN_65 & _GEN_96;
  wire        _GEN_128 = _GEN_65 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_129 = io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_130 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_131 = _GEN_130 | _GEN_97;
  wire        _GEN_132 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_133 = _GEN_132 | _GEN_98;
  wire        _GEN_134 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_135 = _GEN_134 | _GEN_99;
  wire        _GEN_136 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_137 = _GEN_136 | _GEN_100;
  wire        _GEN_138 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_139 = _GEN_138 | _GEN_101;
  wire        _GEN_140 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_141 = _GEN_140 | _GEN_102;
  wire        _GEN_142 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_143 = _GEN_142 | _GEN_103;
  wire        _GEN_144 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_145 = _GEN_144 | _GEN_104;
  wire        _GEN_146 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_147 = _GEN_146 | _GEN_105;
  wire        _GEN_148 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_149 = _GEN_148 | _GEN_106;
  wire        _GEN_150 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_151 = _GEN_150 | _GEN_107;
  wire        _GEN_152 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_153 = _GEN_152 | _GEN_108;
  wire        _GEN_154 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_155 = _GEN_154 | _GEN_109;
  wire        _GEN_156 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_157 = _GEN_156 | _GEN_110;
  wire        _GEN_158 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_159 = _GEN_158 | _GEN_111;
  wire        _GEN_160 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_161 = _GEN_160 | _GEN_112;
  wire        _GEN_162 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_163 = _GEN_162 | _GEN_113;
  wire        _GEN_164 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_165 = _GEN_164 | _GEN_114;
  wire        _GEN_166 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_167 = _GEN_166 | _GEN_115;
  wire        _GEN_168 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_169 = _GEN_168 | _GEN_116;
  wire        _GEN_170 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_171 = _GEN_170 | _GEN_117;
  wire        _GEN_172 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_173 = _GEN_172 | _GEN_118;
  wire        _GEN_174 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_175 = _GEN_174 | _GEN_119;
  wire        _GEN_176 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_177 = _GEN_176 | _GEN_120;
  wire        _GEN_178 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_179 = _GEN_178 | _GEN_121;
  wire        _GEN_180 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_181 = _GEN_180 | _GEN_122;
  wire        _GEN_182 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_183 = _GEN_182 | _GEN_123;
  wire        _GEN_184 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_185 = _GEN_184 | _GEN_124;
  wire        _GEN_186 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_187 = _GEN_186 | _GEN_125;
  wire        _GEN_188 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_189 = _GEN_188 | _GEN_126;
  wire        _GEN_190 = io_wb_resps_1_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_191 = _GEN_190 | _GEN_127;
  wire        _GEN_192 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_128;
  wire        _GEN_193 = io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_194 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_195 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_196 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_197 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_198 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_199 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_200 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_201 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_202 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_203 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_204 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_205 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_206 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_207 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_208 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_209 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_210 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_211 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_212 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_213 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_214 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_215 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_216 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_217 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_218 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_219 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_220 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_221 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_222 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_223 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_224 = io_wb_resps_2_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_225 = _GEN_193 & _GEN_194;
  wire        _GEN_226 = _GEN_193 & _GEN_195;
  wire        _GEN_227 = _GEN_193 & _GEN_196;
  wire        _GEN_228 = _GEN_193 & _GEN_197;
  wire        _GEN_229 = _GEN_193 & _GEN_198;
  wire        _GEN_230 = _GEN_193 & _GEN_199;
  wire        _GEN_231 = _GEN_193 & _GEN_200;
  wire        _GEN_232 = _GEN_193 & _GEN_201;
  wire        _GEN_233 = _GEN_193 & _GEN_202;
  wire        _GEN_234 = _GEN_193 & _GEN_203;
  wire        _GEN_235 = _GEN_193 & _GEN_204;
  wire        _GEN_236 = _GEN_193 & _GEN_205;
  wire        _GEN_237 = _GEN_193 & _GEN_206;
  wire        _GEN_238 = _GEN_193 & _GEN_207;
  wire        _GEN_239 = _GEN_193 & _GEN_208;
  wire        _GEN_240 = _GEN_193 & _GEN_209;
  wire        _GEN_241 = _GEN_193 & _GEN_210;
  wire        _GEN_242 = _GEN_193 & _GEN_211;
  wire        _GEN_243 = _GEN_193 & _GEN_212;
  wire        _GEN_244 = _GEN_193 & _GEN_213;
  wire        _GEN_245 = _GEN_193 & _GEN_214;
  wire        _GEN_246 = _GEN_193 & _GEN_215;
  wire        _GEN_247 = _GEN_193 & _GEN_216;
  wire        _GEN_248 = _GEN_193 & _GEN_217;
  wire        _GEN_249 = _GEN_193 & _GEN_218;
  wire        _GEN_250 = _GEN_193 & _GEN_219;
  wire        _GEN_251 = _GEN_193 & _GEN_220;
  wire        _GEN_252 = _GEN_193 & _GEN_221;
  wire        _GEN_253 = _GEN_193 & _GEN_222;
  wire        _GEN_254 = _GEN_193 & _GEN_223;
  wire        _GEN_255 = _GEN_193 & _GEN_224;
  wire        _GEN_256 = _GEN_193 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_257 = io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_258 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_259 = _GEN_258 | _GEN_225;
  wire        _GEN_260 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_261 = _GEN_260 | _GEN_226;
  wire        _GEN_262 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_263 = _GEN_262 | _GEN_227;
  wire        _GEN_264 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_265 = _GEN_264 | _GEN_228;
  wire        _GEN_266 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_267 = _GEN_266 | _GEN_229;
  wire        _GEN_268 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_269 = _GEN_268 | _GEN_230;
  wire        _GEN_270 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_271 = _GEN_270 | _GEN_231;
  wire        _GEN_272 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_273 = _GEN_272 | _GEN_232;
  wire        _GEN_274 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_275 = _GEN_274 | _GEN_233;
  wire        _GEN_276 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_277 = _GEN_276 | _GEN_234;
  wire        _GEN_278 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_279 = _GEN_278 | _GEN_235;
  wire        _GEN_280 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_281 = _GEN_280 | _GEN_236;
  wire        _GEN_282 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_283 = _GEN_282 | _GEN_237;
  wire        _GEN_284 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_285 = _GEN_284 | _GEN_238;
  wire        _GEN_286 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_287 = _GEN_286 | _GEN_239;
  wire        _GEN_288 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_289 = _GEN_288 | _GEN_240;
  wire        _GEN_290 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_291 = _GEN_290 | _GEN_241;
  wire        _GEN_292 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_293 = _GEN_292 | _GEN_242;
  wire        _GEN_294 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_295 = _GEN_294 | _GEN_243;
  wire        _GEN_296 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_297 = _GEN_296 | _GEN_244;
  wire        _GEN_298 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_299 = _GEN_298 | _GEN_245;
  wire        _GEN_300 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_301 = _GEN_300 | _GEN_246;
  wire        _GEN_302 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_303 = _GEN_302 | _GEN_247;
  wire        _GEN_304 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_305 = _GEN_304 | _GEN_248;
  wire        _GEN_306 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_307 = _GEN_306 | _GEN_249;
  wire        _GEN_308 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_309 = _GEN_308 | _GEN_250;
  wire        _GEN_310 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_311 = _GEN_310 | _GEN_251;
  wire        _GEN_312 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_313 = _GEN_312 | _GEN_252;
  wire        _GEN_314 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_315 = _GEN_314 | _GEN_253;
  wire        _GEN_316 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_317 = _GEN_316 | _GEN_254;
  wire        _GEN_318 = io_wb_resps_3_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_319 = _GEN_318 | _GEN_255;
  wire        _GEN_320 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_256;
  wire        _GEN_321 = io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_322 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_323 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_324 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_325 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_326 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_327 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_328 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_329 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_330 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_331 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_332 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_333 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_334 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_335 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_336 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_337 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_338 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_339 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_340 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_341 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_342 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_343 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_344 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_345 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_346 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_347 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_348 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_349 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_350 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_351 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_352 = io_wb_resps_4_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_353 = _GEN_321 & _GEN_322;
  wire        _GEN_354 = _GEN_321 & _GEN_323;
  wire        _GEN_355 = _GEN_321 & _GEN_324;
  wire        _GEN_356 = _GEN_321 & _GEN_325;
  wire        _GEN_357 = _GEN_321 & _GEN_326;
  wire        _GEN_358 = _GEN_321 & _GEN_327;
  wire        _GEN_359 = _GEN_321 & _GEN_328;
  wire        _GEN_360 = _GEN_321 & _GEN_329;
  wire        _GEN_361 = _GEN_321 & _GEN_330;
  wire        _GEN_362 = _GEN_321 & _GEN_331;
  wire        _GEN_363 = _GEN_321 & _GEN_332;
  wire        _GEN_364 = _GEN_321 & _GEN_333;
  wire        _GEN_365 = _GEN_321 & _GEN_334;
  wire        _GEN_366 = _GEN_321 & _GEN_335;
  wire        _GEN_367 = _GEN_321 & _GEN_336;
  wire        _GEN_368 = _GEN_321 & _GEN_337;
  wire        _GEN_369 = _GEN_321 & _GEN_338;
  wire        _GEN_370 = _GEN_321 & _GEN_339;
  wire        _GEN_371 = _GEN_321 & _GEN_340;
  wire        _GEN_372 = _GEN_321 & _GEN_341;
  wire        _GEN_373 = _GEN_321 & _GEN_342;
  wire        _GEN_374 = _GEN_321 & _GEN_343;
  wire        _GEN_375 = _GEN_321 & _GEN_344;
  wire        _GEN_376 = _GEN_321 & _GEN_345;
  wire        _GEN_377 = _GEN_321 & _GEN_346;
  wire        _GEN_378 = _GEN_321 & _GEN_347;
  wire        _GEN_379 = _GEN_321 & _GEN_348;
  wire        _GEN_380 = _GEN_321 & _GEN_349;
  wire        _GEN_381 = _GEN_321 & _GEN_350;
  wire        _GEN_382 = _GEN_321 & _GEN_351;
  wire        _GEN_383 = _GEN_321 & _GEN_352;
  wire        _GEN_384 = _GEN_321 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_385 = io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_386 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_387 = _GEN_386 | _GEN_353;
  wire        _GEN_388 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_389 = _GEN_388 | _GEN_354;
  wire        _GEN_390 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_391 = _GEN_390 | _GEN_355;
  wire        _GEN_392 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_393 = _GEN_392 | _GEN_356;
  wire        _GEN_394 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_395 = _GEN_394 | _GEN_357;
  wire        _GEN_396 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_397 = _GEN_396 | _GEN_358;
  wire        _GEN_398 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_399 = _GEN_398 | _GEN_359;
  wire        _GEN_400 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_401 = _GEN_400 | _GEN_360;
  wire        _GEN_402 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_403 = _GEN_402 | _GEN_361;
  wire        _GEN_404 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_405 = _GEN_404 | _GEN_362;
  wire        _GEN_406 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_407 = _GEN_406 | _GEN_363;
  wire        _GEN_408 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_409 = _GEN_408 | _GEN_364;
  wire        _GEN_410 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_411 = _GEN_410 | _GEN_365;
  wire        _GEN_412 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_413 = _GEN_412 | _GEN_366;
  wire        _GEN_414 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_415 = _GEN_414 | _GEN_367;
  wire        _GEN_416 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_417 = _GEN_416 | _GEN_368;
  wire        _GEN_418 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_419 = _GEN_418 | _GEN_369;
  wire        _GEN_420 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_421 = _GEN_420 | _GEN_370;
  wire        _GEN_422 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_423 = _GEN_422 | _GEN_371;
  wire        _GEN_424 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_425 = _GEN_424 | _GEN_372;
  wire        _GEN_426 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_427 = _GEN_426 | _GEN_373;
  wire        _GEN_428 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_429 = _GEN_428 | _GEN_374;
  wire        _GEN_430 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_431 = _GEN_430 | _GEN_375;
  wire        _GEN_432 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_433 = _GEN_432 | _GEN_376;
  wire        _GEN_434 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_435 = _GEN_434 | _GEN_377;
  wire        _GEN_436 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_437 = _GEN_436 | _GEN_378;
  wire        _GEN_438 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_439 = _GEN_438 | _GEN_379;
  wire        _GEN_440 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_441 = _GEN_440 | _GEN_380;
  wire        _GEN_442 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_443 = _GEN_442 | _GEN_381;
  wire        _GEN_444 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_445 = _GEN_444 | _GEN_382;
  wire        _GEN_446 = io_wb_resps_5_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_447 = _GEN_446 | _GEN_383;
  wire        _GEN_448 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_384;
  wire        _GEN_449 = io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_450 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_451 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_452 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_453 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_454 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_455 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_456 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_457 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_458 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_459 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_460 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_461 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_462 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_463 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_464 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_465 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_466 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_467 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_468 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_469 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_470 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_471 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_472 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_473 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_474 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_475 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_476 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_477 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_478 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_479 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_480 = io_wb_resps_6_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_481 = _GEN_449 & _GEN_450;
  wire        _GEN_482 = _GEN_449 & _GEN_451;
  wire        _GEN_483 = _GEN_449 & _GEN_452;
  wire        _GEN_484 = _GEN_449 & _GEN_453;
  wire        _GEN_485 = _GEN_449 & _GEN_454;
  wire        _GEN_486 = _GEN_449 & _GEN_455;
  wire        _GEN_487 = _GEN_449 & _GEN_456;
  wire        _GEN_488 = _GEN_449 & _GEN_457;
  wire        _GEN_489 = _GEN_449 & _GEN_458;
  wire        _GEN_490 = _GEN_449 & _GEN_459;
  wire        _GEN_491 = _GEN_449 & _GEN_460;
  wire        _GEN_492 = _GEN_449 & _GEN_461;
  wire        _GEN_493 = _GEN_449 & _GEN_462;
  wire        _GEN_494 = _GEN_449 & _GEN_463;
  wire        _GEN_495 = _GEN_449 & _GEN_464;
  wire        _GEN_496 = _GEN_449 & _GEN_465;
  wire        _GEN_497 = _GEN_449 & _GEN_466;
  wire        _GEN_498 = _GEN_449 & _GEN_467;
  wire        _GEN_499 = _GEN_449 & _GEN_468;
  wire        _GEN_500 = _GEN_449 & _GEN_469;
  wire        _GEN_501 = _GEN_449 & _GEN_470;
  wire        _GEN_502 = _GEN_449 & _GEN_471;
  wire        _GEN_503 = _GEN_449 & _GEN_472;
  wire        _GEN_504 = _GEN_449 & _GEN_473;
  wire        _GEN_505 = _GEN_449 & _GEN_474;
  wire        _GEN_506 = _GEN_449 & _GEN_475;
  wire        _GEN_507 = _GEN_449 & _GEN_476;
  wire        _GEN_508 = _GEN_449 & _GEN_477;
  wire        _GEN_509 = _GEN_449 & _GEN_478;
  wire        _GEN_510 = _GEN_449 & _GEN_479;
  wire        _GEN_511 = _GEN_449 & _GEN_480;
  wire        _GEN_512 = _GEN_449 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_513 = io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_514 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_515 = _GEN_514 | _GEN_481;
  wire        _GEN_516 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_517 = _GEN_516 | _GEN_482;
  wire        _GEN_518 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_519 = _GEN_518 | _GEN_483;
  wire        _GEN_520 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_521 = _GEN_520 | _GEN_484;
  wire        _GEN_522 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_523 = _GEN_522 | _GEN_485;
  wire        _GEN_524 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_525 = _GEN_524 | _GEN_486;
  wire        _GEN_526 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_527 = _GEN_526 | _GEN_487;
  wire        _GEN_528 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_529 = _GEN_528 | _GEN_488;
  wire        _GEN_530 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_531 = _GEN_530 | _GEN_489;
  wire        _GEN_532 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_533 = _GEN_532 | _GEN_490;
  wire        _GEN_534 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_535 = _GEN_534 | _GEN_491;
  wire        _GEN_536 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_537 = _GEN_536 | _GEN_492;
  wire        _GEN_538 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_539 = _GEN_538 | _GEN_493;
  wire        _GEN_540 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_541 = _GEN_540 | _GEN_494;
  wire        _GEN_542 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_543 = _GEN_542 | _GEN_495;
  wire        _GEN_544 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_545 = _GEN_544 | _GEN_496;
  wire        _GEN_546 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_547 = _GEN_546 | _GEN_497;
  wire        _GEN_548 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_549 = _GEN_548 | _GEN_498;
  wire        _GEN_550 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_551 = _GEN_550 | _GEN_499;
  wire        _GEN_552 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_553 = _GEN_552 | _GEN_500;
  wire        _GEN_554 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_555 = _GEN_554 | _GEN_501;
  wire        _GEN_556 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_557 = _GEN_556 | _GEN_502;
  wire        _GEN_558 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_559 = _GEN_558 | _GEN_503;
  wire        _GEN_560 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_561 = _GEN_560 | _GEN_504;
  wire        _GEN_562 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_563 = _GEN_562 | _GEN_505;
  wire        _GEN_564 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_565 = _GEN_564 | _GEN_506;
  wire        _GEN_566 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_567 = _GEN_566 | _GEN_507;
  wire        _GEN_568 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_569 = _GEN_568 | _GEN_508;
  wire        _GEN_570 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_571 = _GEN_570 | _GEN_509;
  wire        _GEN_572 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_573 = _GEN_572 | _GEN_510;
  wire        _GEN_574 = io_wb_resps_7_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_575 = _GEN_574 | _GEN_511;
  wire        _GEN_576 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_512;
  wire        _GEN_577 = io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_578 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_579 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_580 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_581 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_582 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_583 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_584 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_585 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_586 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_587 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_588 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_589 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_590 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_591 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_592 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_593 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_594 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_595 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_596 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_597 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_598 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_599 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_600 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_601 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_602 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_603 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_604 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_605 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_606 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_607 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_608 = io_wb_resps_8_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_609 = _GEN_577 & _GEN_578;
  wire        _GEN_610 = _GEN_577 & _GEN_579;
  wire        _GEN_611 = _GEN_577 & _GEN_580;
  wire        _GEN_612 = _GEN_577 & _GEN_581;
  wire        _GEN_613 = _GEN_577 & _GEN_582;
  wire        _GEN_614 = _GEN_577 & _GEN_583;
  wire        _GEN_615 = _GEN_577 & _GEN_584;
  wire        _GEN_616 = _GEN_577 & _GEN_585;
  wire        _GEN_617 = _GEN_577 & _GEN_586;
  wire        _GEN_618 = _GEN_577 & _GEN_587;
  wire        _GEN_619 = _GEN_577 & _GEN_588;
  wire        _GEN_620 = _GEN_577 & _GEN_589;
  wire        _GEN_621 = _GEN_577 & _GEN_590;
  wire        _GEN_622 = _GEN_577 & _GEN_591;
  wire        _GEN_623 = _GEN_577 & _GEN_592;
  wire        _GEN_624 = _GEN_577 & _GEN_593;
  wire        _GEN_625 = _GEN_577 & _GEN_594;
  wire        _GEN_626 = _GEN_577 & _GEN_595;
  wire        _GEN_627 = _GEN_577 & _GEN_596;
  wire        _GEN_628 = _GEN_577 & _GEN_597;
  wire        _GEN_629 = _GEN_577 & _GEN_598;
  wire        _GEN_630 = _GEN_577 & _GEN_599;
  wire        _GEN_631 = _GEN_577 & _GEN_600;
  wire        _GEN_632 = _GEN_577 & _GEN_601;
  wire        _GEN_633 = _GEN_577 & _GEN_602;
  wire        _GEN_634 = _GEN_577 & _GEN_603;
  wire        _GEN_635 = _GEN_577 & _GEN_604;
  wire        _GEN_636 = _GEN_577 & _GEN_605;
  wire        _GEN_637 = _GEN_577 & _GEN_606;
  wire        _GEN_638 = _GEN_577 & _GEN_607;
  wire        _GEN_639 = _GEN_577 & _GEN_608;
  wire        _GEN_640 = _GEN_577 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_641 = io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_642 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_643 = _GEN_642 | _GEN_609;
  wire        _GEN_644 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_645 = _GEN_644 | _GEN_610;
  wire        _GEN_646 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_647 = _GEN_646 | _GEN_611;
  wire        _GEN_648 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_649 = _GEN_648 | _GEN_612;
  wire        _GEN_650 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_651 = _GEN_650 | _GEN_613;
  wire        _GEN_652 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_653 = _GEN_652 | _GEN_614;
  wire        _GEN_654 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_655 = _GEN_654 | _GEN_615;
  wire        _GEN_656 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_657 = _GEN_656 | _GEN_616;
  wire        _GEN_658 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_659 = _GEN_658 | _GEN_617;
  wire        _GEN_660 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_661 = _GEN_660 | _GEN_618;
  wire        _GEN_662 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_663 = _GEN_662 | _GEN_619;
  wire        _GEN_664 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_665 = _GEN_664 | _GEN_620;
  wire        _GEN_666 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_667 = _GEN_666 | _GEN_621;
  wire        _GEN_668 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_669 = _GEN_668 | _GEN_622;
  wire        _GEN_670 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_671 = _GEN_670 | _GEN_623;
  wire        _GEN_672 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_673 = _GEN_672 | _GEN_624;
  wire        _GEN_674 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_675 = _GEN_674 | _GEN_625;
  wire        _GEN_676 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_677 = _GEN_676 | _GEN_626;
  wire        _GEN_678 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_679 = _GEN_678 | _GEN_627;
  wire        _GEN_680 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_681 = _GEN_680 | _GEN_628;
  wire        _GEN_682 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_683 = _GEN_682 | _GEN_629;
  wire        _GEN_684 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_685 = _GEN_684 | _GEN_630;
  wire        _GEN_686 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_687 = _GEN_686 | _GEN_631;
  wire        _GEN_688 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_689 = _GEN_688 | _GEN_632;
  wire        _GEN_690 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_691 = _GEN_690 | _GEN_633;
  wire        _GEN_692 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_693 = _GEN_692 | _GEN_634;
  wire        _GEN_694 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_695 = _GEN_694 | _GEN_635;
  wire        _GEN_696 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_697 = _GEN_696 | _GEN_636;
  wire        _GEN_698 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_699 = _GEN_698 | _GEN_637;
  wire        _GEN_700 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_701 = _GEN_700 | _GEN_638;
  wire        _GEN_702 = io_wb_resps_9_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_703 = _GEN_702 | _GEN_639;
  wire        _GEN_704 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_640;
  wire        _GEN_705 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h0;
  wire        _GEN_706 = io_lsu_clr_bsy_0_bits[6:2] == 5'h0;
  wire        _GEN_707 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1;
  wire        _GEN_708 = io_lsu_clr_bsy_0_bits[6:2] == 5'h2;
  wire        _GEN_709 = io_lsu_clr_bsy_0_bits[6:2] == 5'h3;
  wire        _GEN_710 = io_lsu_clr_bsy_0_bits[6:2] == 5'h4;
  wire        _GEN_711 = io_lsu_clr_bsy_0_bits[6:2] == 5'h5;
  wire        _GEN_712 = io_lsu_clr_bsy_0_bits[6:2] == 5'h6;
  wire        _GEN_713 = io_lsu_clr_bsy_0_bits[6:2] == 5'h7;
  wire        _GEN_714 = io_lsu_clr_bsy_0_bits[6:2] == 5'h8;
  wire        _GEN_715 = io_lsu_clr_bsy_0_bits[6:2] == 5'h9;
  wire        _GEN_716 = io_lsu_clr_bsy_0_bits[6:2] == 5'hA;
  wire        _GEN_717 = io_lsu_clr_bsy_0_bits[6:2] == 5'hB;
  wire        _GEN_718 = io_lsu_clr_bsy_0_bits[6:2] == 5'hC;
  wire        _GEN_719 = io_lsu_clr_bsy_0_bits[6:2] == 5'hD;
  wire        _GEN_720 = io_lsu_clr_bsy_0_bits[6:2] == 5'hE;
  wire        _GEN_721 = io_lsu_clr_bsy_0_bits[6:2] == 5'hF;
  wire        _GEN_722 = io_lsu_clr_bsy_0_bits[6:2] == 5'h10;
  wire        _GEN_723 = io_lsu_clr_bsy_0_bits[6:2] == 5'h11;
  wire        _GEN_724 = io_lsu_clr_bsy_0_bits[6:2] == 5'h12;
  wire        _GEN_725 = io_lsu_clr_bsy_0_bits[6:2] == 5'h13;
  wire        _GEN_726 = io_lsu_clr_bsy_0_bits[6:2] == 5'h14;
  wire        _GEN_727 = io_lsu_clr_bsy_0_bits[6:2] == 5'h15;
  wire        _GEN_728 = io_lsu_clr_bsy_0_bits[6:2] == 5'h16;
  wire        _GEN_729 = io_lsu_clr_bsy_0_bits[6:2] == 5'h17;
  wire        _GEN_730 = io_lsu_clr_bsy_0_bits[6:2] == 5'h18;
  wire        _GEN_731 = io_lsu_clr_bsy_0_bits[6:2] == 5'h19;
  wire        _GEN_732 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1A;
  wire        _GEN_733 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1B;
  wire        _GEN_734 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1C;
  wire        _GEN_735 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1D;
  wire        _GEN_736 = io_lsu_clr_bsy_0_bits[6:2] == 5'h1E;
  wire        _GEN_737 = _GEN_705 & _GEN_706;
  wire        _GEN_738 = _GEN_705 & _GEN_707;
  wire        _GEN_739 = _GEN_705 & _GEN_708;
  wire        _GEN_740 = _GEN_705 & _GEN_709;
  wire        _GEN_741 = _GEN_705 & _GEN_710;
  wire        _GEN_742 = _GEN_705 & _GEN_711;
  wire        _GEN_743 = _GEN_705 & _GEN_712;
  wire        _GEN_744 = _GEN_705 & _GEN_713;
  wire        _GEN_745 = _GEN_705 & _GEN_714;
  wire        _GEN_746 = _GEN_705 & _GEN_715;
  wire        _GEN_747 = _GEN_705 & _GEN_716;
  wire        _GEN_748 = _GEN_705 & _GEN_717;
  wire        _GEN_749 = _GEN_705 & _GEN_718;
  wire        _GEN_750 = _GEN_705 & _GEN_719;
  wire        _GEN_751 = _GEN_705 & _GEN_720;
  wire        _GEN_752 = _GEN_705 & _GEN_721;
  wire        _GEN_753 = _GEN_705 & _GEN_722;
  wire        _GEN_754 = _GEN_705 & _GEN_723;
  wire        _GEN_755 = _GEN_705 & _GEN_724;
  wire        _GEN_756 = _GEN_705 & _GEN_725;
  wire        _GEN_757 = _GEN_705 & _GEN_726;
  wire        _GEN_758 = _GEN_705 & _GEN_727;
  wire        _GEN_759 = _GEN_705 & _GEN_728;
  wire        _GEN_760 = _GEN_705 & _GEN_729;
  wire        _GEN_761 = _GEN_705 & _GEN_730;
  wire        _GEN_762 = _GEN_705 & _GEN_731;
  wire        _GEN_763 = _GEN_705 & _GEN_732;
  wire        _GEN_764 = _GEN_705 & _GEN_733;
  wire        _GEN_765 = _GEN_705 & _GEN_734;
  wire        _GEN_766 = _GEN_705 & _GEN_735;
  wire        _GEN_767 = _GEN_705 & _GEN_736;
  wire        _GEN_768 = _GEN_705 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_769 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h0;
  wire        _GEN_770 = io_lsu_clr_bsy_1_bits[6:2] == 5'h0;
  wire        _GEN_771 = _GEN_770 | _GEN_737;
  wire        _GEN_772 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1;
  wire        _GEN_773 = _GEN_772 | _GEN_738;
  wire        _GEN_774 = io_lsu_clr_bsy_1_bits[6:2] == 5'h2;
  wire        _GEN_775 = _GEN_774 | _GEN_739;
  wire        _GEN_776 = io_lsu_clr_bsy_1_bits[6:2] == 5'h3;
  wire        _GEN_777 = _GEN_776 | _GEN_740;
  wire        _GEN_778 = io_lsu_clr_bsy_1_bits[6:2] == 5'h4;
  wire        _GEN_779 = _GEN_778 | _GEN_741;
  wire        _GEN_780 = io_lsu_clr_bsy_1_bits[6:2] == 5'h5;
  wire        _GEN_781 = _GEN_780 | _GEN_742;
  wire        _GEN_782 = io_lsu_clr_bsy_1_bits[6:2] == 5'h6;
  wire        _GEN_783 = _GEN_782 | _GEN_743;
  wire        _GEN_784 = io_lsu_clr_bsy_1_bits[6:2] == 5'h7;
  wire        _GEN_785 = _GEN_784 | _GEN_744;
  wire        _GEN_786 = io_lsu_clr_bsy_1_bits[6:2] == 5'h8;
  wire        _GEN_787 = _GEN_786 | _GEN_745;
  wire        _GEN_788 = io_lsu_clr_bsy_1_bits[6:2] == 5'h9;
  wire        _GEN_789 = _GEN_788 | _GEN_746;
  wire        _GEN_790 = io_lsu_clr_bsy_1_bits[6:2] == 5'hA;
  wire        _GEN_791 = _GEN_790 | _GEN_747;
  wire        _GEN_792 = io_lsu_clr_bsy_1_bits[6:2] == 5'hB;
  wire        _GEN_793 = _GEN_792 | _GEN_748;
  wire        _GEN_794 = io_lsu_clr_bsy_1_bits[6:2] == 5'hC;
  wire        _GEN_795 = _GEN_794 | _GEN_749;
  wire        _GEN_796 = io_lsu_clr_bsy_1_bits[6:2] == 5'hD;
  wire        _GEN_797 = _GEN_796 | _GEN_750;
  wire        _GEN_798 = io_lsu_clr_bsy_1_bits[6:2] == 5'hE;
  wire        _GEN_799 = _GEN_798 | _GEN_751;
  wire        _GEN_800 = io_lsu_clr_bsy_1_bits[6:2] == 5'hF;
  wire        _GEN_801 = _GEN_800 | _GEN_752;
  wire        _GEN_802 = io_lsu_clr_bsy_1_bits[6:2] == 5'h10;
  wire        _GEN_803 = _GEN_802 | _GEN_753;
  wire        _GEN_804 = io_lsu_clr_bsy_1_bits[6:2] == 5'h11;
  wire        _GEN_805 = _GEN_804 | _GEN_754;
  wire        _GEN_806 = io_lsu_clr_bsy_1_bits[6:2] == 5'h12;
  wire        _GEN_807 = _GEN_806 | _GEN_755;
  wire        _GEN_808 = io_lsu_clr_bsy_1_bits[6:2] == 5'h13;
  wire        _GEN_809 = _GEN_808 | _GEN_756;
  wire        _GEN_810 = io_lsu_clr_bsy_1_bits[6:2] == 5'h14;
  wire        _GEN_811 = _GEN_810 | _GEN_757;
  wire        _GEN_812 = io_lsu_clr_bsy_1_bits[6:2] == 5'h15;
  wire        _GEN_813 = _GEN_812 | _GEN_758;
  wire        _GEN_814 = io_lsu_clr_bsy_1_bits[6:2] == 5'h16;
  wire        _GEN_815 = _GEN_814 | _GEN_759;
  wire        _GEN_816 = io_lsu_clr_bsy_1_bits[6:2] == 5'h17;
  wire        _GEN_817 = _GEN_816 | _GEN_760;
  wire        _GEN_818 = io_lsu_clr_bsy_1_bits[6:2] == 5'h18;
  wire        _GEN_819 = _GEN_818 | _GEN_761;
  wire        _GEN_820 = io_lsu_clr_bsy_1_bits[6:2] == 5'h19;
  wire        _GEN_821 = _GEN_820 | _GEN_762;
  wire        _GEN_822 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1A;
  wire        _GEN_823 = _GEN_822 | _GEN_763;
  wire        _GEN_824 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1B;
  wire        _GEN_825 = _GEN_824 | _GEN_764;
  wire        _GEN_826 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1C;
  wire        _GEN_827 = _GEN_826 | _GEN_765;
  wire        _GEN_828 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1D;
  wire        _GEN_829 = _GEN_828 | _GEN_766;
  wire        _GEN_830 = io_lsu_clr_bsy_1_bits[6:2] == 5'h1E;
  wire        _GEN_831 = _GEN_830 | _GEN_767;
  wire        _GEN_832 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_768;
  wire        _GEN_833 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h0;
  wire        _GEN_834 = io_lsu_clr_bsy_2_bits[6:2] == 5'h0;
  wire        _GEN_835 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1;
  wire        _GEN_836 = io_lsu_clr_bsy_2_bits[6:2] == 5'h2;
  wire        _GEN_837 = io_lsu_clr_bsy_2_bits[6:2] == 5'h3;
  wire        _GEN_838 = io_lsu_clr_bsy_2_bits[6:2] == 5'h4;
  wire        _GEN_839 = io_lsu_clr_bsy_2_bits[6:2] == 5'h5;
  wire        _GEN_840 = io_lsu_clr_bsy_2_bits[6:2] == 5'h6;
  wire        _GEN_841 = io_lsu_clr_bsy_2_bits[6:2] == 5'h7;
  wire        _GEN_842 = io_lsu_clr_bsy_2_bits[6:2] == 5'h8;
  wire        _GEN_843 = io_lsu_clr_bsy_2_bits[6:2] == 5'h9;
  wire        _GEN_844 = io_lsu_clr_bsy_2_bits[6:2] == 5'hA;
  wire        _GEN_845 = io_lsu_clr_bsy_2_bits[6:2] == 5'hB;
  wire        _GEN_846 = io_lsu_clr_bsy_2_bits[6:2] == 5'hC;
  wire        _GEN_847 = io_lsu_clr_bsy_2_bits[6:2] == 5'hD;
  wire        _GEN_848 = io_lsu_clr_bsy_2_bits[6:2] == 5'hE;
  wire        _GEN_849 = io_lsu_clr_bsy_2_bits[6:2] == 5'hF;
  wire        _GEN_850 = io_lsu_clr_bsy_2_bits[6:2] == 5'h10;
  wire        _GEN_851 = io_lsu_clr_bsy_2_bits[6:2] == 5'h11;
  wire        _GEN_852 = io_lsu_clr_bsy_2_bits[6:2] == 5'h12;
  wire        _GEN_853 = io_lsu_clr_bsy_2_bits[6:2] == 5'h13;
  wire        _GEN_854 = io_lsu_clr_bsy_2_bits[6:2] == 5'h14;
  wire        _GEN_855 = io_lsu_clr_bsy_2_bits[6:2] == 5'h15;
  wire        _GEN_856 = io_lsu_clr_bsy_2_bits[6:2] == 5'h16;
  wire        _GEN_857 = io_lsu_clr_bsy_2_bits[6:2] == 5'h17;
  wire        _GEN_858 = io_lsu_clr_bsy_2_bits[6:2] == 5'h18;
  wire        _GEN_859 = io_lsu_clr_bsy_2_bits[6:2] == 5'h19;
  wire        _GEN_860 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1A;
  wire        _GEN_861 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1B;
  wire        _GEN_862 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1C;
  wire        _GEN_863 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1D;
  wire        _GEN_864 = io_lsu_clr_bsy_2_bits[6:2] == 5'h1E;
  wire        _GEN_865 = _GEN_833 & _GEN_834;
  wire        _GEN_866 = _GEN_833 & _GEN_835;
  wire        _GEN_867 = _GEN_833 & _GEN_836;
  wire        _GEN_868 = _GEN_833 & _GEN_837;
  wire        _GEN_869 = _GEN_833 & _GEN_838;
  wire        _GEN_870 = _GEN_833 & _GEN_839;
  wire        _GEN_871 = _GEN_833 & _GEN_840;
  wire        _GEN_872 = _GEN_833 & _GEN_841;
  wire        _GEN_873 = _GEN_833 & _GEN_842;
  wire        _GEN_874 = _GEN_833 & _GEN_843;
  wire        _GEN_875 = _GEN_833 & _GEN_844;
  wire        _GEN_876 = _GEN_833 & _GEN_845;
  wire        _GEN_877 = _GEN_833 & _GEN_846;
  wire        _GEN_878 = _GEN_833 & _GEN_847;
  wire        _GEN_879 = _GEN_833 & _GEN_848;
  wire        _GEN_880 = _GEN_833 & _GEN_849;
  wire        _GEN_881 = _GEN_833 & _GEN_850;
  wire        _GEN_882 = _GEN_833 & _GEN_851;
  wire        _GEN_883 = _GEN_833 & _GEN_852;
  wire        _GEN_884 = _GEN_833 & _GEN_853;
  wire        _GEN_885 = _GEN_833 & _GEN_854;
  wire        _GEN_886 = _GEN_833 & _GEN_855;
  wire        _GEN_887 = _GEN_833 & _GEN_856;
  wire        _GEN_888 = _GEN_833 & _GEN_857;
  wire        _GEN_889 = _GEN_833 & _GEN_858;
  wire        _GEN_890 = _GEN_833 & _GEN_859;
  wire        _GEN_891 = _GEN_833 & _GEN_860;
  wire        _GEN_892 = _GEN_833 & _GEN_861;
  wire        _GEN_893 = _GEN_833 & _GEN_862;
  wire        _GEN_894 = _GEN_833 & _GEN_863;
  wire        _GEN_895 = _GEN_833 & _GEN_864;
  wire        _GEN_896 = _GEN_833 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_897 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h0;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_11 = rob_predicated__0;
      5'b00001:
        casez_tmp_11 = rob_predicated__1;
      5'b00010:
        casez_tmp_11 = rob_predicated__2;
      5'b00011:
        casez_tmp_11 = rob_predicated__3;
      5'b00100:
        casez_tmp_11 = rob_predicated__4;
      5'b00101:
        casez_tmp_11 = rob_predicated__5;
      5'b00110:
        casez_tmp_11 = rob_predicated__6;
      5'b00111:
        casez_tmp_11 = rob_predicated__7;
      5'b01000:
        casez_tmp_11 = rob_predicated__8;
      5'b01001:
        casez_tmp_11 = rob_predicated__9;
      5'b01010:
        casez_tmp_11 = rob_predicated__10;
      5'b01011:
        casez_tmp_11 = rob_predicated__11;
      5'b01100:
        casez_tmp_11 = rob_predicated__12;
      5'b01101:
        casez_tmp_11 = rob_predicated__13;
      5'b01110:
        casez_tmp_11 = rob_predicated__14;
      5'b01111:
        casez_tmp_11 = rob_predicated__15;
      5'b10000:
        casez_tmp_11 = rob_predicated__16;
      5'b10001:
        casez_tmp_11 = rob_predicated__17;
      5'b10010:
        casez_tmp_11 = rob_predicated__18;
      5'b10011:
        casez_tmp_11 = rob_predicated__19;
      5'b10100:
        casez_tmp_11 = rob_predicated__20;
      5'b10101:
        casez_tmp_11 = rob_predicated__21;
      5'b10110:
        casez_tmp_11 = rob_predicated__22;
      5'b10111:
        casez_tmp_11 = rob_predicated__23;
      5'b11000:
        casez_tmp_11 = rob_predicated__24;
      5'b11001:
        casez_tmp_11 = rob_predicated__25;
      5'b11010:
        casez_tmp_11 = rob_predicated__26;
      5'b11011:
        casez_tmp_11 = rob_predicated__27;
      5'b11100:
        casez_tmp_11 = rob_predicated__28;
      5'b11101:
        casez_tmp_11 = rob_predicated__29;
      5'b11110:
        casez_tmp_11 = rob_predicated__30;
      default:
        casez_tmp_11 = rob_predicated__31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_12 = rob_uop__0_uopc;
      5'b00001:
        casez_tmp_12 = rob_uop__1_uopc;
      5'b00010:
        casez_tmp_12 = rob_uop__2_uopc;
      5'b00011:
        casez_tmp_12 = rob_uop__3_uopc;
      5'b00100:
        casez_tmp_12 = rob_uop__4_uopc;
      5'b00101:
        casez_tmp_12 = rob_uop__5_uopc;
      5'b00110:
        casez_tmp_12 = rob_uop__6_uopc;
      5'b00111:
        casez_tmp_12 = rob_uop__7_uopc;
      5'b01000:
        casez_tmp_12 = rob_uop__8_uopc;
      5'b01001:
        casez_tmp_12 = rob_uop__9_uopc;
      5'b01010:
        casez_tmp_12 = rob_uop__10_uopc;
      5'b01011:
        casez_tmp_12 = rob_uop__11_uopc;
      5'b01100:
        casez_tmp_12 = rob_uop__12_uopc;
      5'b01101:
        casez_tmp_12 = rob_uop__13_uopc;
      5'b01110:
        casez_tmp_12 = rob_uop__14_uopc;
      5'b01111:
        casez_tmp_12 = rob_uop__15_uopc;
      5'b10000:
        casez_tmp_12 = rob_uop__16_uopc;
      5'b10001:
        casez_tmp_12 = rob_uop__17_uopc;
      5'b10010:
        casez_tmp_12 = rob_uop__18_uopc;
      5'b10011:
        casez_tmp_12 = rob_uop__19_uopc;
      5'b10100:
        casez_tmp_12 = rob_uop__20_uopc;
      5'b10101:
        casez_tmp_12 = rob_uop__21_uopc;
      5'b10110:
        casez_tmp_12 = rob_uop__22_uopc;
      5'b10111:
        casez_tmp_12 = rob_uop__23_uopc;
      5'b11000:
        casez_tmp_12 = rob_uop__24_uopc;
      5'b11001:
        casez_tmp_12 = rob_uop__25_uopc;
      5'b11010:
        casez_tmp_12 = rob_uop__26_uopc;
      5'b11011:
        casez_tmp_12 = rob_uop__27_uopc;
      5'b11100:
        casez_tmp_12 = rob_uop__28_uopc;
      5'b11101:
        casez_tmp_12 = rob_uop__29_uopc;
      5'b11110:
        casez_tmp_12 = rob_uop__30_uopc;
      default:
        casez_tmp_12 = rob_uop__31_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_13 = rob_uop__0_is_rvc;
      5'b00001:
        casez_tmp_13 = rob_uop__1_is_rvc;
      5'b00010:
        casez_tmp_13 = rob_uop__2_is_rvc;
      5'b00011:
        casez_tmp_13 = rob_uop__3_is_rvc;
      5'b00100:
        casez_tmp_13 = rob_uop__4_is_rvc;
      5'b00101:
        casez_tmp_13 = rob_uop__5_is_rvc;
      5'b00110:
        casez_tmp_13 = rob_uop__6_is_rvc;
      5'b00111:
        casez_tmp_13 = rob_uop__7_is_rvc;
      5'b01000:
        casez_tmp_13 = rob_uop__8_is_rvc;
      5'b01001:
        casez_tmp_13 = rob_uop__9_is_rvc;
      5'b01010:
        casez_tmp_13 = rob_uop__10_is_rvc;
      5'b01011:
        casez_tmp_13 = rob_uop__11_is_rvc;
      5'b01100:
        casez_tmp_13 = rob_uop__12_is_rvc;
      5'b01101:
        casez_tmp_13 = rob_uop__13_is_rvc;
      5'b01110:
        casez_tmp_13 = rob_uop__14_is_rvc;
      5'b01111:
        casez_tmp_13 = rob_uop__15_is_rvc;
      5'b10000:
        casez_tmp_13 = rob_uop__16_is_rvc;
      5'b10001:
        casez_tmp_13 = rob_uop__17_is_rvc;
      5'b10010:
        casez_tmp_13 = rob_uop__18_is_rvc;
      5'b10011:
        casez_tmp_13 = rob_uop__19_is_rvc;
      5'b10100:
        casez_tmp_13 = rob_uop__20_is_rvc;
      5'b10101:
        casez_tmp_13 = rob_uop__21_is_rvc;
      5'b10110:
        casez_tmp_13 = rob_uop__22_is_rvc;
      5'b10111:
        casez_tmp_13 = rob_uop__23_is_rvc;
      5'b11000:
        casez_tmp_13 = rob_uop__24_is_rvc;
      5'b11001:
        casez_tmp_13 = rob_uop__25_is_rvc;
      5'b11010:
        casez_tmp_13 = rob_uop__26_is_rvc;
      5'b11011:
        casez_tmp_13 = rob_uop__27_is_rvc;
      5'b11100:
        casez_tmp_13 = rob_uop__28_is_rvc;
      5'b11101:
        casez_tmp_13 = rob_uop__29_is_rvc;
      5'b11110:
        casez_tmp_13 = rob_uop__30_is_rvc;
      default:
        casez_tmp_13 = rob_uop__31_is_rvc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_14 = rob_uop__0_ftq_idx;
      5'b00001:
        casez_tmp_14 = rob_uop__1_ftq_idx;
      5'b00010:
        casez_tmp_14 = rob_uop__2_ftq_idx;
      5'b00011:
        casez_tmp_14 = rob_uop__3_ftq_idx;
      5'b00100:
        casez_tmp_14 = rob_uop__4_ftq_idx;
      5'b00101:
        casez_tmp_14 = rob_uop__5_ftq_idx;
      5'b00110:
        casez_tmp_14 = rob_uop__6_ftq_idx;
      5'b00111:
        casez_tmp_14 = rob_uop__7_ftq_idx;
      5'b01000:
        casez_tmp_14 = rob_uop__8_ftq_idx;
      5'b01001:
        casez_tmp_14 = rob_uop__9_ftq_idx;
      5'b01010:
        casez_tmp_14 = rob_uop__10_ftq_idx;
      5'b01011:
        casez_tmp_14 = rob_uop__11_ftq_idx;
      5'b01100:
        casez_tmp_14 = rob_uop__12_ftq_idx;
      5'b01101:
        casez_tmp_14 = rob_uop__13_ftq_idx;
      5'b01110:
        casez_tmp_14 = rob_uop__14_ftq_idx;
      5'b01111:
        casez_tmp_14 = rob_uop__15_ftq_idx;
      5'b10000:
        casez_tmp_14 = rob_uop__16_ftq_idx;
      5'b10001:
        casez_tmp_14 = rob_uop__17_ftq_idx;
      5'b10010:
        casez_tmp_14 = rob_uop__18_ftq_idx;
      5'b10011:
        casez_tmp_14 = rob_uop__19_ftq_idx;
      5'b10100:
        casez_tmp_14 = rob_uop__20_ftq_idx;
      5'b10101:
        casez_tmp_14 = rob_uop__21_ftq_idx;
      5'b10110:
        casez_tmp_14 = rob_uop__22_ftq_idx;
      5'b10111:
        casez_tmp_14 = rob_uop__23_ftq_idx;
      5'b11000:
        casez_tmp_14 = rob_uop__24_ftq_idx;
      5'b11001:
        casez_tmp_14 = rob_uop__25_ftq_idx;
      5'b11010:
        casez_tmp_14 = rob_uop__26_ftq_idx;
      5'b11011:
        casez_tmp_14 = rob_uop__27_ftq_idx;
      5'b11100:
        casez_tmp_14 = rob_uop__28_ftq_idx;
      5'b11101:
        casez_tmp_14 = rob_uop__29_ftq_idx;
      5'b11110:
        casez_tmp_14 = rob_uop__30_ftq_idx;
      default:
        casez_tmp_14 = rob_uop__31_ftq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_15 = rob_uop__0_edge_inst;
      5'b00001:
        casez_tmp_15 = rob_uop__1_edge_inst;
      5'b00010:
        casez_tmp_15 = rob_uop__2_edge_inst;
      5'b00011:
        casez_tmp_15 = rob_uop__3_edge_inst;
      5'b00100:
        casez_tmp_15 = rob_uop__4_edge_inst;
      5'b00101:
        casez_tmp_15 = rob_uop__5_edge_inst;
      5'b00110:
        casez_tmp_15 = rob_uop__6_edge_inst;
      5'b00111:
        casez_tmp_15 = rob_uop__7_edge_inst;
      5'b01000:
        casez_tmp_15 = rob_uop__8_edge_inst;
      5'b01001:
        casez_tmp_15 = rob_uop__9_edge_inst;
      5'b01010:
        casez_tmp_15 = rob_uop__10_edge_inst;
      5'b01011:
        casez_tmp_15 = rob_uop__11_edge_inst;
      5'b01100:
        casez_tmp_15 = rob_uop__12_edge_inst;
      5'b01101:
        casez_tmp_15 = rob_uop__13_edge_inst;
      5'b01110:
        casez_tmp_15 = rob_uop__14_edge_inst;
      5'b01111:
        casez_tmp_15 = rob_uop__15_edge_inst;
      5'b10000:
        casez_tmp_15 = rob_uop__16_edge_inst;
      5'b10001:
        casez_tmp_15 = rob_uop__17_edge_inst;
      5'b10010:
        casez_tmp_15 = rob_uop__18_edge_inst;
      5'b10011:
        casez_tmp_15 = rob_uop__19_edge_inst;
      5'b10100:
        casez_tmp_15 = rob_uop__20_edge_inst;
      5'b10101:
        casez_tmp_15 = rob_uop__21_edge_inst;
      5'b10110:
        casez_tmp_15 = rob_uop__22_edge_inst;
      5'b10111:
        casez_tmp_15 = rob_uop__23_edge_inst;
      5'b11000:
        casez_tmp_15 = rob_uop__24_edge_inst;
      5'b11001:
        casez_tmp_15 = rob_uop__25_edge_inst;
      5'b11010:
        casez_tmp_15 = rob_uop__26_edge_inst;
      5'b11011:
        casez_tmp_15 = rob_uop__27_edge_inst;
      5'b11100:
        casez_tmp_15 = rob_uop__28_edge_inst;
      5'b11101:
        casez_tmp_15 = rob_uop__29_edge_inst;
      5'b11110:
        casez_tmp_15 = rob_uop__30_edge_inst;
      default:
        casez_tmp_15 = rob_uop__31_edge_inst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_16 = rob_uop__0_pc_lob;
      5'b00001:
        casez_tmp_16 = rob_uop__1_pc_lob;
      5'b00010:
        casez_tmp_16 = rob_uop__2_pc_lob;
      5'b00011:
        casez_tmp_16 = rob_uop__3_pc_lob;
      5'b00100:
        casez_tmp_16 = rob_uop__4_pc_lob;
      5'b00101:
        casez_tmp_16 = rob_uop__5_pc_lob;
      5'b00110:
        casez_tmp_16 = rob_uop__6_pc_lob;
      5'b00111:
        casez_tmp_16 = rob_uop__7_pc_lob;
      5'b01000:
        casez_tmp_16 = rob_uop__8_pc_lob;
      5'b01001:
        casez_tmp_16 = rob_uop__9_pc_lob;
      5'b01010:
        casez_tmp_16 = rob_uop__10_pc_lob;
      5'b01011:
        casez_tmp_16 = rob_uop__11_pc_lob;
      5'b01100:
        casez_tmp_16 = rob_uop__12_pc_lob;
      5'b01101:
        casez_tmp_16 = rob_uop__13_pc_lob;
      5'b01110:
        casez_tmp_16 = rob_uop__14_pc_lob;
      5'b01111:
        casez_tmp_16 = rob_uop__15_pc_lob;
      5'b10000:
        casez_tmp_16 = rob_uop__16_pc_lob;
      5'b10001:
        casez_tmp_16 = rob_uop__17_pc_lob;
      5'b10010:
        casez_tmp_16 = rob_uop__18_pc_lob;
      5'b10011:
        casez_tmp_16 = rob_uop__19_pc_lob;
      5'b10100:
        casez_tmp_16 = rob_uop__20_pc_lob;
      5'b10101:
        casez_tmp_16 = rob_uop__21_pc_lob;
      5'b10110:
        casez_tmp_16 = rob_uop__22_pc_lob;
      5'b10111:
        casez_tmp_16 = rob_uop__23_pc_lob;
      5'b11000:
        casez_tmp_16 = rob_uop__24_pc_lob;
      5'b11001:
        casez_tmp_16 = rob_uop__25_pc_lob;
      5'b11010:
        casez_tmp_16 = rob_uop__26_pc_lob;
      5'b11011:
        casez_tmp_16 = rob_uop__27_pc_lob;
      5'b11100:
        casez_tmp_16 = rob_uop__28_pc_lob;
      5'b11101:
        casez_tmp_16 = rob_uop__29_pc_lob;
      5'b11110:
        casez_tmp_16 = rob_uop__30_pc_lob;
      default:
        casez_tmp_16 = rob_uop__31_pc_lob;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_17 = rob_uop__0_pdst;
      5'b00001:
        casez_tmp_17 = rob_uop__1_pdst;
      5'b00010:
        casez_tmp_17 = rob_uop__2_pdst;
      5'b00011:
        casez_tmp_17 = rob_uop__3_pdst;
      5'b00100:
        casez_tmp_17 = rob_uop__4_pdst;
      5'b00101:
        casez_tmp_17 = rob_uop__5_pdst;
      5'b00110:
        casez_tmp_17 = rob_uop__6_pdst;
      5'b00111:
        casez_tmp_17 = rob_uop__7_pdst;
      5'b01000:
        casez_tmp_17 = rob_uop__8_pdst;
      5'b01001:
        casez_tmp_17 = rob_uop__9_pdst;
      5'b01010:
        casez_tmp_17 = rob_uop__10_pdst;
      5'b01011:
        casez_tmp_17 = rob_uop__11_pdst;
      5'b01100:
        casez_tmp_17 = rob_uop__12_pdst;
      5'b01101:
        casez_tmp_17 = rob_uop__13_pdst;
      5'b01110:
        casez_tmp_17 = rob_uop__14_pdst;
      5'b01111:
        casez_tmp_17 = rob_uop__15_pdst;
      5'b10000:
        casez_tmp_17 = rob_uop__16_pdst;
      5'b10001:
        casez_tmp_17 = rob_uop__17_pdst;
      5'b10010:
        casez_tmp_17 = rob_uop__18_pdst;
      5'b10011:
        casez_tmp_17 = rob_uop__19_pdst;
      5'b10100:
        casez_tmp_17 = rob_uop__20_pdst;
      5'b10101:
        casez_tmp_17 = rob_uop__21_pdst;
      5'b10110:
        casez_tmp_17 = rob_uop__22_pdst;
      5'b10111:
        casez_tmp_17 = rob_uop__23_pdst;
      5'b11000:
        casez_tmp_17 = rob_uop__24_pdst;
      5'b11001:
        casez_tmp_17 = rob_uop__25_pdst;
      5'b11010:
        casez_tmp_17 = rob_uop__26_pdst;
      5'b11011:
        casez_tmp_17 = rob_uop__27_pdst;
      5'b11100:
        casez_tmp_17 = rob_uop__28_pdst;
      5'b11101:
        casez_tmp_17 = rob_uop__29_pdst;
      5'b11110:
        casez_tmp_17 = rob_uop__30_pdst;
      default:
        casez_tmp_17 = rob_uop__31_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_18 = rob_uop__0_stale_pdst;
      5'b00001:
        casez_tmp_18 = rob_uop__1_stale_pdst;
      5'b00010:
        casez_tmp_18 = rob_uop__2_stale_pdst;
      5'b00011:
        casez_tmp_18 = rob_uop__3_stale_pdst;
      5'b00100:
        casez_tmp_18 = rob_uop__4_stale_pdst;
      5'b00101:
        casez_tmp_18 = rob_uop__5_stale_pdst;
      5'b00110:
        casez_tmp_18 = rob_uop__6_stale_pdst;
      5'b00111:
        casez_tmp_18 = rob_uop__7_stale_pdst;
      5'b01000:
        casez_tmp_18 = rob_uop__8_stale_pdst;
      5'b01001:
        casez_tmp_18 = rob_uop__9_stale_pdst;
      5'b01010:
        casez_tmp_18 = rob_uop__10_stale_pdst;
      5'b01011:
        casez_tmp_18 = rob_uop__11_stale_pdst;
      5'b01100:
        casez_tmp_18 = rob_uop__12_stale_pdst;
      5'b01101:
        casez_tmp_18 = rob_uop__13_stale_pdst;
      5'b01110:
        casez_tmp_18 = rob_uop__14_stale_pdst;
      5'b01111:
        casez_tmp_18 = rob_uop__15_stale_pdst;
      5'b10000:
        casez_tmp_18 = rob_uop__16_stale_pdst;
      5'b10001:
        casez_tmp_18 = rob_uop__17_stale_pdst;
      5'b10010:
        casez_tmp_18 = rob_uop__18_stale_pdst;
      5'b10011:
        casez_tmp_18 = rob_uop__19_stale_pdst;
      5'b10100:
        casez_tmp_18 = rob_uop__20_stale_pdst;
      5'b10101:
        casez_tmp_18 = rob_uop__21_stale_pdst;
      5'b10110:
        casez_tmp_18 = rob_uop__22_stale_pdst;
      5'b10111:
        casez_tmp_18 = rob_uop__23_stale_pdst;
      5'b11000:
        casez_tmp_18 = rob_uop__24_stale_pdst;
      5'b11001:
        casez_tmp_18 = rob_uop__25_stale_pdst;
      5'b11010:
        casez_tmp_18 = rob_uop__26_stale_pdst;
      5'b11011:
        casez_tmp_18 = rob_uop__27_stale_pdst;
      5'b11100:
        casez_tmp_18 = rob_uop__28_stale_pdst;
      5'b11101:
        casez_tmp_18 = rob_uop__29_stale_pdst;
      5'b11110:
        casez_tmp_18 = rob_uop__30_stale_pdst;
      default:
        casez_tmp_18 = rob_uop__31_stale_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_19 = rob_uop__0_is_fencei;
      5'b00001:
        casez_tmp_19 = rob_uop__1_is_fencei;
      5'b00010:
        casez_tmp_19 = rob_uop__2_is_fencei;
      5'b00011:
        casez_tmp_19 = rob_uop__3_is_fencei;
      5'b00100:
        casez_tmp_19 = rob_uop__4_is_fencei;
      5'b00101:
        casez_tmp_19 = rob_uop__5_is_fencei;
      5'b00110:
        casez_tmp_19 = rob_uop__6_is_fencei;
      5'b00111:
        casez_tmp_19 = rob_uop__7_is_fencei;
      5'b01000:
        casez_tmp_19 = rob_uop__8_is_fencei;
      5'b01001:
        casez_tmp_19 = rob_uop__9_is_fencei;
      5'b01010:
        casez_tmp_19 = rob_uop__10_is_fencei;
      5'b01011:
        casez_tmp_19 = rob_uop__11_is_fencei;
      5'b01100:
        casez_tmp_19 = rob_uop__12_is_fencei;
      5'b01101:
        casez_tmp_19 = rob_uop__13_is_fencei;
      5'b01110:
        casez_tmp_19 = rob_uop__14_is_fencei;
      5'b01111:
        casez_tmp_19 = rob_uop__15_is_fencei;
      5'b10000:
        casez_tmp_19 = rob_uop__16_is_fencei;
      5'b10001:
        casez_tmp_19 = rob_uop__17_is_fencei;
      5'b10010:
        casez_tmp_19 = rob_uop__18_is_fencei;
      5'b10011:
        casez_tmp_19 = rob_uop__19_is_fencei;
      5'b10100:
        casez_tmp_19 = rob_uop__20_is_fencei;
      5'b10101:
        casez_tmp_19 = rob_uop__21_is_fencei;
      5'b10110:
        casez_tmp_19 = rob_uop__22_is_fencei;
      5'b10111:
        casez_tmp_19 = rob_uop__23_is_fencei;
      5'b11000:
        casez_tmp_19 = rob_uop__24_is_fencei;
      5'b11001:
        casez_tmp_19 = rob_uop__25_is_fencei;
      5'b11010:
        casez_tmp_19 = rob_uop__26_is_fencei;
      5'b11011:
        casez_tmp_19 = rob_uop__27_is_fencei;
      5'b11100:
        casez_tmp_19 = rob_uop__28_is_fencei;
      5'b11101:
        casez_tmp_19 = rob_uop__29_is_fencei;
      5'b11110:
        casez_tmp_19 = rob_uop__30_is_fencei;
      default:
        casez_tmp_19 = rob_uop__31_is_fencei;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_20 = rob_uop__0_uses_ldq;
      5'b00001:
        casez_tmp_20 = rob_uop__1_uses_ldq;
      5'b00010:
        casez_tmp_20 = rob_uop__2_uses_ldq;
      5'b00011:
        casez_tmp_20 = rob_uop__3_uses_ldq;
      5'b00100:
        casez_tmp_20 = rob_uop__4_uses_ldq;
      5'b00101:
        casez_tmp_20 = rob_uop__5_uses_ldq;
      5'b00110:
        casez_tmp_20 = rob_uop__6_uses_ldq;
      5'b00111:
        casez_tmp_20 = rob_uop__7_uses_ldq;
      5'b01000:
        casez_tmp_20 = rob_uop__8_uses_ldq;
      5'b01001:
        casez_tmp_20 = rob_uop__9_uses_ldq;
      5'b01010:
        casez_tmp_20 = rob_uop__10_uses_ldq;
      5'b01011:
        casez_tmp_20 = rob_uop__11_uses_ldq;
      5'b01100:
        casez_tmp_20 = rob_uop__12_uses_ldq;
      5'b01101:
        casez_tmp_20 = rob_uop__13_uses_ldq;
      5'b01110:
        casez_tmp_20 = rob_uop__14_uses_ldq;
      5'b01111:
        casez_tmp_20 = rob_uop__15_uses_ldq;
      5'b10000:
        casez_tmp_20 = rob_uop__16_uses_ldq;
      5'b10001:
        casez_tmp_20 = rob_uop__17_uses_ldq;
      5'b10010:
        casez_tmp_20 = rob_uop__18_uses_ldq;
      5'b10011:
        casez_tmp_20 = rob_uop__19_uses_ldq;
      5'b10100:
        casez_tmp_20 = rob_uop__20_uses_ldq;
      5'b10101:
        casez_tmp_20 = rob_uop__21_uses_ldq;
      5'b10110:
        casez_tmp_20 = rob_uop__22_uses_ldq;
      5'b10111:
        casez_tmp_20 = rob_uop__23_uses_ldq;
      5'b11000:
        casez_tmp_20 = rob_uop__24_uses_ldq;
      5'b11001:
        casez_tmp_20 = rob_uop__25_uses_ldq;
      5'b11010:
        casez_tmp_20 = rob_uop__26_uses_ldq;
      5'b11011:
        casez_tmp_20 = rob_uop__27_uses_ldq;
      5'b11100:
        casez_tmp_20 = rob_uop__28_uses_ldq;
      5'b11101:
        casez_tmp_20 = rob_uop__29_uses_ldq;
      5'b11110:
        casez_tmp_20 = rob_uop__30_uses_ldq;
      default:
        casez_tmp_20 = rob_uop__31_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_21 = rob_uop__0_uses_stq;
      5'b00001:
        casez_tmp_21 = rob_uop__1_uses_stq;
      5'b00010:
        casez_tmp_21 = rob_uop__2_uses_stq;
      5'b00011:
        casez_tmp_21 = rob_uop__3_uses_stq;
      5'b00100:
        casez_tmp_21 = rob_uop__4_uses_stq;
      5'b00101:
        casez_tmp_21 = rob_uop__5_uses_stq;
      5'b00110:
        casez_tmp_21 = rob_uop__6_uses_stq;
      5'b00111:
        casez_tmp_21 = rob_uop__7_uses_stq;
      5'b01000:
        casez_tmp_21 = rob_uop__8_uses_stq;
      5'b01001:
        casez_tmp_21 = rob_uop__9_uses_stq;
      5'b01010:
        casez_tmp_21 = rob_uop__10_uses_stq;
      5'b01011:
        casez_tmp_21 = rob_uop__11_uses_stq;
      5'b01100:
        casez_tmp_21 = rob_uop__12_uses_stq;
      5'b01101:
        casez_tmp_21 = rob_uop__13_uses_stq;
      5'b01110:
        casez_tmp_21 = rob_uop__14_uses_stq;
      5'b01111:
        casez_tmp_21 = rob_uop__15_uses_stq;
      5'b10000:
        casez_tmp_21 = rob_uop__16_uses_stq;
      5'b10001:
        casez_tmp_21 = rob_uop__17_uses_stq;
      5'b10010:
        casez_tmp_21 = rob_uop__18_uses_stq;
      5'b10011:
        casez_tmp_21 = rob_uop__19_uses_stq;
      5'b10100:
        casez_tmp_21 = rob_uop__20_uses_stq;
      5'b10101:
        casez_tmp_21 = rob_uop__21_uses_stq;
      5'b10110:
        casez_tmp_21 = rob_uop__22_uses_stq;
      5'b10111:
        casez_tmp_21 = rob_uop__23_uses_stq;
      5'b11000:
        casez_tmp_21 = rob_uop__24_uses_stq;
      5'b11001:
        casez_tmp_21 = rob_uop__25_uses_stq;
      5'b11010:
        casez_tmp_21 = rob_uop__26_uses_stq;
      5'b11011:
        casez_tmp_21 = rob_uop__27_uses_stq;
      5'b11100:
        casez_tmp_21 = rob_uop__28_uses_stq;
      5'b11101:
        casez_tmp_21 = rob_uop__29_uses_stq;
      5'b11110:
        casez_tmp_21 = rob_uop__30_uses_stq;
      default:
        casez_tmp_21 = rob_uop__31_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_22 = rob_uop__0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_22 = rob_uop__1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_22 = rob_uop__2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_22 = rob_uop__3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_22 = rob_uop__4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_22 = rob_uop__5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_22 = rob_uop__6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_22 = rob_uop__7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_22 = rob_uop__8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_22 = rob_uop__9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_22 = rob_uop__10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_22 = rob_uop__11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_22 = rob_uop__12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_22 = rob_uop__13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_22 = rob_uop__14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_22 = rob_uop__15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_22 = rob_uop__16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_22 = rob_uop__17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_22 = rob_uop__18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_22 = rob_uop__19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_22 = rob_uop__20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_22 = rob_uop__21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_22 = rob_uop__22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_22 = rob_uop__23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_22 = rob_uop__24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_22 = rob_uop__25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_22 = rob_uop__26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_22 = rob_uop__27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_22 = rob_uop__28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_22 = rob_uop__29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_22 = rob_uop__30_is_sys_pc2epc;
      default:
        casez_tmp_22 = rob_uop__31_is_sys_pc2epc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_23 = rob_uop__0_flush_on_commit;
      5'b00001:
        casez_tmp_23 = rob_uop__1_flush_on_commit;
      5'b00010:
        casez_tmp_23 = rob_uop__2_flush_on_commit;
      5'b00011:
        casez_tmp_23 = rob_uop__3_flush_on_commit;
      5'b00100:
        casez_tmp_23 = rob_uop__4_flush_on_commit;
      5'b00101:
        casez_tmp_23 = rob_uop__5_flush_on_commit;
      5'b00110:
        casez_tmp_23 = rob_uop__6_flush_on_commit;
      5'b00111:
        casez_tmp_23 = rob_uop__7_flush_on_commit;
      5'b01000:
        casez_tmp_23 = rob_uop__8_flush_on_commit;
      5'b01001:
        casez_tmp_23 = rob_uop__9_flush_on_commit;
      5'b01010:
        casez_tmp_23 = rob_uop__10_flush_on_commit;
      5'b01011:
        casez_tmp_23 = rob_uop__11_flush_on_commit;
      5'b01100:
        casez_tmp_23 = rob_uop__12_flush_on_commit;
      5'b01101:
        casez_tmp_23 = rob_uop__13_flush_on_commit;
      5'b01110:
        casez_tmp_23 = rob_uop__14_flush_on_commit;
      5'b01111:
        casez_tmp_23 = rob_uop__15_flush_on_commit;
      5'b10000:
        casez_tmp_23 = rob_uop__16_flush_on_commit;
      5'b10001:
        casez_tmp_23 = rob_uop__17_flush_on_commit;
      5'b10010:
        casez_tmp_23 = rob_uop__18_flush_on_commit;
      5'b10011:
        casez_tmp_23 = rob_uop__19_flush_on_commit;
      5'b10100:
        casez_tmp_23 = rob_uop__20_flush_on_commit;
      5'b10101:
        casez_tmp_23 = rob_uop__21_flush_on_commit;
      5'b10110:
        casez_tmp_23 = rob_uop__22_flush_on_commit;
      5'b10111:
        casez_tmp_23 = rob_uop__23_flush_on_commit;
      5'b11000:
        casez_tmp_23 = rob_uop__24_flush_on_commit;
      5'b11001:
        casez_tmp_23 = rob_uop__25_flush_on_commit;
      5'b11010:
        casez_tmp_23 = rob_uop__26_flush_on_commit;
      5'b11011:
        casez_tmp_23 = rob_uop__27_flush_on_commit;
      5'b11100:
        casez_tmp_23 = rob_uop__28_flush_on_commit;
      5'b11101:
        casez_tmp_23 = rob_uop__29_flush_on_commit;
      5'b11110:
        casez_tmp_23 = rob_uop__30_flush_on_commit;
      default:
        casez_tmp_23 = rob_uop__31_flush_on_commit;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_24 = rob_uop__0_ldst;
      5'b00001:
        casez_tmp_24 = rob_uop__1_ldst;
      5'b00010:
        casez_tmp_24 = rob_uop__2_ldst;
      5'b00011:
        casez_tmp_24 = rob_uop__3_ldst;
      5'b00100:
        casez_tmp_24 = rob_uop__4_ldst;
      5'b00101:
        casez_tmp_24 = rob_uop__5_ldst;
      5'b00110:
        casez_tmp_24 = rob_uop__6_ldst;
      5'b00111:
        casez_tmp_24 = rob_uop__7_ldst;
      5'b01000:
        casez_tmp_24 = rob_uop__8_ldst;
      5'b01001:
        casez_tmp_24 = rob_uop__9_ldst;
      5'b01010:
        casez_tmp_24 = rob_uop__10_ldst;
      5'b01011:
        casez_tmp_24 = rob_uop__11_ldst;
      5'b01100:
        casez_tmp_24 = rob_uop__12_ldst;
      5'b01101:
        casez_tmp_24 = rob_uop__13_ldst;
      5'b01110:
        casez_tmp_24 = rob_uop__14_ldst;
      5'b01111:
        casez_tmp_24 = rob_uop__15_ldst;
      5'b10000:
        casez_tmp_24 = rob_uop__16_ldst;
      5'b10001:
        casez_tmp_24 = rob_uop__17_ldst;
      5'b10010:
        casez_tmp_24 = rob_uop__18_ldst;
      5'b10011:
        casez_tmp_24 = rob_uop__19_ldst;
      5'b10100:
        casez_tmp_24 = rob_uop__20_ldst;
      5'b10101:
        casez_tmp_24 = rob_uop__21_ldst;
      5'b10110:
        casez_tmp_24 = rob_uop__22_ldst;
      5'b10111:
        casez_tmp_24 = rob_uop__23_ldst;
      5'b11000:
        casez_tmp_24 = rob_uop__24_ldst;
      5'b11001:
        casez_tmp_24 = rob_uop__25_ldst;
      5'b11010:
        casez_tmp_24 = rob_uop__26_ldst;
      5'b11011:
        casez_tmp_24 = rob_uop__27_ldst;
      5'b11100:
        casez_tmp_24 = rob_uop__28_ldst;
      5'b11101:
        casez_tmp_24 = rob_uop__29_ldst;
      5'b11110:
        casez_tmp_24 = rob_uop__30_ldst;
      default:
        casez_tmp_24 = rob_uop__31_ldst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_25 = rob_uop__0_ldst_val;
      5'b00001:
        casez_tmp_25 = rob_uop__1_ldst_val;
      5'b00010:
        casez_tmp_25 = rob_uop__2_ldst_val;
      5'b00011:
        casez_tmp_25 = rob_uop__3_ldst_val;
      5'b00100:
        casez_tmp_25 = rob_uop__4_ldst_val;
      5'b00101:
        casez_tmp_25 = rob_uop__5_ldst_val;
      5'b00110:
        casez_tmp_25 = rob_uop__6_ldst_val;
      5'b00111:
        casez_tmp_25 = rob_uop__7_ldst_val;
      5'b01000:
        casez_tmp_25 = rob_uop__8_ldst_val;
      5'b01001:
        casez_tmp_25 = rob_uop__9_ldst_val;
      5'b01010:
        casez_tmp_25 = rob_uop__10_ldst_val;
      5'b01011:
        casez_tmp_25 = rob_uop__11_ldst_val;
      5'b01100:
        casez_tmp_25 = rob_uop__12_ldst_val;
      5'b01101:
        casez_tmp_25 = rob_uop__13_ldst_val;
      5'b01110:
        casez_tmp_25 = rob_uop__14_ldst_val;
      5'b01111:
        casez_tmp_25 = rob_uop__15_ldst_val;
      5'b10000:
        casez_tmp_25 = rob_uop__16_ldst_val;
      5'b10001:
        casez_tmp_25 = rob_uop__17_ldst_val;
      5'b10010:
        casez_tmp_25 = rob_uop__18_ldst_val;
      5'b10011:
        casez_tmp_25 = rob_uop__19_ldst_val;
      5'b10100:
        casez_tmp_25 = rob_uop__20_ldst_val;
      5'b10101:
        casez_tmp_25 = rob_uop__21_ldst_val;
      5'b10110:
        casez_tmp_25 = rob_uop__22_ldst_val;
      5'b10111:
        casez_tmp_25 = rob_uop__23_ldst_val;
      5'b11000:
        casez_tmp_25 = rob_uop__24_ldst_val;
      5'b11001:
        casez_tmp_25 = rob_uop__25_ldst_val;
      5'b11010:
        casez_tmp_25 = rob_uop__26_ldst_val;
      5'b11011:
        casez_tmp_25 = rob_uop__27_ldst_val;
      5'b11100:
        casez_tmp_25 = rob_uop__28_ldst_val;
      5'b11101:
        casez_tmp_25 = rob_uop__29_ldst_val;
      5'b11110:
        casez_tmp_25 = rob_uop__30_ldst_val;
      default:
        casez_tmp_25 = rob_uop__31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_26 = rob_uop__0_dst_rtype;
      5'b00001:
        casez_tmp_26 = rob_uop__1_dst_rtype;
      5'b00010:
        casez_tmp_26 = rob_uop__2_dst_rtype;
      5'b00011:
        casez_tmp_26 = rob_uop__3_dst_rtype;
      5'b00100:
        casez_tmp_26 = rob_uop__4_dst_rtype;
      5'b00101:
        casez_tmp_26 = rob_uop__5_dst_rtype;
      5'b00110:
        casez_tmp_26 = rob_uop__6_dst_rtype;
      5'b00111:
        casez_tmp_26 = rob_uop__7_dst_rtype;
      5'b01000:
        casez_tmp_26 = rob_uop__8_dst_rtype;
      5'b01001:
        casez_tmp_26 = rob_uop__9_dst_rtype;
      5'b01010:
        casez_tmp_26 = rob_uop__10_dst_rtype;
      5'b01011:
        casez_tmp_26 = rob_uop__11_dst_rtype;
      5'b01100:
        casez_tmp_26 = rob_uop__12_dst_rtype;
      5'b01101:
        casez_tmp_26 = rob_uop__13_dst_rtype;
      5'b01110:
        casez_tmp_26 = rob_uop__14_dst_rtype;
      5'b01111:
        casez_tmp_26 = rob_uop__15_dst_rtype;
      5'b10000:
        casez_tmp_26 = rob_uop__16_dst_rtype;
      5'b10001:
        casez_tmp_26 = rob_uop__17_dst_rtype;
      5'b10010:
        casez_tmp_26 = rob_uop__18_dst_rtype;
      5'b10011:
        casez_tmp_26 = rob_uop__19_dst_rtype;
      5'b10100:
        casez_tmp_26 = rob_uop__20_dst_rtype;
      5'b10101:
        casez_tmp_26 = rob_uop__21_dst_rtype;
      5'b10110:
        casez_tmp_26 = rob_uop__22_dst_rtype;
      5'b10111:
        casez_tmp_26 = rob_uop__23_dst_rtype;
      5'b11000:
        casez_tmp_26 = rob_uop__24_dst_rtype;
      5'b11001:
        casez_tmp_26 = rob_uop__25_dst_rtype;
      5'b11010:
        casez_tmp_26 = rob_uop__26_dst_rtype;
      5'b11011:
        casez_tmp_26 = rob_uop__27_dst_rtype;
      5'b11100:
        casez_tmp_26 = rob_uop__28_dst_rtype;
      5'b11101:
        casez_tmp_26 = rob_uop__29_dst_rtype;
      5'b11110:
        casez_tmp_26 = rob_uop__30_dst_rtype;
      default:
        casez_tmp_26 = rob_uop__31_dst_rtype;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_27 = rob_uop__0_fp_val;
      5'b00001:
        casez_tmp_27 = rob_uop__1_fp_val;
      5'b00010:
        casez_tmp_27 = rob_uop__2_fp_val;
      5'b00011:
        casez_tmp_27 = rob_uop__3_fp_val;
      5'b00100:
        casez_tmp_27 = rob_uop__4_fp_val;
      5'b00101:
        casez_tmp_27 = rob_uop__5_fp_val;
      5'b00110:
        casez_tmp_27 = rob_uop__6_fp_val;
      5'b00111:
        casez_tmp_27 = rob_uop__7_fp_val;
      5'b01000:
        casez_tmp_27 = rob_uop__8_fp_val;
      5'b01001:
        casez_tmp_27 = rob_uop__9_fp_val;
      5'b01010:
        casez_tmp_27 = rob_uop__10_fp_val;
      5'b01011:
        casez_tmp_27 = rob_uop__11_fp_val;
      5'b01100:
        casez_tmp_27 = rob_uop__12_fp_val;
      5'b01101:
        casez_tmp_27 = rob_uop__13_fp_val;
      5'b01110:
        casez_tmp_27 = rob_uop__14_fp_val;
      5'b01111:
        casez_tmp_27 = rob_uop__15_fp_val;
      5'b10000:
        casez_tmp_27 = rob_uop__16_fp_val;
      5'b10001:
        casez_tmp_27 = rob_uop__17_fp_val;
      5'b10010:
        casez_tmp_27 = rob_uop__18_fp_val;
      5'b10011:
        casez_tmp_27 = rob_uop__19_fp_val;
      5'b10100:
        casez_tmp_27 = rob_uop__20_fp_val;
      5'b10101:
        casez_tmp_27 = rob_uop__21_fp_val;
      5'b10110:
        casez_tmp_27 = rob_uop__22_fp_val;
      5'b10111:
        casez_tmp_27 = rob_uop__23_fp_val;
      5'b11000:
        casez_tmp_27 = rob_uop__24_fp_val;
      5'b11001:
        casez_tmp_27 = rob_uop__25_fp_val;
      5'b11010:
        casez_tmp_27 = rob_uop__26_fp_val;
      5'b11011:
        casez_tmp_27 = rob_uop__27_fp_val;
      5'b11100:
        casez_tmp_27 = rob_uop__28_fp_val;
      5'b11101:
        casez_tmp_27 = rob_uop__29_fp_val;
      5'b11110:
        casez_tmp_27 = rob_uop__30_fp_val;
      default:
        casez_tmp_27 = rob_uop__31_fp_val;
    endcase
  end // always @(*)
  wire        _full_T = rob_tail == rob_head;
  wire        full = _full_T & maybe_full;
  wire        rbk_row = _io_commit_rollback_T_3 & ~full;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_28 = rob_val__0;
      5'b00001:
        casez_tmp_28 = rob_val__1;
      5'b00010:
        casez_tmp_28 = rob_val__2;
      5'b00011:
        casez_tmp_28 = rob_val__3;
      5'b00100:
        casez_tmp_28 = rob_val__4;
      5'b00101:
        casez_tmp_28 = rob_val__5;
      5'b00110:
        casez_tmp_28 = rob_val__6;
      5'b00111:
        casez_tmp_28 = rob_val__7;
      5'b01000:
        casez_tmp_28 = rob_val__8;
      5'b01001:
        casez_tmp_28 = rob_val__9;
      5'b01010:
        casez_tmp_28 = rob_val__10;
      5'b01011:
        casez_tmp_28 = rob_val__11;
      5'b01100:
        casez_tmp_28 = rob_val__12;
      5'b01101:
        casez_tmp_28 = rob_val__13;
      5'b01110:
        casez_tmp_28 = rob_val__14;
      5'b01111:
        casez_tmp_28 = rob_val__15;
      5'b10000:
        casez_tmp_28 = rob_val__16;
      5'b10001:
        casez_tmp_28 = rob_val__17;
      5'b10010:
        casez_tmp_28 = rob_val__18;
      5'b10011:
        casez_tmp_28 = rob_val__19;
      5'b10100:
        casez_tmp_28 = rob_val__20;
      5'b10101:
        casez_tmp_28 = rob_val__21;
      5'b10110:
        casez_tmp_28 = rob_val__22;
      5'b10111:
        casez_tmp_28 = rob_val__23;
      5'b11000:
        casez_tmp_28 = rob_val__24;
      5'b11001:
        casez_tmp_28 = rob_val__25;
      5'b11010:
        casez_tmp_28 = rob_val__26;
      5'b11011:
        casez_tmp_28 = rob_val__27;
      5'b11100:
        casez_tmp_28 = rob_val__28;
      5'b11101:
        casez_tmp_28 = rob_val__29;
      5'b11110:
        casez_tmp_28 = rob_val__30;
      default:
        casez_tmp_28 = rob_val__31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_0_output = rbk_row & casez_tmp_28;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_29 = rob_fflags_0_0;
      5'b00001:
        casez_tmp_29 = rob_fflags_0_1;
      5'b00010:
        casez_tmp_29 = rob_fflags_0_2;
      5'b00011:
        casez_tmp_29 = rob_fflags_0_3;
      5'b00100:
        casez_tmp_29 = rob_fflags_0_4;
      5'b00101:
        casez_tmp_29 = rob_fflags_0_5;
      5'b00110:
        casez_tmp_29 = rob_fflags_0_6;
      5'b00111:
        casez_tmp_29 = rob_fflags_0_7;
      5'b01000:
        casez_tmp_29 = rob_fflags_0_8;
      5'b01001:
        casez_tmp_29 = rob_fflags_0_9;
      5'b01010:
        casez_tmp_29 = rob_fflags_0_10;
      5'b01011:
        casez_tmp_29 = rob_fflags_0_11;
      5'b01100:
        casez_tmp_29 = rob_fflags_0_12;
      5'b01101:
        casez_tmp_29 = rob_fflags_0_13;
      5'b01110:
        casez_tmp_29 = rob_fflags_0_14;
      5'b01111:
        casez_tmp_29 = rob_fflags_0_15;
      5'b10000:
        casez_tmp_29 = rob_fflags_0_16;
      5'b10001:
        casez_tmp_29 = rob_fflags_0_17;
      5'b10010:
        casez_tmp_29 = rob_fflags_0_18;
      5'b10011:
        casez_tmp_29 = rob_fflags_0_19;
      5'b10100:
        casez_tmp_29 = rob_fflags_0_20;
      5'b10101:
        casez_tmp_29 = rob_fflags_0_21;
      5'b10110:
        casez_tmp_29 = rob_fflags_0_22;
      5'b10111:
        casez_tmp_29 = rob_fflags_0_23;
      5'b11000:
        casez_tmp_29 = rob_fflags_0_24;
      5'b11001:
        casez_tmp_29 = rob_fflags_0_25;
      5'b11010:
        casez_tmp_29 = rob_fflags_0_26;
      5'b11011:
        casez_tmp_29 = rob_fflags_0_27;
      5'b11100:
        casez_tmp_29 = rob_fflags_0_28;
      5'b11101:
        casez_tmp_29 = rob_fflags_0_29;
      5'b11110:
        casez_tmp_29 = rob_fflags_0_30;
      default:
        casez_tmp_29 = rob_fflags_0_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_30 = rob_uop__0_uses_ldq;
      5'b00001:
        casez_tmp_30 = rob_uop__1_uses_ldq;
      5'b00010:
        casez_tmp_30 = rob_uop__2_uses_ldq;
      5'b00011:
        casez_tmp_30 = rob_uop__3_uses_ldq;
      5'b00100:
        casez_tmp_30 = rob_uop__4_uses_ldq;
      5'b00101:
        casez_tmp_30 = rob_uop__5_uses_ldq;
      5'b00110:
        casez_tmp_30 = rob_uop__6_uses_ldq;
      5'b00111:
        casez_tmp_30 = rob_uop__7_uses_ldq;
      5'b01000:
        casez_tmp_30 = rob_uop__8_uses_ldq;
      5'b01001:
        casez_tmp_30 = rob_uop__9_uses_ldq;
      5'b01010:
        casez_tmp_30 = rob_uop__10_uses_ldq;
      5'b01011:
        casez_tmp_30 = rob_uop__11_uses_ldq;
      5'b01100:
        casez_tmp_30 = rob_uop__12_uses_ldq;
      5'b01101:
        casez_tmp_30 = rob_uop__13_uses_ldq;
      5'b01110:
        casez_tmp_30 = rob_uop__14_uses_ldq;
      5'b01111:
        casez_tmp_30 = rob_uop__15_uses_ldq;
      5'b10000:
        casez_tmp_30 = rob_uop__16_uses_ldq;
      5'b10001:
        casez_tmp_30 = rob_uop__17_uses_ldq;
      5'b10010:
        casez_tmp_30 = rob_uop__18_uses_ldq;
      5'b10011:
        casez_tmp_30 = rob_uop__19_uses_ldq;
      5'b10100:
        casez_tmp_30 = rob_uop__20_uses_ldq;
      5'b10101:
        casez_tmp_30 = rob_uop__21_uses_ldq;
      5'b10110:
        casez_tmp_30 = rob_uop__22_uses_ldq;
      5'b10111:
        casez_tmp_30 = rob_uop__23_uses_ldq;
      5'b11000:
        casez_tmp_30 = rob_uop__24_uses_ldq;
      5'b11001:
        casez_tmp_30 = rob_uop__25_uses_ldq;
      5'b11010:
        casez_tmp_30 = rob_uop__26_uses_ldq;
      5'b11011:
        casez_tmp_30 = rob_uop__27_uses_ldq;
      5'b11100:
        casez_tmp_30 = rob_uop__28_uses_ldq;
      5'b11101:
        casez_tmp_30 = rob_uop__29_uses_ldq;
      5'b11110:
        casez_tmp_30 = rob_uop__30_uses_ldq;
      default:
        casez_tmp_30 = rob_uop__31_uses_ldq;
    endcase
  end // always @(*)
  reg  [6:0]  rob_uop_1_0_uopc;
  reg         rob_uop_1_0_is_rvc;
  reg  [19:0] rob_uop_1_0_br_mask;
  reg  [5:0]  rob_uop_1_0_ftq_idx;
  reg         rob_uop_1_0_edge_inst;
  reg  [5:0]  rob_uop_1_0_pc_lob;
  reg  [6:0]  rob_uop_1_0_pdst;
  reg  [6:0]  rob_uop_1_0_stale_pdst;
  reg         rob_uop_1_0_is_fencei;
  reg         rob_uop_1_0_uses_ldq;
  reg         rob_uop_1_0_uses_stq;
  reg         rob_uop_1_0_is_sys_pc2epc;
  reg         rob_uop_1_0_flush_on_commit;
  reg  [5:0]  rob_uop_1_0_ldst;
  reg         rob_uop_1_0_ldst_val;
  reg  [1:0]  rob_uop_1_0_dst_rtype;
  reg         rob_uop_1_0_fp_val;
  reg  [6:0]  rob_uop_1_1_uopc;
  reg         rob_uop_1_1_is_rvc;
  reg  [19:0] rob_uop_1_1_br_mask;
  reg  [5:0]  rob_uop_1_1_ftq_idx;
  reg         rob_uop_1_1_edge_inst;
  reg  [5:0]  rob_uop_1_1_pc_lob;
  reg  [6:0]  rob_uop_1_1_pdst;
  reg  [6:0]  rob_uop_1_1_stale_pdst;
  reg         rob_uop_1_1_is_fencei;
  reg         rob_uop_1_1_uses_ldq;
  reg         rob_uop_1_1_uses_stq;
  reg         rob_uop_1_1_is_sys_pc2epc;
  reg         rob_uop_1_1_flush_on_commit;
  reg  [5:0]  rob_uop_1_1_ldst;
  reg         rob_uop_1_1_ldst_val;
  reg  [1:0]  rob_uop_1_1_dst_rtype;
  reg         rob_uop_1_1_fp_val;
  reg  [6:0]  rob_uop_1_2_uopc;
  reg         rob_uop_1_2_is_rvc;
  reg  [19:0] rob_uop_1_2_br_mask;
  reg  [5:0]  rob_uop_1_2_ftq_idx;
  reg         rob_uop_1_2_edge_inst;
  reg  [5:0]  rob_uop_1_2_pc_lob;
  reg  [6:0]  rob_uop_1_2_pdst;
  reg  [6:0]  rob_uop_1_2_stale_pdst;
  reg         rob_uop_1_2_is_fencei;
  reg         rob_uop_1_2_uses_ldq;
  reg         rob_uop_1_2_uses_stq;
  reg         rob_uop_1_2_is_sys_pc2epc;
  reg         rob_uop_1_2_flush_on_commit;
  reg  [5:0]  rob_uop_1_2_ldst;
  reg         rob_uop_1_2_ldst_val;
  reg  [1:0]  rob_uop_1_2_dst_rtype;
  reg         rob_uop_1_2_fp_val;
  reg  [6:0]  rob_uop_1_3_uopc;
  reg         rob_uop_1_3_is_rvc;
  reg  [19:0] rob_uop_1_3_br_mask;
  reg  [5:0]  rob_uop_1_3_ftq_idx;
  reg         rob_uop_1_3_edge_inst;
  reg  [5:0]  rob_uop_1_3_pc_lob;
  reg  [6:0]  rob_uop_1_3_pdst;
  reg  [6:0]  rob_uop_1_3_stale_pdst;
  reg         rob_uop_1_3_is_fencei;
  reg         rob_uop_1_3_uses_ldq;
  reg         rob_uop_1_3_uses_stq;
  reg         rob_uop_1_3_is_sys_pc2epc;
  reg         rob_uop_1_3_flush_on_commit;
  reg  [5:0]  rob_uop_1_3_ldst;
  reg         rob_uop_1_3_ldst_val;
  reg  [1:0]  rob_uop_1_3_dst_rtype;
  reg         rob_uop_1_3_fp_val;
  reg  [6:0]  rob_uop_1_4_uopc;
  reg         rob_uop_1_4_is_rvc;
  reg  [19:0] rob_uop_1_4_br_mask;
  reg  [5:0]  rob_uop_1_4_ftq_idx;
  reg         rob_uop_1_4_edge_inst;
  reg  [5:0]  rob_uop_1_4_pc_lob;
  reg  [6:0]  rob_uop_1_4_pdst;
  reg  [6:0]  rob_uop_1_4_stale_pdst;
  reg         rob_uop_1_4_is_fencei;
  reg         rob_uop_1_4_uses_ldq;
  reg         rob_uop_1_4_uses_stq;
  reg         rob_uop_1_4_is_sys_pc2epc;
  reg         rob_uop_1_4_flush_on_commit;
  reg  [5:0]  rob_uop_1_4_ldst;
  reg         rob_uop_1_4_ldst_val;
  reg  [1:0]  rob_uop_1_4_dst_rtype;
  reg         rob_uop_1_4_fp_val;
  reg  [6:0]  rob_uop_1_5_uopc;
  reg         rob_uop_1_5_is_rvc;
  reg  [19:0] rob_uop_1_5_br_mask;
  reg  [5:0]  rob_uop_1_5_ftq_idx;
  reg         rob_uop_1_5_edge_inst;
  reg  [5:0]  rob_uop_1_5_pc_lob;
  reg  [6:0]  rob_uop_1_5_pdst;
  reg  [6:0]  rob_uop_1_5_stale_pdst;
  reg         rob_uop_1_5_is_fencei;
  reg         rob_uop_1_5_uses_ldq;
  reg         rob_uop_1_5_uses_stq;
  reg         rob_uop_1_5_is_sys_pc2epc;
  reg         rob_uop_1_5_flush_on_commit;
  reg  [5:0]  rob_uop_1_5_ldst;
  reg         rob_uop_1_5_ldst_val;
  reg  [1:0]  rob_uop_1_5_dst_rtype;
  reg         rob_uop_1_5_fp_val;
  reg  [6:0]  rob_uop_1_6_uopc;
  reg         rob_uop_1_6_is_rvc;
  reg  [19:0] rob_uop_1_6_br_mask;
  reg  [5:0]  rob_uop_1_6_ftq_idx;
  reg         rob_uop_1_6_edge_inst;
  reg  [5:0]  rob_uop_1_6_pc_lob;
  reg  [6:0]  rob_uop_1_6_pdst;
  reg  [6:0]  rob_uop_1_6_stale_pdst;
  reg         rob_uop_1_6_is_fencei;
  reg         rob_uop_1_6_uses_ldq;
  reg         rob_uop_1_6_uses_stq;
  reg         rob_uop_1_6_is_sys_pc2epc;
  reg         rob_uop_1_6_flush_on_commit;
  reg  [5:0]  rob_uop_1_6_ldst;
  reg         rob_uop_1_6_ldst_val;
  reg  [1:0]  rob_uop_1_6_dst_rtype;
  reg         rob_uop_1_6_fp_val;
  reg  [6:0]  rob_uop_1_7_uopc;
  reg         rob_uop_1_7_is_rvc;
  reg  [19:0] rob_uop_1_7_br_mask;
  reg  [5:0]  rob_uop_1_7_ftq_idx;
  reg         rob_uop_1_7_edge_inst;
  reg  [5:0]  rob_uop_1_7_pc_lob;
  reg  [6:0]  rob_uop_1_7_pdst;
  reg  [6:0]  rob_uop_1_7_stale_pdst;
  reg         rob_uop_1_7_is_fencei;
  reg         rob_uop_1_7_uses_ldq;
  reg         rob_uop_1_7_uses_stq;
  reg         rob_uop_1_7_is_sys_pc2epc;
  reg         rob_uop_1_7_flush_on_commit;
  reg  [5:0]  rob_uop_1_7_ldst;
  reg         rob_uop_1_7_ldst_val;
  reg  [1:0]  rob_uop_1_7_dst_rtype;
  reg         rob_uop_1_7_fp_val;
  reg  [6:0]  rob_uop_1_8_uopc;
  reg         rob_uop_1_8_is_rvc;
  reg  [19:0] rob_uop_1_8_br_mask;
  reg  [5:0]  rob_uop_1_8_ftq_idx;
  reg         rob_uop_1_8_edge_inst;
  reg  [5:0]  rob_uop_1_8_pc_lob;
  reg  [6:0]  rob_uop_1_8_pdst;
  reg  [6:0]  rob_uop_1_8_stale_pdst;
  reg         rob_uop_1_8_is_fencei;
  reg         rob_uop_1_8_uses_ldq;
  reg         rob_uop_1_8_uses_stq;
  reg         rob_uop_1_8_is_sys_pc2epc;
  reg         rob_uop_1_8_flush_on_commit;
  reg  [5:0]  rob_uop_1_8_ldst;
  reg         rob_uop_1_8_ldst_val;
  reg  [1:0]  rob_uop_1_8_dst_rtype;
  reg         rob_uop_1_8_fp_val;
  reg  [6:0]  rob_uop_1_9_uopc;
  reg         rob_uop_1_9_is_rvc;
  reg  [19:0] rob_uop_1_9_br_mask;
  reg  [5:0]  rob_uop_1_9_ftq_idx;
  reg         rob_uop_1_9_edge_inst;
  reg  [5:0]  rob_uop_1_9_pc_lob;
  reg  [6:0]  rob_uop_1_9_pdst;
  reg  [6:0]  rob_uop_1_9_stale_pdst;
  reg         rob_uop_1_9_is_fencei;
  reg         rob_uop_1_9_uses_ldq;
  reg         rob_uop_1_9_uses_stq;
  reg         rob_uop_1_9_is_sys_pc2epc;
  reg         rob_uop_1_9_flush_on_commit;
  reg  [5:0]  rob_uop_1_9_ldst;
  reg         rob_uop_1_9_ldst_val;
  reg  [1:0]  rob_uop_1_9_dst_rtype;
  reg         rob_uop_1_9_fp_val;
  reg  [6:0]  rob_uop_1_10_uopc;
  reg         rob_uop_1_10_is_rvc;
  reg  [19:0] rob_uop_1_10_br_mask;
  reg  [5:0]  rob_uop_1_10_ftq_idx;
  reg         rob_uop_1_10_edge_inst;
  reg  [5:0]  rob_uop_1_10_pc_lob;
  reg  [6:0]  rob_uop_1_10_pdst;
  reg  [6:0]  rob_uop_1_10_stale_pdst;
  reg         rob_uop_1_10_is_fencei;
  reg         rob_uop_1_10_uses_ldq;
  reg         rob_uop_1_10_uses_stq;
  reg         rob_uop_1_10_is_sys_pc2epc;
  reg         rob_uop_1_10_flush_on_commit;
  reg  [5:0]  rob_uop_1_10_ldst;
  reg         rob_uop_1_10_ldst_val;
  reg  [1:0]  rob_uop_1_10_dst_rtype;
  reg         rob_uop_1_10_fp_val;
  reg  [6:0]  rob_uop_1_11_uopc;
  reg         rob_uop_1_11_is_rvc;
  reg  [19:0] rob_uop_1_11_br_mask;
  reg  [5:0]  rob_uop_1_11_ftq_idx;
  reg         rob_uop_1_11_edge_inst;
  reg  [5:0]  rob_uop_1_11_pc_lob;
  reg  [6:0]  rob_uop_1_11_pdst;
  reg  [6:0]  rob_uop_1_11_stale_pdst;
  reg         rob_uop_1_11_is_fencei;
  reg         rob_uop_1_11_uses_ldq;
  reg         rob_uop_1_11_uses_stq;
  reg         rob_uop_1_11_is_sys_pc2epc;
  reg         rob_uop_1_11_flush_on_commit;
  reg  [5:0]  rob_uop_1_11_ldst;
  reg         rob_uop_1_11_ldst_val;
  reg  [1:0]  rob_uop_1_11_dst_rtype;
  reg         rob_uop_1_11_fp_val;
  reg  [6:0]  rob_uop_1_12_uopc;
  reg         rob_uop_1_12_is_rvc;
  reg  [19:0] rob_uop_1_12_br_mask;
  reg  [5:0]  rob_uop_1_12_ftq_idx;
  reg         rob_uop_1_12_edge_inst;
  reg  [5:0]  rob_uop_1_12_pc_lob;
  reg  [6:0]  rob_uop_1_12_pdst;
  reg  [6:0]  rob_uop_1_12_stale_pdst;
  reg         rob_uop_1_12_is_fencei;
  reg         rob_uop_1_12_uses_ldq;
  reg         rob_uop_1_12_uses_stq;
  reg         rob_uop_1_12_is_sys_pc2epc;
  reg         rob_uop_1_12_flush_on_commit;
  reg  [5:0]  rob_uop_1_12_ldst;
  reg         rob_uop_1_12_ldst_val;
  reg  [1:0]  rob_uop_1_12_dst_rtype;
  reg         rob_uop_1_12_fp_val;
  reg  [6:0]  rob_uop_1_13_uopc;
  reg         rob_uop_1_13_is_rvc;
  reg  [19:0] rob_uop_1_13_br_mask;
  reg  [5:0]  rob_uop_1_13_ftq_idx;
  reg         rob_uop_1_13_edge_inst;
  reg  [5:0]  rob_uop_1_13_pc_lob;
  reg  [6:0]  rob_uop_1_13_pdst;
  reg  [6:0]  rob_uop_1_13_stale_pdst;
  reg         rob_uop_1_13_is_fencei;
  reg         rob_uop_1_13_uses_ldq;
  reg         rob_uop_1_13_uses_stq;
  reg         rob_uop_1_13_is_sys_pc2epc;
  reg         rob_uop_1_13_flush_on_commit;
  reg  [5:0]  rob_uop_1_13_ldst;
  reg         rob_uop_1_13_ldst_val;
  reg  [1:0]  rob_uop_1_13_dst_rtype;
  reg         rob_uop_1_13_fp_val;
  reg  [6:0]  rob_uop_1_14_uopc;
  reg         rob_uop_1_14_is_rvc;
  reg  [19:0] rob_uop_1_14_br_mask;
  reg  [5:0]  rob_uop_1_14_ftq_idx;
  reg         rob_uop_1_14_edge_inst;
  reg  [5:0]  rob_uop_1_14_pc_lob;
  reg  [6:0]  rob_uop_1_14_pdst;
  reg  [6:0]  rob_uop_1_14_stale_pdst;
  reg         rob_uop_1_14_is_fencei;
  reg         rob_uop_1_14_uses_ldq;
  reg         rob_uop_1_14_uses_stq;
  reg         rob_uop_1_14_is_sys_pc2epc;
  reg         rob_uop_1_14_flush_on_commit;
  reg  [5:0]  rob_uop_1_14_ldst;
  reg         rob_uop_1_14_ldst_val;
  reg  [1:0]  rob_uop_1_14_dst_rtype;
  reg         rob_uop_1_14_fp_val;
  reg  [6:0]  rob_uop_1_15_uopc;
  reg         rob_uop_1_15_is_rvc;
  reg  [19:0] rob_uop_1_15_br_mask;
  reg  [5:0]  rob_uop_1_15_ftq_idx;
  reg         rob_uop_1_15_edge_inst;
  reg  [5:0]  rob_uop_1_15_pc_lob;
  reg  [6:0]  rob_uop_1_15_pdst;
  reg  [6:0]  rob_uop_1_15_stale_pdst;
  reg         rob_uop_1_15_is_fencei;
  reg         rob_uop_1_15_uses_ldq;
  reg         rob_uop_1_15_uses_stq;
  reg         rob_uop_1_15_is_sys_pc2epc;
  reg         rob_uop_1_15_flush_on_commit;
  reg  [5:0]  rob_uop_1_15_ldst;
  reg         rob_uop_1_15_ldst_val;
  reg  [1:0]  rob_uop_1_15_dst_rtype;
  reg         rob_uop_1_15_fp_val;
  reg  [6:0]  rob_uop_1_16_uopc;
  reg         rob_uop_1_16_is_rvc;
  reg  [19:0] rob_uop_1_16_br_mask;
  reg  [5:0]  rob_uop_1_16_ftq_idx;
  reg         rob_uop_1_16_edge_inst;
  reg  [5:0]  rob_uop_1_16_pc_lob;
  reg  [6:0]  rob_uop_1_16_pdst;
  reg  [6:0]  rob_uop_1_16_stale_pdst;
  reg         rob_uop_1_16_is_fencei;
  reg         rob_uop_1_16_uses_ldq;
  reg         rob_uop_1_16_uses_stq;
  reg         rob_uop_1_16_is_sys_pc2epc;
  reg         rob_uop_1_16_flush_on_commit;
  reg  [5:0]  rob_uop_1_16_ldst;
  reg         rob_uop_1_16_ldst_val;
  reg  [1:0]  rob_uop_1_16_dst_rtype;
  reg         rob_uop_1_16_fp_val;
  reg  [6:0]  rob_uop_1_17_uopc;
  reg         rob_uop_1_17_is_rvc;
  reg  [19:0] rob_uop_1_17_br_mask;
  reg  [5:0]  rob_uop_1_17_ftq_idx;
  reg         rob_uop_1_17_edge_inst;
  reg  [5:0]  rob_uop_1_17_pc_lob;
  reg  [6:0]  rob_uop_1_17_pdst;
  reg  [6:0]  rob_uop_1_17_stale_pdst;
  reg         rob_uop_1_17_is_fencei;
  reg         rob_uop_1_17_uses_ldq;
  reg         rob_uop_1_17_uses_stq;
  reg         rob_uop_1_17_is_sys_pc2epc;
  reg         rob_uop_1_17_flush_on_commit;
  reg  [5:0]  rob_uop_1_17_ldst;
  reg         rob_uop_1_17_ldst_val;
  reg  [1:0]  rob_uop_1_17_dst_rtype;
  reg         rob_uop_1_17_fp_val;
  reg  [6:0]  rob_uop_1_18_uopc;
  reg         rob_uop_1_18_is_rvc;
  reg  [19:0] rob_uop_1_18_br_mask;
  reg  [5:0]  rob_uop_1_18_ftq_idx;
  reg         rob_uop_1_18_edge_inst;
  reg  [5:0]  rob_uop_1_18_pc_lob;
  reg  [6:0]  rob_uop_1_18_pdst;
  reg  [6:0]  rob_uop_1_18_stale_pdst;
  reg         rob_uop_1_18_is_fencei;
  reg         rob_uop_1_18_uses_ldq;
  reg         rob_uop_1_18_uses_stq;
  reg         rob_uop_1_18_is_sys_pc2epc;
  reg         rob_uop_1_18_flush_on_commit;
  reg  [5:0]  rob_uop_1_18_ldst;
  reg         rob_uop_1_18_ldst_val;
  reg  [1:0]  rob_uop_1_18_dst_rtype;
  reg         rob_uop_1_18_fp_val;
  reg  [6:0]  rob_uop_1_19_uopc;
  reg         rob_uop_1_19_is_rvc;
  reg  [19:0] rob_uop_1_19_br_mask;
  reg  [5:0]  rob_uop_1_19_ftq_idx;
  reg         rob_uop_1_19_edge_inst;
  reg  [5:0]  rob_uop_1_19_pc_lob;
  reg  [6:0]  rob_uop_1_19_pdst;
  reg  [6:0]  rob_uop_1_19_stale_pdst;
  reg         rob_uop_1_19_is_fencei;
  reg         rob_uop_1_19_uses_ldq;
  reg         rob_uop_1_19_uses_stq;
  reg         rob_uop_1_19_is_sys_pc2epc;
  reg         rob_uop_1_19_flush_on_commit;
  reg  [5:0]  rob_uop_1_19_ldst;
  reg         rob_uop_1_19_ldst_val;
  reg  [1:0]  rob_uop_1_19_dst_rtype;
  reg         rob_uop_1_19_fp_val;
  reg  [6:0]  rob_uop_1_20_uopc;
  reg         rob_uop_1_20_is_rvc;
  reg  [19:0] rob_uop_1_20_br_mask;
  reg  [5:0]  rob_uop_1_20_ftq_idx;
  reg         rob_uop_1_20_edge_inst;
  reg  [5:0]  rob_uop_1_20_pc_lob;
  reg  [6:0]  rob_uop_1_20_pdst;
  reg  [6:0]  rob_uop_1_20_stale_pdst;
  reg         rob_uop_1_20_is_fencei;
  reg         rob_uop_1_20_uses_ldq;
  reg         rob_uop_1_20_uses_stq;
  reg         rob_uop_1_20_is_sys_pc2epc;
  reg         rob_uop_1_20_flush_on_commit;
  reg  [5:0]  rob_uop_1_20_ldst;
  reg         rob_uop_1_20_ldst_val;
  reg  [1:0]  rob_uop_1_20_dst_rtype;
  reg         rob_uop_1_20_fp_val;
  reg  [6:0]  rob_uop_1_21_uopc;
  reg         rob_uop_1_21_is_rvc;
  reg  [19:0] rob_uop_1_21_br_mask;
  reg  [5:0]  rob_uop_1_21_ftq_idx;
  reg         rob_uop_1_21_edge_inst;
  reg  [5:0]  rob_uop_1_21_pc_lob;
  reg  [6:0]  rob_uop_1_21_pdst;
  reg  [6:0]  rob_uop_1_21_stale_pdst;
  reg         rob_uop_1_21_is_fencei;
  reg         rob_uop_1_21_uses_ldq;
  reg         rob_uop_1_21_uses_stq;
  reg         rob_uop_1_21_is_sys_pc2epc;
  reg         rob_uop_1_21_flush_on_commit;
  reg  [5:0]  rob_uop_1_21_ldst;
  reg         rob_uop_1_21_ldst_val;
  reg  [1:0]  rob_uop_1_21_dst_rtype;
  reg         rob_uop_1_21_fp_val;
  reg  [6:0]  rob_uop_1_22_uopc;
  reg         rob_uop_1_22_is_rvc;
  reg  [19:0] rob_uop_1_22_br_mask;
  reg  [5:0]  rob_uop_1_22_ftq_idx;
  reg         rob_uop_1_22_edge_inst;
  reg  [5:0]  rob_uop_1_22_pc_lob;
  reg  [6:0]  rob_uop_1_22_pdst;
  reg  [6:0]  rob_uop_1_22_stale_pdst;
  reg         rob_uop_1_22_is_fencei;
  reg         rob_uop_1_22_uses_ldq;
  reg         rob_uop_1_22_uses_stq;
  reg         rob_uop_1_22_is_sys_pc2epc;
  reg         rob_uop_1_22_flush_on_commit;
  reg  [5:0]  rob_uop_1_22_ldst;
  reg         rob_uop_1_22_ldst_val;
  reg  [1:0]  rob_uop_1_22_dst_rtype;
  reg         rob_uop_1_22_fp_val;
  reg  [6:0]  rob_uop_1_23_uopc;
  reg         rob_uop_1_23_is_rvc;
  reg  [19:0] rob_uop_1_23_br_mask;
  reg  [5:0]  rob_uop_1_23_ftq_idx;
  reg         rob_uop_1_23_edge_inst;
  reg  [5:0]  rob_uop_1_23_pc_lob;
  reg  [6:0]  rob_uop_1_23_pdst;
  reg  [6:0]  rob_uop_1_23_stale_pdst;
  reg         rob_uop_1_23_is_fencei;
  reg         rob_uop_1_23_uses_ldq;
  reg         rob_uop_1_23_uses_stq;
  reg         rob_uop_1_23_is_sys_pc2epc;
  reg         rob_uop_1_23_flush_on_commit;
  reg  [5:0]  rob_uop_1_23_ldst;
  reg         rob_uop_1_23_ldst_val;
  reg  [1:0]  rob_uop_1_23_dst_rtype;
  reg         rob_uop_1_23_fp_val;
  reg  [6:0]  rob_uop_1_24_uopc;
  reg         rob_uop_1_24_is_rvc;
  reg  [19:0] rob_uop_1_24_br_mask;
  reg  [5:0]  rob_uop_1_24_ftq_idx;
  reg         rob_uop_1_24_edge_inst;
  reg  [5:0]  rob_uop_1_24_pc_lob;
  reg  [6:0]  rob_uop_1_24_pdst;
  reg  [6:0]  rob_uop_1_24_stale_pdst;
  reg         rob_uop_1_24_is_fencei;
  reg         rob_uop_1_24_uses_ldq;
  reg         rob_uop_1_24_uses_stq;
  reg         rob_uop_1_24_is_sys_pc2epc;
  reg         rob_uop_1_24_flush_on_commit;
  reg  [5:0]  rob_uop_1_24_ldst;
  reg         rob_uop_1_24_ldst_val;
  reg  [1:0]  rob_uop_1_24_dst_rtype;
  reg         rob_uop_1_24_fp_val;
  reg  [6:0]  rob_uop_1_25_uopc;
  reg         rob_uop_1_25_is_rvc;
  reg  [19:0] rob_uop_1_25_br_mask;
  reg  [5:0]  rob_uop_1_25_ftq_idx;
  reg         rob_uop_1_25_edge_inst;
  reg  [5:0]  rob_uop_1_25_pc_lob;
  reg  [6:0]  rob_uop_1_25_pdst;
  reg  [6:0]  rob_uop_1_25_stale_pdst;
  reg         rob_uop_1_25_is_fencei;
  reg         rob_uop_1_25_uses_ldq;
  reg         rob_uop_1_25_uses_stq;
  reg         rob_uop_1_25_is_sys_pc2epc;
  reg         rob_uop_1_25_flush_on_commit;
  reg  [5:0]  rob_uop_1_25_ldst;
  reg         rob_uop_1_25_ldst_val;
  reg  [1:0]  rob_uop_1_25_dst_rtype;
  reg         rob_uop_1_25_fp_val;
  reg  [6:0]  rob_uop_1_26_uopc;
  reg         rob_uop_1_26_is_rvc;
  reg  [19:0] rob_uop_1_26_br_mask;
  reg  [5:0]  rob_uop_1_26_ftq_idx;
  reg         rob_uop_1_26_edge_inst;
  reg  [5:0]  rob_uop_1_26_pc_lob;
  reg  [6:0]  rob_uop_1_26_pdst;
  reg  [6:0]  rob_uop_1_26_stale_pdst;
  reg         rob_uop_1_26_is_fencei;
  reg         rob_uop_1_26_uses_ldq;
  reg         rob_uop_1_26_uses_stq;
  reg         rob_uop_1_26_is_sys_pc2epc;
  reg         rob_uop_1_26_flush_on_commit;
  reg  [5:0]  rob_uop_1_26_ldst;
  reg         rob_uop_1_26_ldst_val;
  reg  [1:0]  rob_uop_1_26_dst_rtype;
  reg         rob_uop_1_26_fp_val;
  reg  [6:0]  rob_uop_1_27_uopc;
  reg         rob_uop_1_27_is_rvc;
  reg  [19:0] rob_uop_1_27_br_mask;
  reg  [5:0]  rob_uop_1_27_ftq_idx;
  reg         rob_uop_1_27_edge_inst;
  reg  [5:0]  rob_uop_1_27_pc_lob;
  reg  [6:0]  rob_uop_1_27_pdst;
  reg  [6:0]  rob_uop_1_27_stale_pdst;
  reg         rob_uop_1_27_is_fencei;
  reg         rob_uop_1_27_uses_ldq;
  reg         rob_uop_1_27_uses_stq;
  reg         rob_uop_1_27_is_sys_pc2epc;
  reg         rob_uop_1_27_flush_on_commit;
  reg  [5:0]  rob_uop_1_27_ldst;
  reg         rob_uop_1_27_ldst_val;
  reg  [1:0]  rob_uop_1_27_dst_rtype;
  reg         rob_uop_1_27_fp_val;
  reg  [6:0]  rob_uop_1_28_uopc;
  reg         rob_uop_1_28_is_rvc;
  reg  [19:0] rob_uop_1_28_br_mask;
  reg  [5:0]  rob_uop_1_28_ftq_idx;
  reg         rob_uop_1_28_edge_inst;
  reg  [5:0]  rob_uop_1_28_pc_lob;
  reg  [6:0]  rob_uop_1_28_pdst;
  reg  [6:0]  rob_uop_1_28_stale_pdst;
  reg         rob_uop_1_28_is_fencei;
  reg         rob_uop_1_28_uses_ldq;
  reg         rob_uop_1_28_uses_stq;
  reg         rob_uop_1_28_is_sys_pc2epc;
  reg         rob_uop_1_28_flush_on_commit;
  reg  [5:0]  rob_uop_1_28_ldst;
  reg         rob_uop_1_28_ldst_val;
  reg  [1:0]  rob_uop_1_28_dst_rtype;
  reg         rob_uop_1_28_fp_val;
  reg  [6:0]  rob_uop_1_29_uopc;
  reg         rob_uop_1_29_is_rvc;
  reg  [19:0] rob_uop_1_29_br_mask;
  reg  [5:0]  rob_uop_1_29_ftq_idx;
  reg         rob_uop_1_29_edge_inst;
  reg  [5:0]  rob_uop_1_29_pc_lob;
  reg  [6:0]  rob_uop_1_29_pdst;
  reg  [6:0]  rob_uop_1_29_stale_pdst;
  reg         rob_uop_1_29_is_fencei;
  reg         rob_uop_1_29_uses_ldq;
  reg         rob_uop_1_29_uses_stq;
  reg         rob_uop_1_29_is_sys_pc2epc;
  reg         rob_uop_1_29_flush_on_commit;
  reg  [5:0]  rob_uop_1_29_ldst;
  reg         rob_uop_1_29_ldst_val;
  reg  [1:0]  rob_uop_1_29_dst_rtype;
  reg         rob_uop_1_29_fp_val;
  reg  [6:0]  rob_uop_1_30_uopc;
  reg         rob_uop_1_30_is_rvc;
  reg  [19:0] rob_uop_1_30_br_mask;
  reg  [5:0]  rob_uop_1_30_ftq_idx;
  reg         rob_uop_1_30_edge_inst;
  reg  [5:0]  rob_uop_1_30_pc_lob;
  reg  [6:0]  rob_uop_1_30_pdst;
  reg  [6:0]  rob_uop_1_30_stale_pdst;
  reg         rob_uop_1_30_is_fencei;
  reg         rob_uop_1_30_uses_ldq;
  reg         rob_uop_1_30_uses_stq;
  reg         rob_uop_1_30_is_sys_pc2epc;
  reg         rob_uop_1_30_flush_on_commit;
  reg  [5:0]  rob_uop_1_30_ldst;
  reg         rob_uop_1_30_ldst_val;
  reg  [1:0]  rob_uop_1_30_dst_rtype;
  reg         rob_uop_1_30_fp_val;
  reg  [6:0]  rob_uop_1_31_uopc;
  reg         rob_uop_1_31_is_rvc;
  reg  [19:0] rob_uop_1_31_br_mask;
  reg  [5:0]  rob_uop_1_31_ftq_idx;
  reg         rob_uop_1_31_edge_inst;
  reg  [5:0]  rob_uop_1_31_pc_lob;
  reg  [6:0]  rob_uop_1_31_pdst;
  reg  [6:0]  rob_uop_1_31_stale_pdst;
  reg         rob_uop_1_31_is_fencei;
  reg         rob_uop_1_31_uses_ldq;
  reg         rob_uop_1_31_uses_stq;
  reg         rob_uop_1_31_is_sys_pc2epc;
  reg         rob_uop_1_31_flush_on_commit;
  reg  [5:0]  rob_uop_1_31_ldst;
  reg         rob_uop_1_31_ldst_val;
  reg  [1:0]  rob_uop_1_31_dst_rtype;
  reg         rob_uop_1_31_fp_val;
  reg         rob_predicated_1_0;
  reg         rob_predicated_1_1;
  reg         rob_predicated_1_2;
  reg         rob_predicated_1_3;
  reg         rob_predicated_1_4;
  reg         rob_predicated_1_5;
  reg         rob_predicated_1_6;
  reg         rob_predicated_1_7;
  reg         rob_predicated_1_8;
  reg         rob_predicated_1_9;
  reg         rob_predicated_1_10;
  reg         rob_predicated_1_11;
  reg         rob_predicated_1_12;
  reg         rob_predicated_1_13;
  reg         rob_predicated_1_14;
  reg         rob_predicated_1_15;
  reg         rob_predicated_1_16;
  reg         rob_predicated_1_17;
  reg         rob_predicated_1_18;
  reg         rob_predicated_1_19;
  reg         rob_predicated_1_20;
  reg         rob_predicated_1_21;
  reg         rob_predicated_1_22;
  reg         rob_predicated_1_23;
  reg         rob_predicated_1_24;
  reg         rob_predicated_1_25;
  reg         rob_predicated_1_26;
  reg         rob_predicated_1_27;
  reg         rob_predicated_1_28;
  reg         rob_predicated_1_29;
  reg         rob_predicated_1_30;
  reg         rob_predicated_1_31;
  wire        _GEN_898 = io_enq_valids_1 & _GEN_2;
  wire        _GEN_899 = io_enq_valids_1 & _GEN_3;
  wire        _GEN_900 = io_enq_valids_1 & _GEN_4;
  wire        _GEN_901 = io_enq_valids_1 & _GEN_5;
  wire        _GEN_902 = io_enq_valids_1 & _GEN_6;
  wire        _GEN_903 = io_enq_valids_1 & _GEN_7;
  wire        _GEN_904 = io_enq_valids_1 & _GEN_8;
  wire        _GEN_905 = io_enq_valids_1 & _GEN_9;
  wire        _GEN_906 = io_enq_valids_1 & _GEN_10;
  wire        _GEN_907 = io_enq_valids_1 & _GEN_11;
  wire        _GEN_908 = io_enq_valids_1 & _GEN_12;
  wire        _GEN_909 = io_enq_valids_1 & _GEN_13;
  wire        _GEN_910 = io_enq_valids_1 & _GEN_14;
  wire        _GEN_911 = io_enq_valids_1 & _GEN_15;
  wire        _GEN_912 = io_enq_valids_1 & _GEN_16;
  wire        _GEN_913 = io_enq_valids_1 & _GEN_17;
  wire        _GEN_914 = io_enq_valids_1 & _GEN_18;
  wire        _GEN_915 = io_enq_valids_1 & _GEN_19;
  wire        _GEN_916 = io_enq_valids_1 & _GEN_20;
  wire        _GEN_917 = io_enq_valids_1 & _GEN_21;
  wire        _GEN_918 = io_enq_valids_1 & _GEN_22;
  wire        _GEN_919 = io_enq_valids_1 & _GEN_23;
  wire        _GEN_920 = io_enq_valids_1 & _GEN_24;
  wire        _GEN_921 = io_enq_valids_1 & _GEN_25;
  wire        _GEN_922 = io_enq_valids_1 & _GEN_26;
  wire        _GEN_923 = io_enq_valids_1 & _GEN_27;
  wire        _GEN_924 = io_enq_valids_1 & _GEN_28;
  wire        _GEN_925 = io_enq_valids_1 & _GEN_29;
  wire        _GEN_926 = io_enq_valids_1 & _GEN_30;
  wire        _GEN_927 = io_enq_valids_1 & _GEN_31;
  wire        _GEN_928 = io_enq_valids_1 & _GEN_32;
  wire        _GEN_929 = io_enq_valids_1 & (&rob_tail);
  wire        _GEN_930 = io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_931 = _GEN_930 & _GEN_66;
  wire        _GEN_932 = _GEN_930 & _GEN_67;
  wire        _GEN_933 = _GEN_930 & _GEN_68;
  wire        _GEN_934 = _GEN_930 & _GEN_69;
  wire        _GEN_935 = _GEN_930 & _GEN_70;
  wire        _GEN_936 = _GEN_930 & _GEN_71;
  wire        _GEN_937 = _GEN_930 & _GEN_72;
  wire        _GEN_938 = _GEN_930 & _GEN_73;
  wire        _GEN_939 = _GEN_930 & _GEN_74;
  wire        _GEN_940 = _GEN_930 & _GEN_75;
  wire        _GEN_941 = _GEN_930 & _GEN_76;
  wire        _GEN_942 = _GEN_930 & _GEN_77;
  wire        _GEN_943 = _GEN_930 & _GEN_78;
  wire        _GEN_944 = _GEN_930 & _GEN_79;
  wire        _GEN_945 = _GEN_930 & _GEN_80;
  wire        _GEN_946 = _GEN_930 & _GEN_81;
  wire        _GEN_947 = _GEN_930 & _GEN_82;
  wire        _GEN_948 = _GEN_930 & _GEN_83;
  wire        _GEN_949 = _GEN_930 & _GEN_84;
  wire        _GEN_950 = _GEN_930 & _GEN_85;
  wire        _GEN_951 = _GEN_930 & _GEN_86;
  wire        _GEN_952 = _GEN_930 & _GEN_87;
  wire        _GEN_953 = _GEN_930 & _GEN_88;
  wire        _GEN_954 = _GEN_930 & _GEN_89;
  wire        _GEN_955 = _GEN_930 & _GEN_90;
  wire        _GEN_956 = _GEN_930 & _GEN_91;
  wire        _GEN_957 = _GEN_930 & _GEN_92;
  wire        _GEN_958 = _GEN_930 & _GEN_93;
  wire        _GEN_959 = _GEN_930 & _GEN_94;
  wire        _GEN_960 = _GEN_930 & _GEN_95;
  wire        _GEN_961 = _GEN_930 & _GEN_96;
  wire        _GEN_962 = _GEN_930 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_963 = io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_964 = _GEN_130 | _GEN_931;
  wire        _GEN_965 = _GEN_132 | _GEN_932;
  wire        _GEN_966 = _GEN_134 | _GEN_933;
  wire        _GEN_967 = _GEN_136 | _GEN_934;
  wire        _GEN_968 = _GEN_138 | _GEN_935;
  wire        _GEN_969 = _GEN_140 | _GEN_936;
  wire        _GEN_970 = _GEN_142 | _GEN_937;
  wire        _GEN_971 = _GEN_144 | _GEN_938;
  wire        _GEN_972 = _GEN_146 | _GEN_939;
  wire        _GEN_973 = _GEN_148 | _GEN_940;
  wire        _GEN_974 = _GEN_150 | _GEN_941;
  wire        _GEN_975 = _GEN_152 | _GEN_942;
  wire        _GEN_976 = _GEN_154 | _GEN_943;
  wire        _GEN_977 = _GEN_156 | _GEN_944;
  wire        _GEN_978 = _GEN_158 | _GEN_945;
  wire        _GEN_979 = _GEN_160 | _GEN_946;
  wire        _GEN_980 = _GEN_162 | _GEN_947;
  wire        _GEN_981 = _GEN_164 | _GEN_948;
  wire        _GEN_982 = _GEN_166 | _GEN_949;
  wire        _GEN_983 = _GEN_168 | _GEN_950;
  wire        _GEN_984 = _GEN_170 | _GEN_951;
  wire        _GEN_985 = _GEN_172 | _GEN_952;
  wire        _GEN_986 = _GEN_174 | _GEN_953;
  wire        _GEN_987 = _GEN_176 | _GEN_954;
  wire        _GEN_988 = _GEN_178 | _GEN_955;
  wire        _GEN_989 = _GEN_180 | _GEN_956;
  wire        _GEN_990 = _GEN_182 | _GEN_957;
  wire        _GEN_991 = _GEN_184 | _GEN_958;
  wire        _GEN_992 = _GEN_186 | _GEN_959;
  wire        _GEN_993 = _GEN_188 | _GEN_960;
  wire        _GEN_994 = _GEN_190 | _GEN_961;
  wire        _GEN_995 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_962;
  wire        _GEN_996 = io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_997 = _GEN_996 & _GEN_194;
  wire        _GEN_998 = _GEN_996 & _GEN_195;
  wire        _GEN_999 = _GEN_996 & _GEN_196;
  wire        _GEN_1000 = _GEN_996 & _GEN_197;
  wire        _GEN_1001 = _GEN_996 & _GEN_198;
  wire        _GEN_1002 = _GEN_996 & _GEN_199;
  wire        _GEN_1003 = _GEN_996 & _GEN_200;
  wire        _GEN_1004 = _GEN_996 & _GEN_201;
  wire        _GEN_1005 = _GEN_996 & _GEN_202;
  wire        _GEN_1006 = _GEN_996 & _GEN_203;
  wire        _GEN_1007 = _GEN_996 & _GEN_204;
  wire        _GEN_1008 = _GEN_996 & _GEN_205;
  wire        _GEN_1009 = _GEN_996 & _GEN_206;
  wire        _GEN_1010 = _GEN_996 & _GEN_207;
  wire        _GEN_1011 = _GEN_996 & _GEN_208;
  wire        _GEN_1012 = _GEN_996 & _GEN_209;
  wire        _GEN_1013 = _GEN_996 & _GEN_210;
  wire        _GEN_1014 = _GEN_996 & _GEN_211;
  wire        _GEN_1015 = _GEN_996 & _GEN_212;
  wire        _GEN_1016 = _GEN_996 & _GEN_213;
  wire        _GEN_1017 = _GEN_996 & _GEN_214;
  wire        _GEN_1018 = _GEN_996 & _GEN_215;
  wire        _GEN_1019 = _GEN_996 & _GEN_216;
  wire        _GEN_1020 = _GEN_996 & _GEN_217;
  wire        _GEN_1021 = _GEN_996 & _GEN_218;
  wire        _GEN_1022 = _GEN_996 & _GEN_219;
  wire        _GEN_1023 = _GEN_996 & _GEN_220;
  wire        _GEN_1024 = _GEN_996 & _GEN_221;
  wire        _GEN_1025 = _GEN_996 & _GEN_222;
  wire        _GEN_1026 = _GEN_996 & _GEN_223;
  wire        _GEN_1027 = _GEN_996 & _GEN_224;
  wire        _GEN_1028 = _GEN_996 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_1029 = io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_1030 = _GEN_258 | _GEN_997;
  wire        _GEN_1031 = _GEN_260 | _GEN_998;
  wire        _GEN_1032 = _GEN_262 | _GEN_999;
  wire        _GEN_1033 = _GEN_264 | _GEN_1000;
  wire        _GEN_1034 = _GEN_266 | _GEN_1001;
  wire        _GEN_1035 = _GEN_268 | _GEN_1002;
  wire        _GEN_1036 = _GEN_270 | _GEN_1003;
  wire        _GEN_1037 = _GEN_272 | _GEN_1004;
  wire        _GEN_1038 = _GEN_274 | _GEN_1005;
  wire        _GEN_1039 = _GEN_276 | _GEN_1006;
  wire        _GEN_1040 = _GEN_278 | _GEN_1007;
  wire        _GEN_1041 = _GEN_280 | _GEN_1008;
  wire        _GEN_1042 = _GEN_282 | _GEN_1009;
  wire        _GEN_1043 = _GEN_284 | _GEN_1010;
  wire        _GEN_1044 = _GEN_286 | _GEN_1011;
  wire        _GEN_1045 = _GEN_288 | _GEN_1012;
  wire        _GEN_1046 = _GEN_290 | _GEN_1013;
  wire        _GEN_1047 = _GEN_292 | _GEN_1014;
  wire        _GEN_1048 = _GEN_294 | _GEN_1015;
  wire        _GEN_1049 = _GEN_296 | _GEN_1016;
  wire        _GEN_1050 = _GEN_298 | _GEN_1017;
  wire        _GEN_1051 = _GEN_300 | _GEN_1018;
  wire        _GEN_1052 = _GEN_302 | _GEN_1019;
  wire        _GEN_1053 = _GEN_304 | _GEN_1020;
  wire        _GEN_1054 = _GEN_306 | _GEN_1021;
  wire        _GEN_1055 = _GEN_308 | _GEN_1022;
  wire        _GEN_1056 = _GEN_310 | _GEN_1023;
  wire        _GEN_1057 = _GEN_312 | _GEN_1024;
  wire        _GEN_1058 = _GEN_314 | _GEN_1025;
  wire        _GEN_1059 = _GEN_316 | _GEN_1026;
  wire        _GEN_1060 = _GEN_318 | _GEN_1027;
  wire        _GEN_1061 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1028;
  wire        _GEN_1062 = io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_1063 = _GEN_1062 & _GEN_322;
  wire        _GEN_1064 = _GEN_1062 & _GEN_323;
  wire        _GEN_1065 = _GEN_1062 & _GEN_324;
  wire        _GEN_1066 = _GEN_1062 & _GEN_325;
  wire        _GEN_1067 = _GEN_1062 & _GEN_326;
  wire        _GEN_1068 = _GEN_1062 & _GEN_327;
  wire        _GEN_1069 = _GEN_1062 & _GEN_328;
  wire        _GEN_1070 = _GEN_1062 & _GEN_329;
  wire        _GEN_1071 = _GEN_1062 & _GEN_330;
  wire        _GEN_1072 = _GEN_1062 & _GEN_331;
  wire        _GEN_1073 = _GEN_1062 & _GEN_332;
  wire        _GEN_1074 = _GEN_1062 & _GEN_333;
  wire        _GEN_1075 = _GEN_1062 & _GEN_334;
  wire        _GEN_1076 = _GEN_1062 & _GEN_335;
  wire        _GEN_1077 = _GEN_1062 & _GEN_336;
  wire        _GEN_1078 = _GEN_1062 & _GEN_337;
  wire        _GEN_1079 = _GEN_1062 & _GEN_338;
  wire        _GEN_1080 = _GEN_1062 & _GEN_339;
  wire        _GEN_1081 = _GEN_1062 & _GEN_340;
  wire        _GEN_1082 = _GEN_1062 & _GEN_341;
  wire        _GEN_1083 = _GEN_1062 & _GEN_342;
  wire        _GEN_1084 = _GEN_1062 & _GEN_343;
  wire        _GEN_1085 = _GEN_1062 & _GEN_344;
  wire        _GEN_1086 = _GEN_1062 & _GEN_345;
  wire        _GEN_1087 = _GEN_1062 & _GEN_346;
  wire        _GEN_1088 = _GEN_1062 & _GEN_347;
  wire        _GEN_1089 = _GEN_1062 & _GEN_348;
  wire        _GEN_1090 = _GEN_1062 & _GEN_349;
  wire        _GEN_1091 = _GEN_1062 & _GEN_350;
  wire        _GEN_1092 = _GEN_1062 & _GEN_351;
  wire        _GEN_1093 = _GEN_1062 & _GEN_352;
  wire        _GEN_1094 = _GEN_1062 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_1095 = io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_1096 = _GEN_386 | _GEN_1063;
  wire        _GEN_1097 = _GEN_388 | _GEN_1064;
  wire        _GEN_1098 = _GEN_390 | _GEN_1065;
  wire        _GEN_1099 = _GEN_392 | _GEN_1066;
  wire        _GEN_1100 = _GEN_394 | _GEN_1067;
  wire        _GEN_1101 = _GEN_396 | _GEN_1068;
  wire        _GEN_1102 = _GEN_398 | _GEN_1069;
  wire        _GEN_1103 = _GEN_400 | _GEN_1070;
  wire        _GEN_1104 = _GEN_402 | _GEN_1071;
  wire        _GEN_1105 = _GEN_404 | _GEN_1072;
  wire        _GEN_1106 = _GEN_406 | _GEN_1073;
  wire        _GEN_1107 = _GEN_408 | _GEN_1074;
  wire        _GEN_1108 = _GEN_410 | _GEN_1075;
  wire        _GEN_1109 = _GEN_412 | _GEN_1076;
  wire        _GEN_1110 = _GEN_414 | _GEN_1077;
  wire        _GEN_1111 = _GEN_416 | _GEN_1078;
  wire        _GEN_1112 = _GEN_418 | _GEN_1079;
  wire        _GEN_1113 = _GEN_420 | _GEN_1080;
  wire        _GEN_1114 = _GEN_422 | _GEN_1081;
  wire        _GEN_1115 = _GEN_424 | _GEN_1082;
  wire        _GEN_1116 = _GEN_426 | _GEN_1083;
  wire        _GEN_1117 = _GEN_428 | _GEN_1084;
  wire        _GEN_1118 = _GEN_430 | _GEN_1085;
  wire        _GEN_1119 = _GEN_432 | _GEN_1086;
  wire        _GEN_1120 = _GEN_434 | _GEN_1087;
  wire        _GEN_1121 = _GEN_436 | _GEN_1088;
  wire        _GEN_1122 = _GEN_438 | _GEN_1089;
  wire        _GEN_1123 = _GEN_440 | _GEN_1090;
  wire        _GEN_1124 = _GEN_442 | _GEN_1091;
  wire        _GEN_1125 = _GEN_444 | _GEN_1092;
  wire        _GEN_1126 = _GEN_446 | _GEN_1093;
  wire        _GEN_1127 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1094;
  wire        _GEN_1128 = io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_1129 = _GEN_1128 & _GEN_450;
  wire        _GEN_1130 = _GEN_1128 & _GEN_451;
  wire        _GEN_1131 = _GEN_1128 & _GEN_452;
  wire        _GEN_1132 = _GEN_1128 & _GEN_453;
  wire        _GEN_1133 = _GEN_1128 & _GEN_454;
  wire        _GEN_1134 = _GEN_1128 & _GEN_455;
  wire        _GEN_1135 = _GEN_1128 & _GEN_456;
  wire        _GEN_1136 = _GEN_1128 & _GEN_457;
  wire        _GEN_1137 = _GEN_1128 & _GEN_458;
  wire        _GEN_1138 = _GEN_1128 & _GEN_459;
  wire        _GEN_1139 = _GEN_1128 & _GEN_460;
  wire        _GEN_1140 = _GEN_1128 & _GEN_461;
  wire        _GEN_1141 = _GEN_1128 & _GEN_462;
  wire        _GEN_1142 = _GEN_1128 & _GEN_463;
  wire        _GEN_1143 = _GEN_1128 & _GEN_464;
  wire        _GEN_1144 = _GEN_1128 & _GEN_465;
  wire        _GEN_1145 = _GEN_1128 & _GEN_466;
  wire        _GEN_1146 = _GEN_1128 & _GEN_467;
  wire        _GEN_1147 = _GEN_1128 & _GEN_468;
  wire        _GEN_1148 = _GEN_1128 & _GEN_469;
  wire        _GEN_1149 = _GEN_1128 & _GEN_470;
  wire        _GEN_1150 = _GEN_1128 & _GEN_471;
  wire        _GEN_1151 = _GEN_1128 & _GEN_472;
  wire        _GEN_1152 = _GEN_1128 & _GEN_473;
  wire        _GEN_1153 = _GEN_1128 & _GEN_474;
  wire        _GEN_1154 = _GEN_1128 & _GEN_475;
  wire        _GEN_1155 = _GEN_1128 & _GEN_476;
  wire        _GEN_1156 = _GEN_1128 & _GEN_477;
  wire        _GEN_1157 = _GEN_1128 & _GEN_478;
  wire        _GEN_1158 = _GEN_1128 & _GEN_479;
  wire        _GEN_1159 = _GEN_1128 & _GEN_480;
  wire        _GEN_1160 = _GEN_1128 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_1161 = io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_1162 = _GEN_514 | _GEN_1129;
  wire        _GEN_1163 = _GEN_516 | _GEN_1130;
  wire        _GEN_1164 = _GEN_518 | _GEN_1131;
  wire        _GEN_1165 = _GEN_520 | _GEN_1132;
  wire        _GEN_1166 = _GEN_522 | _GEN_1133;
  wire        _GEN_1167 = _GEN_524 | _GEN_1134;
  wire        _GEN_1168 = _GEN_526 | _GEN_1135;
  wire        _GEN_1169 = _GEN_528 | _GEN_1136;
  wire        _GEN_1170 = _GEN_530 | _GEN_1137;
  wire        _GEN_1171 = _GEN_532 | _GEN_1138;
  wire        _GEN_1172 = _GEN_534 | _GEN_1139;
  wire        _GEN_1173 = _GEN_536 | _GEN_1140;
  wire        _GEN_1174 = _GEN_538 | _GEN_1141;
  wire        _GEN_1175 = _GEN_540 | _GEN_1142;
  wire        _GEN_1176 = _GEN_542 | _GEN_1143;
  wire        _GEN_1177 = _GEN_544 | _GEN_1144;
  wire        _GEN_1178 = _GEN_546 | _GEN_1145;
  wire        _GEN_1179 = _GEN_548 | _GEN_1146;
  wire        _GEN_1180 = _GEN_550 | _GEN_1147;
  wire        _GEN_1181 = _GEN_552 | _GEN_1148;
  wire        _GEN_1182 = _GEN_554 | _GEN_1149;
  wire        _GEN_1183 = _GEN_556 | _GEN_1150;
  wire        _GEN_1184 = _GEN_558 | _GEN_1151;
  wire        _GEN_1185 = _GEN_560 | _GEN_1152;
  wire        _GEN_1186 = _GEN_562 | _GEN_1153;
  wire        _GEN_1187 = _GEN_564 | _GEN_1154;
  wire        _GEN_1188 = _GEN_566 | _GEN_1155;
  wire        _GEN_1189 = _GEN_568 | _GEN_1156;
  wire        _GEN_1190 = _GEN_570 | _GEN_1157;
  wire        _GEN_1191 = _GEN_572 | _GEN_1158;
  wire        _GEN_1192 = _GEN_574 | _GEN_1159;
  wire        _GEN_1193 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_1160;
  wire        _GEN_1194 = io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_1195 = _GEN_1194 & _GEN_578;
  wire        _GEN_1196 = _GEN_1194 & _GEN_579;
  wire        _GEN_1197 = _GEN_1194 & _GEN_580;
  wire        _GEN_1198 = _GEN_1194 & _GEN_581;
  wire        _GEN_1199 = _GEN_1194 & _GEN_582;
  wire        _GEN_1200 = _GEN_1194 & _GEN_583;
  wire        _GEN_1201 = _GEN_1194 & _GEN_584;
  wire        _GEN_1202 = _GEN_1194 & _GEN_585;
  wire        _GEN_1203 = _GEN_1194 & _GEN_586;
  wire        _GEN_1204 = _GEN_1194 & _GEN_587;
  wire        _GEN_1205 = _GEN_1194 & _GEN_588;
  wire        _GEN_1206 = _GEN_1194 & _GEN_589;
  wire        _GEN_1207 = _GEN_1194 & _GEN_590;
  wire        _GEN_1208 = _GEN_1194 & _GEN_591;
  wire        _GEN_1209 = _GEN_1194 & _GEN_592;
  wire        _GEN_1210 = _GEN_1194 & _GEN_593;
  wire        _GEN_1211 = _GEN_1194 & _GEN_594;
  wire        _GEN_1212 = _GEN_1194 & _GEN_595;
  wire        _GEN_1213 = _GEN_1194 & _GEN_596;
  wire        _GEN_1214 = _GEN_1194 & _GEN_597;
  wire        _GEN_1215 = _GEN_1194 & _GEN_598;
  wire        _GEN_1216 = _GEN_1194 & _GEN_599;
  wire        _GEN_1217 = _GEN_1194 & _GEN_600;
  wire        _GEN_1218 = _GEN_1194 & _GEN_601;
  wire        _GEN_1219 = _GEN_1194 & _GEN_602;
  wire        _GEN_1220 = _GEN_1194 & _GEN_603;
  wire        _GEN_1221 = _GEN_1194 & _GEN_604;
  wire        _GEN_1222 = _GEN_1194 & _GEN_605;
  wire        _GEN_1223 = _GEN_1194 & _GEN_606;
  wire        _GEN_1224 = _GEN_1194 & _GEN_607;
  wire        _GEN_1225 = _GEN_1194 & _GEN_608;
  wire        _GEN_1226 = _GEN_1194 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_1227 = io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_1228 = _GEN_642 | _GEN_1195;
  wire        _GEN_1229 = _GEN_644 | _GEN_1196;
  wire        _GEN_1230 = _GEN_646 | _GEN_1197;
  wire        _GEN_1231 = _GEN_648 | _GEN_1198;
  wire        _GEN_1232 = _GEN_650 | _GEN_1199;
  wire        _GEN_1233 = _GEN_652 | _GEN_1200;
  wire        _GEN_1234 = _GEN_654 | _GEN_1201;
  wire        _GEN_1235 = _GEN_656 | _GEN_1202;
  wire        _GEN_1236 = _GEN_658 | _GEN_1203;
  wire        _GEN_1237 = _GEN_660 | _GEN_1204;
  wire        _GEN_1238 = _GEN_662 | _GEN_1205;
  wire        _GEN_1239 = _GEN_664 | _GEN_1206;
  wire        _GEN_1240 = _GEN_666 | _GEN_1207;
  wire        _GEN_1241 = _GEN_668 | _GEN_1208;
  wire        _GEN_1242 = _GEN_670 | _GEN_1209;
  wire        _GEN_1243 = _GEN_672 | _GEN_1210;
  wire        _GEN_1244 = _GEN_674 | _GEN_1211;
  wire        _GEN_1245 = _GEN_676 | _GEN_1212;
  wire        _GEN_1246 = _GEN_678 | _GEN_1213;
  wire        _GEN_1247 = _GEN_680 | _GEN_1214;
  wire        _GEN_1248 = _GEN_682 | _GEN_1215;
  wire        _GEN_1249 = _GEN_684 | _GEN_1216;
  wire        _GEN_1250 = _GEN_686 | _GEN_1217;
  wire        _GEN_1251 = _GEN_688 | _GEN_1218;
  wire        _GEN_1252 = _GEN_690 | _GEN_1219;
  wire        _GEN_1253 = _GEN_692 | _GEN_1220;
  wire        _GEN_1254 = _GEN_694 | _GEN_1221;
  wire        _GEN_1255 = _GEN_696 | _GEN_1222;
  wire        _GEN_1256 = _GEN_698 | _GEN_1223;
  wire        _GEN_1257 = _GEN_700 | _GEN_1224;
  wire        _GEN_1258 = _GEN_702 | _GEN_1225;
  wire        _GEN_1259 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1226;
  wire        _GEN_1260 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h1;
  wire        _GEN_1261 = _GEN_1260 & _GEN_706;
  wire        _GEN_1262 = _GEN_1260 & _GEN_707;
  wire        _GEN_1263 = _GEN_1260 & _GEN_708;
  wire        _GEN_1264 = _GEN_1260 & _GEN_709;
  wire        _GEN_1265 = _GEN_1260 & _GEN_710;
  wire        _GEN_1266 = _GEN_1260 & _GEN_711;
  wire        _GEN_1267 = _GEN_1260 & _GEN_712;
  wire        _GEN_1268 = _GEN_1260 & _GEN_713;
  wire        _GEN_1269 = _GEN_1260 & _GEN_714;
  wire        _GEN_1270 = _GEN_1260 & _GEN_715;
  wire        _GEN_1271 = _GEN_1260 & _GEN_716;
  wire        _GEN_1272 = _GEN_1260 & _GEN_717;
  wire        _GEN_1273 = _GEN_1260 & _GEN_718;
  wire        _GEN_1274 = _GEN_1260 & _GEN_719;
  wire        _GEN_1275 = _GEN_1260 & _GEN_720;
  wire        _GEN_1276 = _GEN_1260 & _GEN_721;
  wire        _GEN_1277 = _GEN_1260 & _GEN_722;
  wire        _GEN_1278 = _GEN_1260 & _GEN_723;
  wire        _GEN_1279 = _GEN_1260 & _GEN_724;
  wire        _GEN_1280 = _GEN_1260 & _GEN_725;
  wire        _GEN_1281 = _GEN_1260 & _GEN_726;
  wire        _GEN_1282 = _GEN_1260 & _GEN_727;
  wire        _GEN_1283 = _GEN_1260 & _GEN_728;
  wire        _GEN_1284 = _GEN_1260 & _GEN_729;
  wire        _GEN_1285 = _GEN_1260 & _GEN_730;
  wire        _GEN_1286 = _GEN_1260 & _GEN_731;
  wire        _GEN_1287 = _GEN_1260 & _GEN_732;
  wire        _GEN_1288 = _GEN_1260 & _GEN_733;
  wire        _GEN_1289 = _GEN_1260 & _GEN_734;
  wire        _GEN_1290 = _GEN_1260 & _GEN_735;
  wire        _GEN_1291 = _GEN_1260 & _GEN_736;
  wire        _GEN_1292 = _GEN_1260 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_1293 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h1;
  wire        _GEN_1294 = _GEN_770 | _GEN_1261;
  wire        _GEN_1295 = _GEN_772 | _GEN_1262;
  wire        _GEN_1296 = _GEN_774 | _GEN_1263;
  wire        _GEN_1297 = _GEN_776 | _GEN_1264;
  wire        _GEN_1298 = _GEN_778 | _GEN_1265;
  wire        _GEN_1299 = _GEN_780 | _GEN_1266;
  wire        _GEN_1300 = _GEN_782 | _GEN_1267;
  wire        _GEN_1301 = _GEN_784 | _GEN_1268;
  wire        _GEN_1302 = _GEN_786 | _GEN_1269;
  wire        _GEN_1303 = _GEN_788 | _GEN_1270;
  wire        _GEN_1304 = _GEN_790 | _GEN_1271;
  wire        _GEN_1305 = _GEN_792 | _GEN_1272;
  wire        _GEN_1306 = _GEN_794 | _GEN_1273;
  wire        _GEN_1307 = _GEN_796 | _GEN_1274;
  wire        _GEN_1308 = _GEN_798 | _GEN_1275;
  wire        _GEN_1309 = _GEN_800 | _GEN_1276;
  wire        _GEN_1310 = _GEN_802 | _GEN_1277;
  wire        _GEN_1311 = _GEN_804 | _GEN_1278;
  wire        _GEN_1312 = _GEN_806 | _GEN_1279;
  wire        _GEN_1313 = _GEN_808 | _GEN_1280;
  wire        _GEN_1314 = _GEN_810 | _GEN_1281;
  wire        _GEN_1315 = _GEN_812 | _GEN_1282;
  wire        _GEN_1316 = _GEN_814 | _GEN_1283;
  wire        _GEN_1317 = _GEN_816 | _GEN_1284;
  wire        _GEN_1318 = _GEN_818 | _GEN_1285;
  wire        _GEN_1319 = _GEN_820 | _GEN_1286;
  wire        _GEN_1320 = _GEN_822 | _GEN_1287;
  wire        _GEN_1321 = _GEN_824 | _GEN_1288;
  wire        _GEN_1322 = _GEN_826 | _GEN_1289;
  wire        _GEN_1323 = _GEN_828 | _GEN_1290;
  wire        _GEN_1324 = _GEN_830 | _GEN_1291;
  wire        _GEN_1325 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_1292;
  wire        _GEN_1326 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h1;
  wire        _GEN_1327 = _GEN_1326 & _GEN_834;
  wire        _GEN_1328 = _GEN_1326 & _GEN_835;
  wire        _GEN_1329 = _GEN_1326 & _GEN_836;
  wire        _GEN_1330 = _GEN_1326 & _GEN_837;
  wire        _GEN_1331 = _GEN_1326 & _GEN_838;
  wire        _GEN_1332 = _GEN_1326 & _GEN_839;
  wire        _GEN_1333 = _GEN_1326 & _GEN_840;
  wire        _GEN_1334 = _GEN_1326 & _GEN_841;
  wire        _GEN_1335 = _GEN_1326 & _GEN_842;
  wire        _GEN_1336 = _GEN_1326 & _GEN_843;
  wire        _GEN_1337 = _GEN_1326 & _GEN_844;
  wire        _GEN_1338 = _GEN_1326 & _GEN_845;
  wire        _GEN_1339 = _GEN_1326 & _GEN_846;
  wire        _GEN_1340 = _GEN_1326 & _GEN_847;
  wire        _GEN_1341 = _GEN_1326 & _GEN_848;
  wire        _GEN_1342 = _GEN_1326 & _GEN_849;
  wire        _GEN_1343 = _GEN_1326 & _GEN_850;
  wire        _GEN_1344 = _GEN_1326 & _GEN_851;
  wire        _GEN_1345 = _GEN_1326 & _GEN_852;
  wire        _GEN_1346 = _GEN_1326 & _GEN_853;
  wire        _GEN_1347 = _GEN_1326 & _GEN_854;
  wire        _GEN_1348 = _GEN_1326 & _GEN_855;
  wire        _GEN_1349 = _GEN_1326 & _GEN_856;
  wire        _GEN_1350 = _GEN_1326 & _GEN_857;
  wire        _GEN_1351 = _GEN_1326 & _GEN_858;
  wire        _GEN_1352 = _GEN_1326 & _GEN_859;
  wire        _GEN_1353 = _GEN_1326 & _GEN_860;
  wire        _GEN_1354 = _GEN_1326 & _GEN_861;
  wire        _GEN_1355 = _GEN_1326 & _GEN_862;
  wire        _GEN_1356 = _GEN_1326 & _GEN_863;
  wire        _GEN_1357 = _GEN_1326 & _GEN_864;
  wire        _GEN_1358 = _GEN_1326 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_1359 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h1;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_31 = rob_predicated_1_0;
      5'b00001:
        casez_tmp_31 = rob_predicated_1_1;
      5'b00010:
        casez_tmp_31 = rob_predicated_1_2;
      5'b00011:
        casez_tmp_31 = rob_predicated_1_3;
      5'b00100:
        casez_tmp_31 = rob_predicated_1_4;
      5'b00101:
        casez_tmp_31 = rob_predicated_1_5;
      5'b00110:
        casez_tmp_31 = rob_predicated_1_6;
      5'b00111:
        casez_tmp_31 = rob_predicated_1_7;
      5'b01000:
        casez_tmp_31 = rob_predicated_1_8;
      5'b01001:
        casez_tmp_31 = rob_predicated_1_9;
      5'b01010:
        casez_tmp_31 = rob_predicated_1_10;
      5'b01011:
        casez_tmp_31 = rob_predicated_1_11;
      5'b01100:
        casez_tmp_31 = rob_predicated_1_12;
      5'b01101:
        casez_tmp_31 = rob_predicated_1_13;
      5'b01110:
        casez_tmp_31 = rob_predicated_1_14;
      5'b01111:
        casez_tmp_31 = rob_predicated_1_15;
      5'b10000:
        casez_tmp_31 = rob_predicated_1_16;
      5'b10001:
        casez_tmp_31 = rob_predicated_1_17;
      5'b10010:
        casez_tmp_31 = rob_predicated_1_18;
      5'b10011:
        casez_tmp_31 = rob_predicated_1_19;
      5'b10100:
        casez_tmp_31 = rob_predicated_1_20;
      5'b10101:
        casez_tmp_31 = rob_predicated_1_21;
      5'b10110:
        casez_tmp_31 = rob_predicated_1_22;
      5'b10111:
        casez_tmp_31 = rob_predicated_1_23;
      5'b11000:
        casez_tmp_31 = rob_predicated_1_24;
      5'b11001:
        casez_tmp_31 = rob_predicated_1_25;
      5'b11010:
        casez_tmp_31 = rob_predicated_1_26;
      5'b11011:
        casez_tmp_31 = rob_predicated_1_27;
      5'b11100:
        casez_tmp_31 = rob_predicated_1_28;
      5'b11101:
        casez_tmp_31 = rob_predicated_1_29;
      5'b11110:
        casez_tmp_31 = rob_predicated_1_30;
      default:
        casez_tmp_31 = rob_predicated_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_32 = rob_uop_1_0_uopc;
      5'b00001:
        casez_tmp_32 = rob_uop_1_1_uopc;
      5'b00010:
        casez_tmp_32 = rob_uop_1_2_uopc;
      5'b00011:
        casez_tmp_32 = rob_uop_1_3_uopc;
      5'b00100:
        casez_tmp_32 = rob_uop_1_4_uopc;
      5'b00101:
        casez_tmp_32 = rob_uop_1_5_uopc;
      5'b00110:
        casez_tmp_32 = rob_uop_1_6_uopc;
      5'b00111:
        casez_tmp_32 = rob_uop_1_7_uopc;
      5'b01000:
        casez_tmp_32 = rob_uop_1_8_uopc;
      5'b01001:
        casez_tmp_32 = rob_uop_1_9_uopc;
      5'b01010:
        casez_tmp_32 = rob_uop_1_10_uopc;
      5'b01011:
        casez_tmp_32 = rob_uop_1_11_uopc;
      5'b01100:
        casez_tmp_32 = rob_uop_1_12_uopc;
      5'b01101:
        casez_tmp_32 = rob_uop_1_13_uopc;
      5'b01110:
        casez_tmp_32 = rob_uop_1_14_uopc;
      5'b01111:
        casez_tmp_32 = rob_uop_1_15_uopc;
      5'b10000:
        casez_tmp_32 = rob_uop_1_16_uopc;
      5'b10001:
        casez_tmp_32 = rob_uop_1_17_uopc;
      5'b10010:
        casez_tmp_32 = rob_uop_1_18_uopc;
      5'b10011:
        casez_tmp_32 = rob_uop_1_19_uopc;
      5'b10100:
        casez_tmp_32 = rob_uop_1_20_uopc;
      5'b10101:
        casez_tmp_32 = rob_uop_1_21_uopc;
      5'b10110:
        casez_tmp_32 = rob_uop_1_22_uopc;
      5'b10111:
        casez_tmp_32 = rob_uop_1_23_uopc;
      5'b11000:
        casez_tmp_32 = rob_uop_1_24_uopc;
      5'b11001:
        casez_tmp_32 = rob_uop_1_25_uopc;
      5'b11010:
        casez_tmp_32 = rob_uop_1_26_uopc;
      5'b11011:
        casez_tmp_32 = rob_uop_1_27_uopc;
      5'b11100:
        casez_tmp_32 = rob_uop_1_28_uopc;
      5'b11101:
        casez_tmp_32 = rob_uop_1_29_uopc;
      5'b11110:
        casez_tmp_32 = rob_uop_1_30_uopc;
      default:
        casez_tmp_32 = rob_uop_1_31_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_33 = rob_uop_1_0_is_rvc;
      5'b00001:
        casez_tmp_33 = rob_uop_1_1_is_rvc;
      5'b00010:
        casez_tmp_33 = rob_uop_1_2_is_rvc;
      5'b00011:
        casez_tmp_33 = rob_uop_1_3_is_rvc;
      5'b00100:
        casez_tmp_33 = rob_uop_1_4_is_rvc;
      5'b00101:
        casez_tmp_33 = rob_uop_1_5_is_rvc;
      5'b00110:
        casez_tmp_33 = rob_uop_1_6_is_rvc;
      5'b00111:
        casez_tmp_33 = rob_uop_1_7_is_rvc;
      5'b01000:
        casez_tmp_33 = rob_uop_1_8_is_rvc;
      5'b01001:
        casez_tmp_33 = rob_uop_1_9_is_rvc;
      5'b01010:
        casez_tmp_33 = rob_uop_1_10_is_rvc;
      5'b01011:
        casez_tmp_33 = rob_uop_1_11_is_rvc;
      5'b01100:
        casez_tmp_33 = rob_uop_1_12_is_rvc;
      5'b01101:
        casez_tmp_33 = rob_uop_1_13_is_rvc;
      5'b01110:
        casez_tmp_33 = rob_uop_1_14_is_rvc;
      5'b01111:
        casez_tmp_33 = rob_uop_1_15_is_rvc;
      5'b10000:
        casez_tmp_33 = rob_uop_1_16_is_rvc;
      5'b10001:
        casez_tmp_33 = rob_uop_1_17_is_rvc;
      5'b10010:
        casez_tmp_33 = rob_uop_1_18_is_rvc;
      5'b10011:
        casez_tmp_33 = rob_uop_1_19_is_rvc;
      5'b10100:
        casez_tmp_33 = rob_uop_1_20_is_rvc;
      5'b10101:
        casez_tmp_33 = rob_uop_1_21_is_rvc;
      5'b10110:
        casez_tmp_33 = rob_uop_1_22_is_rvc;
      5'b10111:
        casez_tmp_33 = rob_uop_1_23_is_rvc;
      5'b11000:
        casez_tmp_33 = rob_uop_1_24_is_rvc;
      5'b11001:
        casez_tmp_33 = rob_uop_1_25_is_rvc;
      5'b11010:
        casez_tmp_33 = rob_uop_1_26_is_rvc;
      5'b11011:
        casez_tmp_33 = rob_uop_1_27_is_rvc;
      5'b11100:
        casez_tmp_33 = rob_uop_1_28_is_rvc;
      5'b11101:
        casez_tmp_33 = rob_uop_1_29_is_rvc;
      5'b11110:
        casez_tmp_33 = rob_uop_1_30_is_rvc;
      default:
        casez_tmp_33 = rob_uop_1_31_is_rvc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_34 = rob_uop_1_0_ftq_idx;
      5'b00001:
        casez_tmp_34 = rob_uop_1_1_ftq_idx;
      5'b00010:
        casez_tmp_34 = rob_uop_1_2_ftq_idx;
      5'b00011:
        casez_tmp_34 = rob_uop_1_3_ftq_idx;
      5'b00100:
        casez_tmp_34 = rob_uop_1_4_ftq_idx;
      5'b00101:
        casez_tmp_34 = rob_uop_1_5_ftq_idx;
      5'b00110:
        casez_tmp_34 = rob_uop_1_6_ftq_idx;
      5'b00111:
        casez_tmp_34 = rob_uop_1_7_ftq_idx;
      5'b01000:
        casez_tmp_34 = rob_uop_1_8_ftq_idx;
      5'b01001:
        casez_tmp_34 = rob_uop_1_9_ftq_idx;
      5'b01010:
        casez_tmp_34 = rob_uop_1_10_ftq_idx;
      5'b01011:
        casez_tmp_34 = rob_uop_1_11_ftq_idx;
      5'b01100:
        casez_tmp_34 = rob_uop_1_12_ftq_idx;
      5'b01101:
        casez_tmp_34 = rob_uop_1_13_ftq_idx;
      5'b01110:
        casez_tmp_34 = rob_uop_1_14_ftq_idx;
      5'b01111:
        casez_tmp_34 = rob_uop_1_15_ftq_idx;
      5'b10000:
        casez_tmp_34 = rob_uop_1_16_ftq_idx;
      5'b10001:
        casez_tmp_34 = rob_uop_1_17_ftq_idx;
      5'b10010:
        casez_tmp_34 = rob_uop_1_18_ftq_idx;
      5'b10011:
        casez_tmp_34 = rob_uop_1_19_ftq_idx;
      5'b10100:
        casez_tmp_34 = rob_uop_1_20_ftq_idx;
      5'b10101:
        casez_tmp_34 = rob_uop_1_21_ftq_idx;
      5'b10110:
        casez_tmp_34 = rob_uop_1_22_ftq_idx;
      5'b10111:
        casez_tmp_34 = rob_uop_1_23_ftq_idx;
      5'b11000:
        casez_tmp_34 = rob_uop_1_24_ftq_idx;
      5'b11001:
        casez_tmp_34 = rob_uop_1_25_ftq_idx;
      5'b11010:
        casez_tmp_34 = rob_uop_1_26_ftq_idx;
      5'b11011:
        casez_tmp_34 = rob_uop_1_27_ftq_idx;
      5'b11100:
        casez_tmp_34 = rob_uop_1_28_ftq_idx;
      5'b11101:
        casez_tmp_34 = rob_uop_1_29_ftq_idx;
      5'b11110:
        casez_tmp_34 = rob_uop_1_30_ftq_idx;
      default:
        casez_tmp_34 = rob_uop_1_31_ftq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_35 = rob_uop_1_0_edge_inst;
      5'b00001:
        casez_tmp_35 = rob_uop_1_1_edge_inst;
      5'b00010:
        casez_tmp_35 = rob_uop_1_2_edge_inst;
      5'b00011:
        casez_tmp_35 = rob_uop_1_3_edge_inst;
      5'b00100:
        casez_tmp_35 = rob_uop_1_4_edge_inst;
      5'b00101:
        casez_tmp_35 = rob_uop_1_5_edge_inst;
      5'b00110:
        casez_tmp_35 = rob_uop_1_6_edge_inst;
      5'b00111:
        casez_tmp_35 = rob_uop_1_7_edge_inst;
      5'b01000:
        casez_tmp_35 = rob_uop_1_8_edge_inst;
      5'b01001:
        casez_tmp_35 = rob_uop_1_9_edge_inst;
      5'b01010:
        casez_tmp_35 = rob_uop_1_10_edge_inst;
      5'b01011:
        casez_tmp_35 = rob_uop_1_11_edge_inst;
      5'b01100:
        casez_tmp_35 = rob_uop_1_12_edge_inst;
      5'b01101:
        casez_tmp_35 = rob_uop_1_13_edge_inst;
      5'b01110:
        casez_tmp_35 = rob_uop_1_14_edge_inst;
      5'b01111:
        casez_tmp_35 = rob_uop_1_15_edge_inst;
      5'b10000:
        casez_tmp_35 = rob_uop_1_16_edge_inst;
      5'b10001:
        casez_tmp_35 = rob_uop_1_17_edge_inst;
      5'b10010:
        casez_tmp_35 = rob_uop_1_18_edge_inst;
      5'b10011:
        casez_tmp_35 = rob_uop_1_19_edge_inst;
      5'b10100:
        casez_tmp_35 = rob_uop_1_20_edge_inst;
      5'b10101:
        casez_tmp_35 = rob_uop_1_21_edge_inst;
      5'b10110:
        casez_tmp_35 = rob_uop_1_22_edge_inst;
      5'b10111:
        casez_tmp_35 = rob_uop_1_23_edge_inst;
      5'b11000:
        casez_tmp_35 = rob_uop_1_24_edge_inst;
      5'b11001:
        casez_tmp_35 = rob_uop_1_25_edge_inst;
      5'b11010:
        casez_tmp_35 = rob_uop_1_26_edge_inst;
      5'b11011:
        casez_tmp_35 = rob_uop_1_27_edge_inst;
      5'b11100:
        casez_tmp_35 = rob_uop_1_28_edge_inst;
      5'b11101:
        casez_tmp_35 = rob_uop_1_29_edge_inst;
      5'b11110:
        casez_tmp_35 = rob_uop_1_30_edge_inst;
      default:
        casez_tmp_35 = rob_uop_1_31_edge_inst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_36 = rob_uop_1_0_pc_lob;
      5'b00001:
        casez_tmp_36 = rob_uop_1_1_pc_lob;
      5'b00010:
        casez_tmp_36 = rob_uop_1_2_pc_lob;
      5'b00011:
        casez_tmp_36 = rob_uop_1_3_pc_lob;
      5'b00100:
        casez_tmp_36 = rob_uop_1_4_pc_lob;
      5'b00101:
        casez_tmp_36 = rob_uop_1_5_pc_lob;
      5'b00110:
        casez_tmp_36 = rob_uop_1_6_pc_lob;
      5'b00111:
        casez_tmp_36 = rob_uop_1_7_pc_lob;
      5'b01000:
        casez_tmp_36 = rob_uop_1_8_pc_lob;
      5'b01001:
        casez_tmp_36 = rob_uop_1_9_pc_lob;
      5'b01010:
        casez_tmp_36 = rob_uop_1_10_pc_lob;
      5'b01011:
        casez_tmp_36 = rob_uop_1_11_pc_lob;
      5'b01100:
        casez_tmp_36 = rob_uop_1_12_pc_lob;
      5'b01101:
        casez_tmp_36 = rob_uop_1_13_pc_lob;
      5'b01110:
        casez_tmp_36 = rob_uop_1_14_pc_lob;
      5'b01111:
        casez_tmp_36 = rob_uop_1_15_pc_lob;
      5'b10000:
        casez_tmp_36 = rob_uop_1_16_pc_lob;
      5'b10001:
        casez_tmp_36 = rob_uop_1_17_pc_lob;
      5'b10010:
        casez_tmp_36 = rob_uop_1_18_pc_lob;
      5'b10011:
        casez_tmp_36 = rob_uop_1_19_pc_lob;
      5'b10100:
        casez_tmp_36 = rob_uop_1_20_pc_lob;
      5'b10101:
        casez_tmp_36 = rob_uop_1_21_pc_lob;
      5'b10110:
        casez_tmp_36 = rob_uop_1_22_pc_lob;
      5'b10111:
        casez_tmp_36 = rob_uop_1_23_pc_lob;
      5'b11000:
        casez_tmp_36 = rob_uop_1_24_pc_lob;
      5'b11001:
        casez_tmp_36 = rob_uop_1_25_pc_lob;
      5'b11010:
        casez_tmp_36 = rob_uop_1_26_pc_lob;
      5'b11011:
        casez_tmp_36 = rob_uop_1_27_pc_lob;
      5'b11100:
        casez_tmp_36 = rob_uop_1_28_pc_lob;
      5'b11101:
        casez_tmp_36 = rob_uop_1_29_pc_lob;
      5'b11110:
        casez_tmp_36 = rob_uop_1_30_pc_lob;
      default:
        casez_tmp_36 = rob_uop_1_31_pc_lob;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_37 = rob_uop_1_0_pdst;
      5'b00001:
        casez_tmp_37 = rob_uop_1_1_pdst;
      5'b00010:
        casez_tmp_37 = rob_uop_1_2_pdst;
      5'b00011:
        casez_tmp_37 = rob_uop_1_3_pdst;
      5'b00100:
        casez_tmp_37 = rob_uop_1_4_pdst;
      5'b00101:
        casez_tmp_37 = rob_uop_1_5_pdst;
      5'b00110:
        casez_tmp_37 = rob_uop_1_6_pdst;
      5'b00111:
        casez_tmp_37 = rob_uop_1_7_pdst;
      5'b01000:
        casez_tmp_37 = rob_uop_1_8_pdst;
      5'b01001:
        casez_tmp_37 = rob_uop_1_9_pdst;
      5'b01010:
        casez_tmp_37 = rob_uop_1_10_pdst;
      5'b01011:
        casez_tmp_37 = rob_uop_1_11_pdst;
      5'b01100:
        casez_tmp_37 = rob_uop_1_12_pdst;
      5'b01101:
        casez_tmp_37 = rob_uop_1_13_pdst;
      5'b01110:
        casez_tmp_37 = rob_uop_1_14_pdst;
      5'b01111:
        casez_tmp_37 = rob_uop_1_15_pdst;
      5'b10000:
        casez_tmp_37 = rob_uop_1_16_pdst;
      5'b10001:
        casez_tmp_37 = rob_uop_1_17_pdst;
      5'b10010:
        casez_tmp_37 = rob_uop_1_18_pdst;
      5'b10011:
        casez_tmp_37 = rob_uop_1_19_pdst;
      5'b10100:
        casez_tmp_37 = rob_uop_1_20_pdst;
      5'b10101:
        casez_tmp_37 = rob_uop_1_21_pdst;
      5'b10110:
        casez_tmp_37 = rob_uop_1_22_pdst;
      5'b10111:
        casez_tmp_37 = rob_uop_1_23_pdst;
      5'b11000:
        casez_tmp_37 = rob_uop_1_24_pdst;
      5'b11001:
        casez_tmp_37 = rob_uop_1_25_pdst;
      5'b11010:
        casez_tmp_37 = rob_uop_1_26_pdst;
      5'b11011:
        casez_tmp_37 = rob_uop_1_27_pdst;
      5'b11100:
        casez_tmp_37 = rob_uop_1_28_pdst;
      5'b11101:
        casez_tmp_37 = rob_uop_1_29_pdst;
      5'b11110:
        casez_tmp_37 = rob_uop_1_30_pdst;
      default:
        casez_tmp_37 = rob_uop_1_31_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_38 = rob_uop_1_0_stale_pdst;
      5'b00001:
        casez_tmp_38 = rob_uop_1_1_stale_pdst;
      5'b00010:
        casez_tmp_38 = rob_uop_1_2_stale_pdst;
      5'b00011:
        casez_tmp_38 = rob_uop_1_3_stale_pdst;
      5'b00100:
        casez_tmp_38 = rob_uop_1_4_stale_pdst;
      5'b00101:
        casez_tmp_38 = rob_uop_1_5_stale_pdst;
      5'b00110:
        casez_tmp_38 = rob_uop_1_6_stale_pdst;
      5'b00111:
        casez_tmp_38 = rob_uop_1_7_stale_pdst;
      5'b01000:
        casez_tmp_38 = rob_uop_1_8_stale_pdst;
      5'b01001:
        casez_tmp_38 = rob_uop_1_9_stale_pdst;
      5'b01010:
        casez_tmp_38 = rob_uop_1_10_stale_pdst;
      5'b01011:
        casez_tmp_38 = rob_uop_1_11_stale_pdst;
      5'b01100:
        casez_tmp_38 = rob_uop_1_12_stale_pdst;
      5'b01101:
        casez_tmp_38 = rob_uop_1_13_stale_pdst;
      5'b01110:
        casez_tmp_38 = rob_uop_1_14_stale_pdst;
      5'b01111:
        casez_tmp_38 = rob_uop_1_15_stale_pdst;
      5'b10000:
        casez_tmp_38 = rob_uop_1_16_stale_pdst;
      5'b10001:
        casez_tmp_38 = rob_uop_1_17_stale_pdst;
      5'b10010:
        casez_tmp_38 = rob_uop_1_18_stale_pdst;
      5'b10011:
        casez_tmp_38 = rob_uop_1_19_stale_pdst;
      5'b10100:
        casez_tmp_38 = rob_uop_1_20_stale_pdst;
      5'b10101:
        casez_tmp_38 = rob_uop_1_21_stale_pdst;
      5'b10110:
        casez_tmp_38 = rob_uop_1_22_stale_pdst;
      5'b10111:
        casez_tmp_38 = rob_uop_1_23_stale_pdst;
      5'b11000:
        casez_tmp_38 = rob_uop_1_24_stale_pdst;
      5'b11001:
        casez_tmp_38 = rob_uop_1_25_stale_pdst;
      5'b11010:
        casez_tmp_38 = rob_uop_1_26_stale_pdst;
      5'b11011:
        casez_tmp_38 = rob_uop_1_27_stale_pdst;
      5'b11100:
        casez_tmp_38 = rob_uop_1_28_stale_pdst;
      5'b11101:
        casez_tmp_38 = rob_uop_1_29_stale_pdst;
      5'b11110:
        casez_tmp_38 = rob_uop_1_30_stale_pdst;
      default:
        casez_tmp_38 = rob_uop_1_31_stale_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_39 = rob_uop_1_0_is_fencei;
      5'b00001:
        casez_tmp_39 = rob_uop_1_1_is_fencei;
      5'b00010:
        casez_tmp_39 = rob_uop_1_2_is_fencei;
      5'b00011:
        casez_tmp_39 = rob_uop_1_3_is_fencei;
      5'b00100:
        casez_tmp_39 = rob_uop_1_4_is_fencei;
      5'b00101:
        casez_tmp_39 = rob_uop_1_5_is_fencei;
      5'b00110:
        casez_tmp_39 = rob_uop_1_6_is_fencei;
      5'b00111:
        casez_tmp_39 = rob_uop_1_7_is_fencei;
      5'b01000:
        casez_tmp_39 = rob_uop_1_8_is_fencei;
      5'b01001:
        casez_tmp_39 = rob_uop_1_9_is_fencei;
      5'b01010:
        casez_tmp_39 = rob_uop_1_10_is_fencei;
      5'b01011:
        casez_tmp_39 = rob_uop_1_11_is_fencei;
      5'b01100:
        casez_tmp_39 = rob_uop_1_12_is_fencei;
      5'b01101:
        casez_tmp_39 = rob_uop_1_13_is_fencei;
      5'b01110:
        casez_tmp_39 = rob_uop_1_14_is_fencei;
      5'b01111:
        casez_tmp_39 = rob_uop_1_15_is_fencei;
      5'b10000:
        casez_tmp_39 = rob_uop_1_16_is_fencei;
      5'b10001:
        casez_tmp_39 = rob_uop_1_17_is_fencei;
      5'b10010:
        casez_tmp_39 = rob_uop_1_18_is_fencei;
      5'b10011:
        casez_tmp_39 = rob_uop_1_19_is_fencei;
      5'b10100:
        casez_tmp_39 = rob_uop_1_20_is_fencei;
      5'b10101:
        casez_tmp_39 = rob_uop_1_21_is_fencei;
      5'b10110:
        casez_tmp_39 = rob_uop_1_22_is_fencei;
      5'b10111:
        casez_tmp_39 = rob_uop_1_23_is_fencei;
      5'b11000:
        casez_tmp_39 = rob_uop_1_24_is_fencei;
      5'b11001:
        casez_tmp_39 = rob_uop_1_25_is_fencei;
      5'b11010:
        casez_tmp_39 = rob_uop_1_26_is_fencei;
      5'b11011:
        casez_tmp_39 = rob_uop_1_27_is_fencei;
      5'b11100:
        casez_tmp_39 = rob_uop_1_28_is_fencei;
      5'b11101:
        casez_tmp_39 = rob_uop_1_29_is_fencei;
      5'b11110:
        casez_tmp_39 = rob_uop_1_30_is_fencei;
      default:
        casez_tmp_39 = rob_uop_1_31_is_fencei;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_40 = rob_uop_1_0_uses_ldq;
      5'b00001:
        casez_tmp_40 = rob_uop_1_1_uses_ldq;
      5'b00010:
        casez_tmp_40 = rob_uop_1_2_uses_ldq;
      5'b00011:
        casez_tmp_40 = rob_uop_1_3_uses_ldq;
      5'b00100:
        casez_tmp_40 = rob_uop_1_4_uses_ldq;
      5'b00101:
        casez_tmp_40 = rob_uop_1_5_uses_ldq;
      5'b00110:
        casez_tmp_40 = rob_uop_1_6_uses_ldq;
      5'b00111:
        casez_tmp_40 = rob_uop_1_7_uses_ldq;
      5'b01000:
        casez_tmp_40 = rob_uop_1_8_uses_ldq;
      5'b01001:
        casez_tmp_40 = rob_uop_1_9_uses_ldq;
      5'b01010:
        casez_tmp_40 = rob_uop_1_10_uses_ldq;
      5'b01011:
        casez_tmp_40 = rob_uop_1_11_uses_ldq;
      5'b01100:
        casez_tmp_40 = rob_uop_1_12_uses_ldq;
      5'b01101:
        casez_tmp_40 = rob_uop_1_13_uses_ldq;
      5'b01110:
        casez_tmp_40 = rob_uop_1_14_uses_ldq;
      5'b01111:
        casez_tmp_40 = rob_uop_1_15_uses_ldq;
      5'b10000:
        casez_tmp_40 = rob_uop_1_16_uses_ldq;
      5'b10001:
        casez_tmp_40 = rob_uop_1_17_uses_ldq;
      5'b10010:
        casez_tmp_40 = rob_uop_1_18_uses_ldq;
      5'b10011:
        casez_tmp_40 = rob_uop_1_19_uses_ldq;
      5'b10100:
        casez_tmp_40 = rob_uop_1_20_uses_ldq;
      5'b10101:
        casez_tmp_40 = rob_uop_1_21_uses_ldq;
      5'b10110:
        casez_tmp_40 = rob_uop_1_22_uses_ldq;
      5'b10111:
        casez_tmp_40 = rob_uop_1_23_uses_ldq;
      5'b11000:
        casez_tmp_40 = rob_uop_1_24_uses_ldq;
      5'b11001:
        casez_tmp_40 = rob_uop_1_25_uses_ldq;
      5'b11010:
        casez_tmp_40 = rob_uop_1_26_uses_ldq;
      5'b11011:
        casez_tmp_40 = rob_uop_1_27_uses_ldq;
      5'b11100:
        casez_tmp_40 = rob_uop_1_28_uses_ldq;
      5'b11101:
        casez_tmp_40 = rob_uop_1_29_uses_ldq;
      5'b11110:
        casez_tmp_40 = rob_uop_1_30_uses_ldq;
      default:
        casez_tmp_40 = rob_uop_1_31_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_41 = rob_uop_1_0_uses_stq;
      5'b00001:
        casez_tmp_41 = rob_uop_1_1_uses_stq;
      5'b00010:
        casez_tmp_41 = rob_uop_1_2_uses_stq;
      5'b00011:
        casez_tmp_41 = rob_uop_1_3_uses_stq;
      5'b00100:
        casez_tmp_41 = rob_uop_1_4_uses_stq;
      5'b00101:
        casez_tmp_41 = rob_uop_1_5_uses_stq;
      5'b00110:
        casez_tmp_41 = rob_uop_1_6_uses_stq;
      5'b00111:
        casez_tmp_41 = rob_uop_1_7_uses_stq;
      5'b01000:
        casez_tmp_41 = rob_uop_1_8_uses_stq;
      5'b01001:
        casez_tmp_41 = rob_uop_1_9_uses_stq;
      5'b01010:
        casez_tmp_41 = rob_uop_1_10_uses_stq;
      5'b01011:
        casez_tmp_41 = rob_uop_1_11_uses_stq;
      5'b01100:
        casez_tmp_41 = rob_uop_1_12_uses_stq;
      5'b01101:
        casez_tmp_41 = rob_uop_1_13_uses_stq;
      5'b01110:
        casez_tmp_41 = rob_uop_1_14_uses_stq;
      5'b01111:
        casez_tmp_41 = rob_uop_1_15_uses_stq;
      5'b10000:
        casez_tmp_41 = rob_uop_1_16_uses_stq;
      5'b10001:
        casez_tmp_41 = rob_uop_1_17_uses_stq;
      5'b10010:
        casez_tmp_41 = rob_uop_1_18_uses_stq;
      5'b10011:
        casez_tmp_41 = rob_uop_1_19_uses_stq;
      5'b10100:
        casez_tmp_41 = rob_uop_1_20_uses_stq;
      5'b10101:
        casez_tmp_41 = rob_uop_1_21_uses_stq;
      5'b10110:
        casez_tmp_41 = rob_uop_1_22_uses_stq;
      5'b10111:
        casez_tmp_41 = rob_uop_1_23_uses_stq;
      5'b11000:
        casez_tmp_41 = rob_uop_1_24_uses_stq;
      5'b11001:
        casez_tmp_41 = rob_uop_1_25_uses_stq;
      5'b11010:
        casez_tmp_41 = rob_uop_1_26_uses_stq;
      5'b11011:
        casez_tmp_41 = rob_uop_1_27_uses_stq;
      5'b11100:
        casez_tmp_41 = rob_uop_1_28_uses_stq;
      5'b11101:
        casez_tmp_41 = rob_uop_1_29_uses_stq;
      5'b11110:
        casez_tmp_41 = rob_uop_1_30_uses_stq;
      default:
        casez_tmp_41 = rob_uop_1_31_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_42 = rob_uop_1_0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_42 = rob_uop_1_1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_42 = rob_uop_1_2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_42 = rob_uop_1_3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_42 = rob_uop_1_4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_42 = rob_uop_1_5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_42 = rob_uop_1_6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_42 = rob_uop_1_7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_42 = rob_uop_1_8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_42 = rob_uop_1_9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_42 = rob_uop_1_10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_42 = rob_uop_1_11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_42 = rob_uop_1_12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_42 = rob_uop_1_13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_42 = rob_uop_1_14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_42 = rob_uop_1_15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_42 = rob_uop_1_16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_42 = rob_uop_1_17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_42 = rob_uop_1_18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_42 = rob_uop_1_19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_42 = rob_uop_1_20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_42 = rob_uop_1_21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_42 = rob_uop_1_22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_42 = rob_uop_1_23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_42 = rob_uop_1_24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_42 = rob_uop_1_25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_42 = rob_uop_1_26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_42 = rob_uop_1_27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_42 = rob_uop_1_28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_42 = rob_uop_1_29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_42 = rob_uop_1_30_is_sys_pc2epc;
      default:
        casez_tmp_42 = rob_uop_1_31_is_sys_pc2epc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_43 = rob_uop_1_0_flush_on_commit;
      5'b00001:
        casez_tmp_43 = rob_uop_1_1_flush_on_commit;
      5'b00010:
        casez_tmp_43 = rob_uop_1_2_flush_on_commit;
      5'b00011:
        casez_tmp_43 = rob_uop_1_3_flush_on_commit;
      5'b00100:
        casez_tmp_43 = rob_uop_1_4_flush_on_commit;
      5'b00101:
        casez_tmp_43 = rob_uop_1_5_flush_on_commit;
      5'b00110:
        casez_tmp_43 = rob_uop_1_6_flush_on_commit;
      5'b00111:
        casez_tmp_43 = rob_uop_1_7_flush_on_commit;
      5'b01000:
        casez_tmp_43 = rob_uop_1_8_flush_on_commit;
      5'b01001:
        casez_tmp_43 = rob_uop_1_9_flush_on_commit;
      5'b01010:
        casez_tmp_43 = rob_uop_1_10_flush_on_commit;
      5'b01011:
        casez_tmp_43 = rob_uop_1_11_flush_on_commit;
      5'b01100:
        casez_tmp_43 = rob_uop_1_12_flush_on_commit;
      5'b01101:
        casez_tmp_43 = rob_uop_1_13_flush_on_commit;
      5'b01110:
        casez_tmp_43 = rob_uop_1_14_flush_on_commit;
      5'b01111:
        casez_tmp_43 = rob_uop_1_15_flush_on_commit;
      5'b10000:
        casez_tmp_43 = rob_uop_1_16_flush_on_commit;
      5'b10001:
        casez_tmp_43 = rob_uop_1_17_flush_on_commit;
      5'b10010:
        casez_tmp_43 = rob_uop_1_18_flush_on_commit;
      5'b10011:
        casez_tmp_43 = rob_uop_1_19_flush_on_commit;
      5'b10100:
        casez_tmp_43 = rob_uop_1_20_flush_on_commit;
      5'b10101:
        casez_tmp_43 = rob_uop_1_21_flush_on_commit;
      5'b10110:
        casez_tmp_43 = rob_uop_1_22_flush_on_commit;
      5'b10111:
        casez_tmp_43 = rob_uop_1_23_flush_on_commit;
      5'b11000:
        casez_tmp_43 = rob_uop_1_24_flush_on_commit;
      5'b11001:
        casez_tmp_43 = rob_uop_1_25_flush_on_commit;
      5'b11010:
        casez_tmp_43 = rob_uop_1_26_flush_on_commit;
      5'b11011:
        casez_tmp_43 = rob_uop_1_27_flush_on_commit;
      5'b11100:
        casez_tmp_43 = rob_uop_1_28_flush_on_commit;
      5'b11101:
        casez_tmp_43 = rob_uop_1_29_flush_on_commit;
      5'b11110:
        casez_tmp_43 = rob_uop_1_30_flush_on_commit;
      default:
        casez_tmp_43 = rob_uop_1_31_flush_on_commit;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_44 = rob_uop_1_0_ldst;
      5'b00001:
        casez_tmp_44 = rob_uop_1_1_ldst;
      5'b00010:
        casez_tmp_44 = rob_uop_1_2_ldst;
      5'b00011:
        casez_tmp_44 = rob_uop_1_3_ldst;
      5'b00100:
        casez_tmp_44 = rob_uop_1_4_ldst;
      5'b00101:
        casez_tmp_44 = rob_uop_1_5_ldst;
      5'b00110:
        casez_tmp_44 = rob_uop_1_6_ldst;
      5'b00111:
        casez_tmp_44 = rob_uop_1_7_ldst;
      5'b01000:
        casez_tmp_44 = rob_uop_1_8_ldst;
      5'b01001:
        casez_tmp_44 = rob_uop_1_9_ldst;
      5'b01010:
        casez_tmp_44 = rob_uop_1_10_ldst;
      5'b01011:
        casez_tmp_44 = rob_uop_1_11_ldst;
      5'b01100:
        casez_tmp_44 = rob_uop_1_12_ldst;
      5'b01101:
        casez_tmp_44 = rob_uop_1_13_ldst;
      5'b01110:
        casez_tmp_44 = rob_uop_1_14_ldst;
      5'b01111:
        casez_tmp_44 = rob_uop_1_15_ldst;
      5'b10000:
        casez_tmp_44 = rob_uop_1_16_ldst;
      5'b10001:
        casez_tmp_44 = rob_uop_1_17_ldst;
      5'b10010:
        casez_tmp_44 = rob_uop_1_18_ldst;
      5'b10011:
        casez_tmp_44 = rob_uop_1_19_ldst;
      5'b10100:
        casez_tmp_44 = rob_uop_1_20_ldst;
      5'b10101:
        casez_tmp_44 = rob_uop_1_21_ldst;
      5'b10110:
        casez_tmp_44 = rob_uop_1_22_ldst;
      5'b10111:
        casez_tmp_44 = rob_uop_1_23_ldst;
      5'b11000:
        casez_tmp_44 = rob_uop_1_24_ldst;
      5'b11001:
        casez_tmp_44 = rob_uop_1_25_ldst;
      5'b11010:
        casez_tmp_44 = rob_uop_1_26_ldst;
      5'b11011:
        casez_tmp_44 = rob_uop_1_27_ldst;
      5'b11100:
        casez_tmp_44 = rob_uop_1_28_ldst;
      5'b11101:
        casez_tmp_44 = rob_uop_1_29_ldst;
      5'b11110:
        casez_tmp_44 = rob_uop_1_30_ldst;
      default:
        casez_tmp_44 = rob_uop_1_31_ldst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_45 = rob_uop_1_0_ldst_val;
      5'b00001:
        casez_tmp_45 = rob_uop_1_1_ldst_val;
      5'b00010:
        casez_tmp_45 = rob_uop_1_2_ldst_val;
      5'b00011:
        casez_tmp_45 = rob_uop_1_3_ldst_val;
      5'b00100:
        casez_tmp_45 = rob_uop_1_4_ldst_val;
      5'b00101:
        casez_tmp_45 = rob_uop_1_5_ldst_val;
      5'b00110:
        casez_tmp_45 = rob_uop_1_6_ldst_val;
      5'b00111:
        casez_tmp_45 = rob_uop_1_7_ldst_val;
      5'b01000:
        casez_tmp_45 = rob_uop_1_8_ldst_val;
      5'b01001:
        casez_tmp_45 = rob_uop_1_9_ldst_val;
      5'b01010:
        casez_tmp_45 = rob_uop_1_10_ldst_val;
      5'b01011:
        casez_tmp_45 = rob_uop_1_11_ldst_val;
      5'b01100:
        casez_tmp_45 = rob_uop_1_12_ldst_val;
      5'b01101:
        casez_tmp_45 = rob_uop_1_13_ldst_val;
      5'b01110:
        casez_tmp_45 = rob_uop_1_14_ldst_val;
      5'b01111:
        casez_tmp_45 = rob_uop_1_15_ldst_val;
      5'b10000:
        casez_tmp_45 = rob_uop_1_16_ldst_val;
      5'b10001:
        casez_tmp_45 = rob_uop_1_17_ldst_val;
      5'b10010:
        casez_tmp_45 = rob_uop_1_18_ldst_val;
      5'b10011:
        casez_tmp_45 = rob_uop_1_19_ldst_val;
      5'b10100:
        casez_tmp_45 = rob_uop_1_20_ldst_val;
      5'b10101:
        casez_tmp_45 = rob_uop_1_21_ldst_val;
      5'b10110:
        casez_tmp_45 = rob_uop_1_22_ldst_val;
      5'b10111:
        casez_tmp_45 = rob_uop_1_23_ldst_val;
      5'b11000:
        casez_tmp_45 = rob_uop_1_24_ldst_val;
      5'b11001:
        casez_tmp_45 = rob_uop_1_25_ldst_val;
      5'b11010:
        casez_tmp_45 = rob_uop_1_26_ldst_val;
      5'b11011:
        casez_tmp_45 = rob_uop_1_27_ldst_val;
      5'b11100:
        casez_tmp_45 = rob_uop_1_28_ldst_val;
      5'b11101:
        casez_tmp_45 = rob_uop_1_29_ldst_val;
      5'b11110:
        casez_tmp_45 = rob_uop_1_30_ldst_val;
      default:
        casez_tmp_45 = rob_uop_1_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_46 = rob_uop_1_0_dst_rtype;
      5'b00001:
        casez_tmp_46 = rob_uop_1_1_dst_rtype;
      5'b00010:
        casez_tmp_46 = rob_uop_1_2_dst_rtype;
      5'b00011:
        casez_tmp_46 = rob_uop_1_3_dst_rtype;
      5'b00100:
        casez_tmp_46 = rob_uop_1_4_dst_rtype;
      5'b00101:
        casez_tmp_46 = rob_uop_1_5_dst_rtype;
      5'b00110:
        casez_tmp_46 = rob_uop_1_6_dst_rtype;
      5'b00111:
        casez_tmp_46 = rob_uop_1_7_dst_rtype;
      5'b01000:
        casez_tmp_46 = rob_uop_1_8_dst_rtype;
      5'b01001:
        casez_tmp_46 = rob_uop_1_9_dst_rtype;
      5'b01010:
        casez_tmp_46 = rob_uop_1_10_dst_rtype;
      5'b01011:
        casez_tmp_46 = rob_uop_1_11_dst_rtype;
      5'b01100:
        casez_tmp_46 = rob_uop_1_12_dst_rtype;
      5'b01101:
        casez_tmp_46 = rob_uop_1_13_dst_rtype;
      5'b01110:
        casez_tmp_46 = rob_uop_1_14_dst_rtype;
      5'b01111:
        casez_tmp_46 = rob_uop_1_15_dst_rtype;
      5'b10000:
        casez_tmp_46 = rob_uop_1_16_dst_rtype;
      5'b10001:
        casez_tmp_46 = rob_uop_1_17_dst_rtype;
      5'b10010:
        casez_tmp_46 = rob_uop_1_18_dst_rtype;
      5'b10011:
        casez_tmp_46 = rob_uop_1_19_dst_rtype;
      5'b10100:
        casez_tmp_46 = rob_uop_1_20_dst_rtype;
      5'b10101:
        casez_tmp_46 = rob_uop_1_21_dst_rtype;
      5'b10110:
        casez_tmp_46 = rob_uop_1_22_dst_rtype;
      5'b10111:
        casez_tmp_46 = rob_uop_1_23_dst_rtype;
      5'b11000:
        casez_tmp_46 = rob_uop_1_24_dst_rtype;
      5'b11001:
        casez_tmp_46 = rob_uop_1_25_dst_rtype;
      5'b11010:
        casez_tmp_46 = rob_uop_1_26_dst_rtype;
      5'b11011:
        casez_tmp_46 = rob_uop_1_27_dst_rtype;
      5'b11100:
        casez_tmp_46 = rob_uop_1_28_dst_rtype;
      5'b11101:
        casez_tmp_46 = rob_uop_1_29_dst_rtype;
      5'b11110:
        casez_tmp_46 = rob_uop_1_30_dst_rtype;
      default:
        casez_tmp_46 = rob_uop_1_31_dst_rtype;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_47 = rob_uop_1_0_fp_val;
      5'b00001:
        casez_tmp_47 = rob_uop_1_1_fp_val;
      5'b00010:
        casez_tmp_47 = rob_uop_1_2_fp_val;
      5'b00011:
        casez_tmp_47 = rob_uop_1_3_fp_val;
      5'b00100:
        casez_tmp_47 = rob_uop_1_4_fp_val;
      5'b00101:
        casez_tmp_47 = rob_uop_1_5_fp_val;
      5'b00110:
        casez_tmp_47 = rob_uop_1_6_fp_val;
      5'b00111:
        casez_tmp_47 = rob_uop_1_7_fp_val;
      5'b01000:
        casez_tmp_47 = rob_uop_1_8_fp_val;
      5'b01001:
        casez_tmp_47 = rob_uop_1_9_fp_val;
      5'b01010:
        casez_tmp_47 = rob_uop_1_10_fp_val;
      5'b01011:
        casez_tmp_47 = rob_uop_1_11_fp_val;
      5'b01100:
        casez_tmp_47 = rob_uop_1_12_fp_val;
      5'b01101:
        casez_tmp_47 = rob_uop_1_13_fp_val;
      5'b01110:
        casez_tmp_47 = rob_uop_1_14_fp_val;
      5'b01111:
        casez_tmp_47 = rob_uop_1_15_fp_val;
      5'b10000:
        casez_tmp_47 = rob_uop_1_16_fp_val;
      5'b10001:
        casez_tmp_47 = rob_uop_1_17_fp_val;
      5'b10010:
        casez_tmp_47 = rob_uop_1_18_fp_val;
      5'b10011:
        casez_tmp_47 = rob_uop_1_19_fp_val;
      5'b10100:
        casez_tmp_47 = rob_uop_1_20_fp_val;
      5'b10101:
        casez_tmp_47 = rob_uop_1_21_fp_val;
      5'b10110:
        casez_tmp_47 = rob_uop_1_22_fp_val;
      5'b10111:
        casez_tmp_47 = rob_uop_1_23_fp_val;
      5'b11000:
        casez_tmp_47 = rob_uop_1_24_fp_val;
      5'b11001:
        casez_tmp_47 = rob_uop_1_25_fp_val;
      5'b11010:
        casez_tmp_47 = rob_uop_1_26_fp_val;
      5'b11011:
        casez_tmp_47 = rob_uop_1_27_fp_val;
      5'b11100:
        casez_tmp_47 = rob_uop_1_28_fp_val;
      5'b11101:
        casez_tmp_47 = rob_uop_1_29_fp_val;
      5'b11110:
        casez_tmp_47 = rob_uop_1_30_fp_val;
      default:
        casez_tmp_47 = rob_uop_1_31_fp_val;
    endcase
  end // always @(*)
  wire        rbk_row_1 = _io_commit_rollback_T_3 & ~full;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_48 = rob_val_1_0;
      5'b00001:
        casez_tmp_48 = rob_val_1_1;
      5'b00010:
        casez_tmp_48 = rob_val_1_2;
      5'b00011:
        casez_tmp_48 = rob_val_1_3;
      5'b00100:
        casez_tmp_48 = rob_val_1_4;
      5'b00101:
        casez_tmp_48 = rob_val_1_5;
      5'b00110:
        casez_tmp_48 = rob_val_1_6;
      5'b00111:
        casez_tmp_48 = rob_val_1_7;
      5'b01000:
        casez_tmp_48 = rob_val_1_8;
      5'b01001:
        casez_tmp_48 = rob_val_1_9;
      5'b01010:
        casez_tmp_48 = rob_val_1_10;
      5'b01011:
        casez_tmp_48 = rob_val_1_11;
      5'b01100:
        casez_tmp_48 = rob_val_1_12;
      5'b01101:
        casez_tmp_48 = rob_val_1_13;
      5'b01110:
        casez_tmp_48 = rob_val_1_14;
      5'b01111:
        casez_tmp_48 = rob_val_1_15;
      5'b10000:
        casez_tmp_48 = rob_val_1_16;
      5'b10001:
        casez_tmp_48 = rob_val_1_17;
      5'b10010:
        casez_tmp_48 = rob_val_1_18;
      5'b10011:
        casez_tmp_48 = rob_val_1_19;
      5'b10100:
        casez_tmp_48 = rob_val_1_20;
      5'b10101:
        casez_tmp_48 = rob_val_1_21;
      5'b10110:
        casez_tmp_48 = rob_val_1_22;
      5'b10111:
        casez_tmp_48 = rob_val_1_23;
      5'b11000:
        casez_tmp_48 = rob_val_1_24;
      5'b11001:
        casez_tmp_48 = rob_val_1_25;
      5'b11010:
        casez_tmp_48 = rob_val_1_26;
      5'b11011:
        casez_tmp_48 = rob_val_1_27;
      5'b11100:
        casez_tmp_48 = rob_val_1_28;
      5'b11101:
        casez_tmp_48 = rob_val_1_29;
      5'b11110:
        casez_tmp_48 = rob_val_1_30;
      default:
        casez_tmp_48 = rob_val_1_31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_1_output = rbk_row_1 & casez_tmp_48;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_49 = rob_fflags_1_0;
      5'b00001:
        casez_tmp_49 = rob_fflags_1_1;
      5'b00010:
        casez_tmp_49 = rob_fflags_1_2;
      5'b00011:
        casez_tmp_49 = rob_fflags_1_3;
      5'b00100:
        casez_tmp_49 = rob_fflags_1_4;
      5'b00101:
        casez_tmp_49 = rob_fflags_1_5;
      5'b00110:
        casez_tmp_49 = rob_fflags_1_6;
      5'b00111:
        casez_tmp_49 = rob_fflags_1_7;
      5'b01000:
        casez_tmp_49 = rob_fflags_1_8;
      5'b01001:
        casez_tmp_49 = rob_fflags_1_9;
      5'b01010:
        casez_tmp_49 = rob_fflags_1_10;
      5'b01011:
        casez_tmp_49 = rob_fflags_1_11;
      5'b01100:
        casez_tmp_49 = rob_fflags_1_12;
      5'b01101:
        casez_tmp_49 = rob_fflags_1_13;
      5'b01110:
        casez_tmp_49 = rob_fflags_1_14;
      5'b01111:
        casez_tmp_49 = rob_fflags_1_15;
      5'b10000:
        casez_tmp_49 = rob_fflags_1_16;
      5'b10001:
        casez_tmp_49 = rob_fflags_1_17;
      5'b10010:
        casez_tmp_49 = rob_fflags_1_18;
      5'b10011:
        casez_tmp_49 = rob_fflags_1_19;
      5'b10100:
        casez_tmp_49 = rob_fflags_1_20;
      5'b10101:
        casez_tmp_49 = rob_fflags_1_21;
      5'b10110:
        casez_tmp_49 = rob_fflags_1_22;
      5'b10111:
        casez_tmp_49 = rob_fflags_1_23;
      5'b11000:
        casez_tmp_49 = rob_fflags_1_24;
      5'b11001:
        casez_tmp_49 = rob_fflags_1_25;
      5'b11010:
        casez_tmp_49 = rob_fflags_1_26;
      5'b11011:
        casez_tmp_49 = rob_fflags_1_27;
      5'b11100:
        casez_tmp_49 = rob_fflags_1_28;
      5'b11101:
        casez_tmp_49 = rob_fflags_1_29;
      5'b11110:
        casez_tmp_49 = rob_fflags_1_30;
      default:
        casez_tmp_49 = rob_fflags_1_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_50 = rob_uop_1_0_uses_ldq;
      5'b00001:
        casez_tmp_50 = rob_uop_1_1_uses_ldq;
      5'b00010:
        casez_tmp_50 = rob_uop_1_2_uses_ldq;
      5'b00011:
        casez_tmp_50 = rob_uop_1_3_uses_ldq;
      5'b00100:
        casez_tmp_50 = rob_uop_1_4_uses_ldq;
      5'b00101:
        casez_tmp_50 = rob_uop_1_5_uses_ldq;
      5'b00110:
        casez_tmp_50 = rob_uop_1_6_uses_ldq;
      5'b00111:
        casez_tmp_50 = rob_uop_1_7_uses_ldq;
      5'b01000:
        casez_tmp_50 = rob_uop_1_8_uses_ldq;
      5'b01001:
        casez_tmp_50 = rob_uop_1_9_uses_ldq;
      5'b01010:
        casez_tmp_50 = rob_uop_1_10_uses_ldq;
      5'b01011:
        casez_tmp_50 = rob_uop_1_11_uses_ldq;
      5'b01100:
        casez_tmp_50 = rob_uop_1_12_uses_ldq;
      5'b01101:
        casez_tmp_50 = rob_uop_1_13_uses_ldq;
      5'b01110:
        casez_tmp_50 = rob_uop_1_14_uses_ldq;
      5'b01111:
        casez_tmp_50 = rob_uop_1_15_uses_ldq;
      5'b10000:
        casez_tmp_50 = rob_uop_1_16_uses_ldq;
      5'b10001:
        casez_tmp_50 = rob_uop_1_17_uses_ldq;
      5'b10010:
        casez_tmp_50 = rob_uop_1_18_uses_ldq;
      5'b10011:
        casez_tmp_50 = rob_uop_1_19_uses_ldq;
      5'b10100:
        casez_tmp_50 = rob_uop_1_20_uses_ldq;
      5'b10101:
        casez_tmp_50 = rob_uop_1_21_uses_ldq;
      5'b10110:
        casez_tmp_50 = rob_uop_1_22_uses_ldq;
      5'b10111:
        casez_tmp_50 = rob_uop_1_23_uses_ldq;
      5'b11000:
        casez_tmp_50 = rob_uop_1_24_uses_ldq;
      5'b11001:
        casez_tmp_50 = rob_uop_1_25_uses_ldq;
      5'b11010:
        casez_tmp_50 = rob_uop_1_26_uses_ldq;
      5'b11011:
        casez_tmp_50 = rob_uop_1_27_uses_ldq;
      5'b11100:
        casez_tmp_50 = rob_uop_1_28_uses_ldq;
      5'b11101:
        casez_tmp_50 = rob_uop_1_29_uses_ldq;
      5'b11110:
        casez_tmp_50 = rob_uop_1_30_uses_ldq;
      default:
        casez_tmp_50 = rob_uop_1_31_uses_ldq;
    endcase
  end // always @(*)
  reg  [6:0]  rob_uop_2_0_uopc;
  reg         rob_uop_2_0_is_rvc;
  reg  [19:0] rob_uop_2_0_br_mask;
  reg  [5:0]  rob_uop_2_0_ftq_idx;
  reg         rob_uop_2_0_edge_inst;
  reg  [5:0]  rob_uop_2_0_pc_lob;
  reg  [6:0]  rob_uop_2_0_pdst;
  reg  [6:0]  rob_uop_2_0_stale_pdst;
  reg         rob_uop_2_0_is_fencei;
  reg         rob_uop_2_0_uses_ldq;
  reg         rob_uop_2_0_uses_stq;
  reg         rob_uop_2_0_is_sys_pc2epc;
  reg         rob_uop_2_0_flush_on_commit;
  reg  [5:0]  rob_uop_2_0_ldst;
  reg         rob_uop_2_0_ldst_val;
  reg  [1:0]  rob_uop_2_0_dst_rtype;
  reg         rob_uop_2_0_fp_val;
  reg  [6:0]  rob_uop_2_1_uopc;
  reg         rob_uop_2_1_is_rvc;
  reg  [19:0] rob_uop_2_1_br_mask;
  reg  [5:0]  rob_uop_2_1_ftq_idx;
  reg         rob_uop_2_1_edge_inst;
  reg  [5:0]  rob_uop_2_1_pc_lob;
  reg  [6:0]  rob_uop_2_1_pdst;
  reg  [6:0]  rob_uop_2_1_stale_pdst;
  reg         rob_uop_2_1_is_fencei;
  reg         rob_uop_2_1_uses_ldq;
  reg         rob_uop_2_1_uses_stq;
  reg         rob_uop_2_1_is_sys_pc2epc;
  reg         rob_uop_2_1_flush_on_commit;
  reg  [5:0]  rob_uop_2_1_ldst;
  reg         rob_uop_2_1_ldst_val;
  reg  [1:0]  rob_uop_2_1_dst_rtype;
  reg         rob_uop_2_1_fp_val;
  reg  [6:0]  rob_uop_2_2_uopc;
  reg         rob_uop_2_2_is_rvc;
  reg  [19:0] rob_uop_2_2_br_mask;
  reg  [5:0]  rob_uop_2_2_ftq_idx;
  reg         rob_uop_2_2_edge_inst;
  reg  [5:0]  rob_uop_2_2_pc_lob;
  reg  [6:0]  rob_uop_2_2_pdst;
  reg  [6:0]  rob_uop_2_2_stale_pdst;
  reg         rob_uop_2_2_is_fencei;
  reg         rob_uop_2_2_uses_ldq;
  reg         rob_uop_2_2_uses_stq;
  reg         rob_uop_2_2_is_sys_pc2epc;
  reg         rob_uop_2_2_flush_on_commit;
  reg  [5:0]  rob_uop_2_2_ldst;
  reg         rob_uop_2_2_ldst_val;
  reg  [1:0]  rob_uop_2_2_dst_rtype;
  reg         rob_uop_2_2_fp_val;
  reg  [6:0]  rob_uop_2_3_uopc;
  reg         rob_uop_2_3_is_rvc;
  reg  [19:0] rob_uop_2_3_br_mask;
  reg  [5:0]  rob_uop_2_3_ftq_idx;
  reg         rob_uop_2_3_edge_inst;
  reg  [5:0]  rob_uop_2_3_pc_lob;
  reg  [6:0]  rob_uop_2_3_pdst;
  reg  [6:0]  rob_uop_2_3_stale_pdst;
  reg         rob_uop_2_3_is_fencei;
  reg         rob_uop_2_3_uses_ldq;
  reg         rob_uop_2_3_uses_stq;
  reg         rob_uop_2_3_is_sys_pc2epc;
  reg         rob_uop_2_3_flush_on_commit;
  reg  [5:0]  rob_uop_2_3_ldst;
  reg         rob_uop_2_3_ldst_val;
  reg  [1:0]  rob_uop_2_3_dst_rtype;
  reg         rob_uop_2_3_fp_val;
  reg  [6:0]  rob_uop_2_4_uopc;
  reg         rob_uop_2_4_is_rvc;
  reg  [19:0] rob_uop_2_4_br_mask;
  reg  [5:0]  rob_uop_2_4_ftq_idx;
  reg         rob_uop_2_4_edge_inst;
  reg  [5:0]  rob_uop_2_4_pc_lob;
  reg  [6:0]  rob_uop_2_4_pdst;
  reg  [6:0]  rob_uop_2_4_stale_pdst;
  reg         rob_uop_2_4_is_fencei;
  reg         rob_uop_2_4_uses_ldq;
  reg         rob_uop_2_4_uses_stq;
  reg         rob_uop_2_4_is_sys_pc2epc;
  reg         rob_uop_2_4_flush_on_commit;
  reg  [5:0]  rob_uop_2_4_ldst;
  reg         rob_uop_2_4_ldst_val;
  reg  [1:0]  rob_uop_2_4_dst_rtype;
  reg         rob_uop_2_4_fp_val;
  reg  [6:0]  rob_uop_2_5_uopc;
  reg         rob_uop_2_5_is_rvc;
  reg  [19:0] rob_uop_2_5_br_mask;
  reg  [5:0]  rob_uop_2_5_ftq_idx;
  reg         rob_uop_2_5_edge_inst;
  reg  [5:0]  rob_uop_2_5_pc_lob;
  reg  [6:0]  rob_uop_2_5_pdst;
  reg  [6:0]  rob_uop_2_5_stale_pdst;
  reg         rob_uop_2_5_is_fencei;
  reg         rob_uop_2_5_uses_ldq;
  reg         rob_uop_2_5_uses_stq;
  reg         rob_uop_2_5_is_sys_pc2epc;
  reg         rob_uop_2_5_flush_on_commit;
  reg  [5:0]  rob_uop_2_5_ldst;
  reg         rob_uop_2_5_ldst_val;
  reg  [1:0]  rob_uop_2_5_dst_rtype;
  reg         rob_uop_2_5_fp_val;
  reg  [6:0]  rob_uop_2_6_uopc;
  reg         rob_uop_2_6_is_rvc;
  reg  [19:0] rob_uop_2_6_br_mask;
  reg  [5:0]  rob_uop_2_6_ftq_idx;
  reg         rob_uop_2_6_edge_inst;
  reg  [5:0]  rob_uop_2_6_pc_lob;
  reg  [6:0]  rob_uop_2_6_pdst;
  reg  [6:0]  rob_uop_2_6_stale_pdst;
  reg         rob_uop_2_6_is_fencei;
  reg         rob_uop_2_6_uses_ldq;
  reg         rob_uop_2_6_uses_stq;
  reg         rob_uop_2_6_is_sys_pc2epc;
  reg         rob_uop_2_6_flush_on_commit;
  reg  [5:0]  rob_uop_2_6_ldst;
  reg         rob_uop_2_6_ldst_val;
  reg  [1:0]  rob_uop_2_6_dst_rtype;
  reg         rob_uop_2_6_fp_val;
  reg  [6:0]  rob_uop_2_7_uopc;
  reg         rob_uop_2_7_is_rvc;
  reg  [19:0] rob_uop_2_7_br_mask;
  reg  [5:0]  rob_uop_2_7_ftq_idx;
  reg         rob_uop_2_7_edge_inst;
  reg  [5:0]  rob_uop_2_7_pc_lob;
  reg  [6:0]  rob_uop_2_7_pdst;
  reg  [6:0]  rob_uop_2_7_stale_pdst;
  reg         rob_uop_2_7_is_fencei;
  reg         rob_uop_2_7_uses_ldq;
  reg         rob_uop_2_7_uses_stq;
  reg         rob_uop_2_7_is_sys_pc2epc;
  reg         rob_uop_2_7_flush_on_commit;
  reg  [5:0]  rob_uop_2_7_ldst;
  reg         rob_uop_2_7_ldst_val;
  reg  [1:0]  rob_uop_2_7_dst_rtype;
  reg         rob_uop_2_7_fp_val;
  reg  [6:0]  rob_uop_2_8_uopc;
  reg         rob_uop_2_8_is_rvc;
  reg  [19:0] rob_uop_2_8_br_mask;
  reg  [5:0]  rob_uop_2_8_ftq_idx;
  reg         rob_uop_2_8_edge_inst;
  reg  [5:0]  rob_uop_2_8_pc_lob;
  reg  [6:0]  rob_uop_2_8_pdst;
  reg  [6:0]  rob_uop_2_8_stale_pdst;
  reg         rob_uop_2_8_is_fencei;
  reg         rob_uop_2_8_uses_ldq;
  reg         rob_uop_2_8_uses_stq;
  reg         rob_uop_2_8_is_sys_pc2epc;
  reg         rob_uop_2_8_flush_on_commit;
  reg  [5:0]  rob_uop_2_8_ldst;
  reg         rob_uop_2_8_ldst_val;
  reg  [1:0]  rob_uop_2_8_dst_rtype;
  reg         rob_uop_2_8_fp_val;
  reg  [6:0]  rob_uop_2_9_uopc;
  reg         rob_uop_2_9_is_rvc;
  reg  [19:0] rob_uop_2_9_br_mask;
  reg  [5:0]  rob_uop_2_9_ftq_idx;
  reg         rob_uop_2_9_edge_inst;
  reg  [5:0]  rob_uop_2_9_pc_lob;
  reg  [6:0]  rob_uop_2_9_pdst;
  reg  [6:0]  rob_uop_2_9_stale_pdst;
  reg         rob_uop_2_9_is_fencei;
  reg         rob_uop_2_9_uses_ldq;
  reg         rob_uop_2_9_uses_stq;
  reg         rob_uop_2_9_is_sys_pc2epc;
  reg         rob_uop_2_9_flush_on_commit;
  reg  [5:0]  rob_uop_2_9_ldst;
  reg         rob_uop_2_9_ldst_val;
  reg  [1:0]  rob_uop_2_9_dst_rtype;
  reg         rob_uop_2_9_fp_val;
  reg  [6:0]  rob_uop_2_10_uopc;
  reg         rob_uop_2_10_is_rvc;
  reg  [19:0] rob_uop_2_10_br_mask;
  reg  [5:0]  rob_uop_2_10_ftq_idx;
  reg         rob_uop_2_10_edge_inst;
  reg  [5:0]  rob_uop_2_10_pc_lob;
  reg  [6:0]  rob_uop_2_10_pdst;
  reg  [6:0]  rob_uop_2_10_stale_pdst;
  reg         rob_uop_2_10_is_fencei;
  reg         rob_uop_2_10_uses_ldq;
  reg         rob_uop_2_10_uses_stq;
  reg         rob_uop_2_10_is_sys_pc2epc;
  reg         rob_uop_2_10_flush_on_commit;
  reg  [5:0]  rob_uop_2_10_ldst;
  reg         rob_uop_2_10_ldst_val;
  reg  [1:0]  rob_uop_2_10_dst_rtype;
  reg         rob_uop_2_10_fp_val;
  reg  [6:0]  rob_uop_2_11_uopc;
  reg         rob_uop_2_11_is_rvc;
  reg  [19:0] rob_uop_2_11_br_mask;
  reg  [5:0]  rob_uop_2_11_ftq_idx;
  reg         rob_uop_2_11_edge_inst;
  reg  [5:0]  rob_uop_2_11_pc_lob;
  reg  [6:0]  rob_uop_2_11_pdst;
  reg  [6:0]  rob_uop_2_11_stale_pdst;
  reg         rob_uop_2_11_is_fencei;
  reg         rob_uop_2_11_uses_ldq;
  reg         rob_uop_2_11_uses_stq;
  reg         rob_uop_2_11_is_sys_pc2epc;
  reg         rob_uop_2_11_flush_on_commit;
  reg  [5:0]  rob_uop_2_11_ldst;
  reg         rob_uop_2_11_ldst_val;
  reg  [1:0]  rob_uop_2_11_dst_rtype;
  reg         rob_uop_2_11_fp_val;
  reg  [6:0]  rob_uop_2_12_uopc;
  reg         rob_uop_2_12_is_rvc;
  reg  [19:0] rob_uop_2_12_br_mask;
  reg  [5:0]  rob_uop_2_12_ftq_idx;
  reg         rob_uop_2_12_edge_inst;
  reg  [5:0]  rob_uop_2_12_pc_lob;
  reg  [6:0]  rob_uop_2_12_pdst;
  reg  [6:0]  rob_uop_2_12_stale_pdst;
  reg         rob_uop_2_12_is_fencei;
  reg         rob_uop_2_12_uses_ldq;
  reg         rob_uop_2_12_uses_stq;
  reg         rob_uop_2_12_is_sys_pc2epc;
  reg         rob_uop_2_12_flush_on_commit;
  reg  [5:0]  rob_uop_2_12_ldst;
  reg         rob_uop_2_12_ldst_val;
  reg  [1:0]  rob_uop_2_12_dst_rtype;
  reg         rob_uop_2_12_fp_val;
  reg  [6:0]  rob_uop_2_13_uopc;
  reg         rob_uop_2_13_is_rvc;
  reg  [19:0] rob_uop_2_13_br_mask;
  reg  [5:0]  rob_uop_2_13_ftq_idx;
  reg         rob_uop_2_13_edge_inst;
  reg  [5:0]  rob_uop_2_13_pc_lob;
  reg  [6:0]  rob_uop_2_13_pdst;
  reg  [6:0]  rob_uop_2_13_stale_pdst;
  reg         rob_uop_2_13_is_fencei;
  reg         rob_uop_2_13_uses_ldq;
  reg         rob_uop_2_13_uses_stq;
  reg         rob_uop_2_13_is_sys_pc2epc;
  reg         rob_uop_2_13_flush_on_commit;
  reg  [5:0]  rob_uop_2_13_ldst;
  reg         rob_uop_2_13_ldst_val;
  reg  [1:0]  rob_uop_2_13_dst_rtype;
  reg         rob_uop_2_13_fp_val;
  reg  [6:0]  rob_uop_2_14_uopc;
  reg         rob_uop_2_14_is_rvc;
  reg  [19:0] rob_uop_2_14_br_mask;
  reg  [5:0]  rob_uop_2_14_ftq_idx;
  reg         rob_uop_2_14_edge_inst;
  reg  [5:0]  rob_uop_2_14_pc_lob;
  reg  [6:0]  rob_uop_2_14_pdst;
  reg  [6:0]  rob_uop_2_14_stale_pdst;
  reg         rob_uop_2_14_is_fencei;
  reg         rob_uop_2_14_uses_ldq;
  reg         rob_uop_2_14_uses_stq;
  reg         rob_uop_2_14_is_sys_pc2epc;
  reg         rob_uop_2_14_flush_on_commit;
  reg  [5:0]  rob_uop_2_14_ldst;
  reg         rob_uop_2_14_ldst_val;
  reg  [1:0]  rob_uop_2_14_dst_rtype;
  reg         rob_uop_2_14_fp_val;
  reg  [6:0]  rob_uop_2_15_uopc;
  reg         rob_uop_2_15_is_rvc;
  reg  [19:0] rob_uop_2_15_br_mask;
  reg  [5:0]  rob_uop_2_15_ftq_idx;
  reg         rob_uop_2_15_edge_inst;
  reg  [5:0]  rob_uop_2_15_pc_lob;
  reg  [6:0]  rob_uop_2_15_pdst;
  reg  [6:0]  rob_uop_2_15_stale_pdst;
  reg         rob_uop_2_15_is_fencei;
  reg         rob_uop_2_15_uses_ldq;
  reg         rob_uop_2_15_uses_stq;
  reg         rob_uop_2_15_is_sys_pc2epc;
  reg         rob_uop_2_15_flush_on_commit;
  reg  [5:0]  rob_uop_2_15_ldst;
  reg         rob_uop_2_15_ldst_val;
  reg  [1:0]  rob_uop_2_15_dst_rtype;
  reg         rob_uop_2_15_fp_val;
  reg  [6:0]  rob_uop_2_16_uopc;
  reg         rob_uop_2_16_is_rvc;
  reg  [19:0] rob_uop_2_16_br_mask;
  reg  [5:0]  rob_uop_2_16_ftq_idx;
  reg         rob_uop_2_16_edge_inst;
  reg  [5:0]  rob_uop_2_16_pc_lob;
  reg  [6:0]  rob_uop_2_16_pdst;
  reg  [6:0]  rob_uop_2_16_stale_pdst;
  reg         rob_uop_2_16_is_fencei;
  reg         rob_uop_2_16_uses_ldq;
  reg         rob_uop_2_16_uses_stq;
  reg         rob_uop_2_16_is_sys_pc2epc;
  reg         rob_uop_2_16_flush_on_commit;
  reg  [5:0]  rob_uop_2_16_ldst;
  reg         rob_uop_2_16_ldst_val;
  reg  [1:0]  rob_uop_2_16_dst_rtype;
  reg         rob_uop_2_16_fp_val;
  reg  [6:0]  rob_uop_2_17_uopc;
  reg         rob_uop_2_17_is_rvc;
  reg  [19:0] rob_uop_2_17_br_mask;
  reg  [5:0]  rob_uop_2_17_ftq_idx;
  reg         rob_uop_2_17_edge_inst;
  reg  [5:0]  rob_uop_2_17_pc_lob;
  reg  [6:0]  rob_uop_2_17_pdst;
  reg  [6:0]  rob_uop_2_17_stale_pdst;
  reg         rob_uop_2_17_is_fencei;
  reg         rob_uop_2_17_uses_ldq;
  reg         rob_uop_2_17_uses_stq;
  reg         rob_uop_2_17_is_sys_pc2epc;
  reg         rob_uop_2_17_flush_on_commit;
  reg  [5:0]  rob_uop_2_17_ldst;
  reg         rob_uop_2_17_ldst_val;
  reg  [1:0]  rob_uop_2_17_dst_rtype;
  reg         rob_uop_2_17_fp_val;
  reg  [6:0]  rob_uop_2_18_uopc;
  reg         rob_uop_2_18_is_rvc;
  reg  [19:0] rob_uop_2_18_br_mask;
  reg  [5:0]  rob_uop_2_18_ftq_idx;
  reg         rob_uop_2_18_edge_inst;
  reg  [5:0]  rob_uop_2_18_pc_lob;
  reg  [6:0]  rob_uop_2_18_pdst;
  reg  [6:0]  rob_uop_2_18_stale_pdst;
  reg         rob_uop_2_18_is_fencei;
  reg         rob_uop_2_18_uses_ldq;
  reg         rob_uop_2_18_uses_stq;
  reg         rob_uop_2_18_is_sys_pc2epc;
  reg         rob_uop_2_18_flush_on_commit;
  reg  [5:0]  rob_uop_2_18_ldst;
  reg         rob_uop_2_18_ldst_val;
  reg  [1:0]  rob_uop_2_18_dst_rtype;
  reg         rob_uop_2_18_fp_val;
  reg  [6:0]  rob_uop_2_19_uopc;
  reg         rob_uop_2_19_is_rvc;
  reg  [19:0] rob_uop_2_19_br_mask;
  reg  [5:0]  rob_uop_2_19_ftq_idx;
  reg         rob_uop_2_19_edge_inst;
  reg  [5:0]  rob_uop_2_19_pc_lob;
  reg  [6:0]  rob_uop_2_19_pdst;
  reg  [6:0]  rob_uop_2_19_stale_pdst;
  reg         rob_uop_2_19_is_fencei;
  reg         rob_uop_2_19_uses_ldq;
  reg         rob_uop_2_19_uses_stq;
  reg         rob_uop_2_19_is_sys_pc2epc;
  reg         rob_uop_2_19_flush_on_commit;
  reg  [5:0]  rob_uop_2_19_ldst;
  reg         rob_uop_2_19_ldst_val;
  reg  [1:0]  rob_uop_2_19_dst_rtype;
  reg         rob_uop_2_19_fp_val;
  reg  [6:0]  rob_uop_2_20_uopc;
  reg         rob_uop_2_20_is_rvc;
  reg  [19:0] rob_uop_2_20_br_mask;
  reg  [5:0]  rob_uop_2_20_ftq_idx;
  reg         rob_uop_2_20_edge_inst;
  reg  [5:0]  rob_uop_2_20_pc_lob;
  reg  [6:0]  rob_uop_2_20_pdst;
  reg  [6:0]  rob_uop_2_20_stale_pdst;
  reg         rob_uop_2_20_is_fencei;
  reg         rob_uop_2_20_uses_ldq;
  reg         rob_uop_2_20_uses_stq;
  reg         rob_uop_2_20_is_sys_pc2epc;
  reg         rob_uop_2_20_flush_on_commit;
  reg  [5:0]  rob_uop_2_20_ldst;
  reg         rob_uop_2_20_ldst_val;
  reg  [1:0]  rob_uop_2_20_dst_rtype;
  reg         rob_uop_2_20_fp_val;
  reg  [6:0]  rob_uop_2_21_uopc;
  reg         rob_uop_2_21_is_rvc;
  reg  [19:0] rob_uop_2_21_br_mask;
  reg  [5:0]  rob_uop_2_21_ftq_idx;
  reg         rob_uop_2_21_edge_inst;
  reg  [5:0]  rob_uop_2_21_pc_lob;
  reg  [6:0]  rob_uop_2_21_pdst;
  reg  [6:0]  rob_uop_2_21_stale_pdst;
  reg         rob_uop_2_21_is_fencei;
  reg         rob_uop_2_21_uses_ldq;
  reg         rob_uop_2_21_uses_stq;
  reg         rob_uop_2_21_is_sys_pc2epc;
  reg         rob_uop_2_21_flush_on_commit;
  reg  [5:0]  rob_uop_2_21_ldst;
  reg         rob_uop_2_21_ldst_val;
  reg  [1:0]  rob_uop_2_21_dst_rtype;
  reg         rob_uop_2_21_fp_val;
  reg  [6:0]  rob_uop_2_22_uopc;
  reg         rob_uop_2_22_is_rvc;
  reg  [19:0] rob_uop_2_22_br_mask;
  reg  [5:0]  rob_uop_2_22_ftq_idx;
  reg         rob_uop_2_22_edge_inst;
  reg  [5:0]  rob_uop_2_22_pc_lob;
  reg  [6:0]  rob_uop_2_22_pdst;
  reg  [6:0]  rob_uop_2_22_stale_pdst;
  reg         rob_uop_2_22_is_fencei;
  reg         rob_uop_2_22_uses_ldq;
  reg         rob_uop_2_22_uses_stq;
  reg         rob_uop_2_22_is_sys_pc2epc;
  reg         rob_uop_2_22_flush_on_commit;
  reg  [5:0]  rob_uop_2_22_ldst;
  reg         rob_uop_2_22_ldst_val;
  reg  [1:0]  rob_uop_2_22_dst_rtype;
  reg         rob_uop_2_22_fp_val;
  reg  [6:0]  rob_uop_2_23_uopc;
  reg         rob_uop_2_23_is_rvc;
  reg  [19:0] rob_uop_2_23_br_mask;
  reg  [5:0]  rob_uop_2_23_ftq_idx;
  reg         rob_uop_2_23_edge_inst;
  reg  [5:0]  rob_uop_2_23_pc_lob;
  reg  [6:0]  rob_uop_2_23_pdst;
  reg  [6:0]  rob_uop_2_23_stale_pdst;
  reg         rob_uop_2_23_is_fencei;
  reg         rob_uop_2_23_uses_ldq;
  reg         rob_uop_2_23_uses_stq;
  reg         rob_uop_2_23_is_sys_pc2epc;
  reg         rob_uop_2_23_flush_on_commit;
  reg  [5:0]  rob_uop_2_23_ldst;
  reg         rob_uop_2_23_ldst_val;
  reg  [1:0]  rob_uop_2_23_dst_rtype;
  reg         rob_uop_2_23_fp_val;
  reg  [6:0]  rob_uop_2_24_uopc;
  reg         rob_uop_2_24_is_rvc;
  reg  [19:0] rob_uop_2_24_br_mask;
  reg  [5:0]  rob_uop_2_24_ftq_idx;
  reg         rob_uop_2_24_edge_inst;
  reg  [5:0]  rob_uop_2_24_pc_lob;
  reg  [6:0]  rob_uop_2_24_pdst;
  reg  [6:0]  rob_uop_2_24_stale_pdst;
  reg         rob_uop_2_24_is_fencei;
  reg         rob_uop_2_24_uses_ldq;
  reg         rob_uop_2_24_uses_stq;
  reg         rob_uop_2_24_is_sys_pc2epc;
  reg         rob_uop_2_24_flush_on_commit;
  reg  [5:0]  rob_uop_2_24_ldst;
  reg         rob_uop_2_24_ldst_val;
  reg  [1:0]  rob_uop_2_24_dst_rtype;
  reg         rob_uop_2_24_fp_val;
  reg  [6:0]  rob_uop_2_25_uopc;
  reg         rob_uop_2_25_is_rvc;
  reg  [19:0] rob_uop_2_25_br_mask;
  reg  [5:0]  rob_uop_2_25_ftq_idx;
  reg         rob_uop_2_25_edge_inst;
  reg  [5:0]  rob_uop_2_25_pc_lob;
  reg  [6:0]  rob_uop_2_25_pdst;
  reg  [6:0]  rob_uop_2_25_stale_pdst;
  reg         rob_uop_2_25_is_fencei;
  reg         rob_uop_2_25_uses_ldq;
  reg         rob_uop_2_25_uses_stq;
  reg         rob_uop_2_25_is_sys_pc2epc;
  reg         rob_uop_2_25_flush_on_commit;
  reg  [5:0]  rob_uop_2_25_ldst;
  reg         rob_uop_2_25_ldst_val;
  reg  [1:0]  rob_uop_2_25_dst_rtype;
  reg         rob_uop_2_25_fp_val;
  reg  [6:0]  rob_uop_2_26_uopc;
  reg         rob_uop_2_26_is_rvc;
  reg  [19:0] rob_uop_2_26_br_mask;
  reg  [5:0]  rob_uop_2_26_ftq_idx;
  reg         rob_uop_2_26_edge_inst;
  reg  [5:0]  rob_uop_2_26_pc_lob;
  reg  [6:0]  rob_uop_2_26_pdst;
  reg  [6:0]  rob_uop_2_26_stale_pdst;
  reg         rob_uop_2_26_is_fencei;
  reg         rob_uop_2_26_uses_ldq;
  reg         rob_uop_2_26_uses_stq;
  reg         rob_uop_2_26_is_sys_pc2epc;
  reg         rob_uop_2_26_flush_on_commit;
  reg  [5:0]  rob_uop_2_26_ldst;
  reg         rob_uop_2_26_ldst_val;
  reg  [1:0]  rob_uop_2_26_dst_rtype;
  reg         rob_uop_2_26_fp_val;
  reg  [6:0]  rob_uop_2_27_uopc;
  reg         rob_uop_2_27_is_rvc;
  reg  [19:0] rob_uop_2_27_br_mask;
  reg  [5:0]  rob_uop_2_27_ftq_idx;
  reg         rob_uop_2_27_edge_inst;
  reg  [5:0]  rob_uop_2_27_pc_lob;
  reg  [6:0]  rob_uop_2_27_pdst;
  reg  [6:0]  rob_uop_2_27_stale_pdst;
  reg         rob_uop_2_27_is_fencei;
  reg         rob_uop_2_27_uses_ldq;
  reg         rob_uop_2_27_uses_stq;
  reg         rob_uop_2_27_is_sys_pc2epc;
  reg         rob_uop_2_27_flush_on_commit;
  reg  [5:0]  rob_uop_2_27_ldst;
  reg         rob_uop_2_27_ldst_val;
  reg  [1:0]  rob_uop_2_27_dst_rtype;
  reg         rob_uop_2_27_fp_val;
  reg  [6:0]  rob_uop_2_28_uopc;
  reg         rob_uop_2_28_is_rvc;
  reg  [19:0] rob_uop_2_28_br_mask;
  reg  [5:0]  rob_uop_2_28_ftq_idx;
  reg         rob_uop_2_28_edge_inst;
  reg  [5:0]  rob_uop_2_28_pc_lob;
  reg  [6:0]  rob_uop_2_28_pdst;
  reg  [6:0]  rob_uop_2_28_stale_pdst;
  reg         rob_uop_2_28_is_fencei;
  reg         rob_uop_2_28_uses_ldq;
  reg         rob_uop_2_28_uses_stq;
  reg         rob_uop_2_28_is_sys_pc2epc;
  reg         rob_uop_2_28_flush_on_commit;
  reg  [5:0]  rob_uop_2_28_ldst;
  reg         rob_uop_2_28_ldst_val;
  reg  [1:0]  rob_uop_2_28_dst_rtype;
  reg         rob_uop_2_28_fp_val;
  reg  [6:0]  rob_uop_2_29_uopc;
  reg         rob_uop_2_29_is_rvc;
  reg  [19:0] rob_uop_2_29_br_mask;
  reg  [5:0]  rob_uop_2_29_ftq_idx;
  reg         rob_uop_2_29_edge_inst;
  reg  [5:0]  rob_uop_2_29_pc_lob;
  reg  [6:0]  rob_uop_2_29_pdst;
  reg  [6:0]  rob_uop_2_29_stale_pdst;
  reg         rob_uop_2_29_is_fencei;
  reg         rob_uop_2_29_uses_ldq;
  reg         rob_uop_2_29_uses_stq;
  reg         rob_uop_2_29_is_sys_pc2epc;
  reg         rob_uop_2_29_flush_on_commit;
  reg  [5:0]  rob_uop_2_29_ldst;
  reg         rob_uop_2_29_ldst_val;
  reg  [1:0]  rob_uop_2_29_dst_rtype;
  reg         rob_uop_2_29_fp_val;
  reg  [6:0]  rob_uop_2_30_uopc;
  reg         rob_uop_2_30_is_rvc;
  reg  [19:0] rob_uop_2_30_br_mask;
  reg  [5:0]  rob_uop_2_30_ftq_idx;
  reg         rob_uop_2_30_edge_inst;
  reg  [5:0]  rob_uop_2_30_pc_lob;
  reg  [6:0]  rob_uop_2_30_pdst;
  reg  [6:0]  rob_uop_2_30_stale_pdst;
  reg         rob_uop_2_30_is_fencei;
  reg         rob_uop_2_30_uses_ldq;
  reg         rob_uop_2_30_uses_stq;
  reg         rob_uop_2_30_is_sys_pc2epc;
  reg         rob_uop_2_30_flush_on_commit;
  reg  [5:0]  rob_uop_2_30_ldst;
  reg         rob_uop_2_30_ldst_val;
  reg  [1:0]  rob_uop_2_30_dst_rtype;
  reg         rob_uop_2_30_fp_val;
  reg  [6:0]  rob_uop_2_31_uopc;
  reg         rob_uop_2_31_is_rvc;
  reg  [19:0] rob_uop_2_31_br_mask;
  reg  [5:0]  rob_uop_2_31_ftq_idx;
  reg         rob_uop_2_31_edge_inst;
  reg  [5:0]  rob_uop_2_31_pc_lob;
  reg  [6:0]  rob_uop_2_31_pdst;
  reg  [6:0]  rob_uop_2_31_stale_pdst;
  reg         rob_uop_2_31_is_fencei;
  reg         rob_uop_2_31_uses_ldq;
  reg         rob_uop_2_31_uses_stq;
  reg         rob_uop_2_31_is_sys_pc2epc;
  reg         rob_uop_2_31_flush_on_commit;
  reg  [5:0]  rob_uop_2_31_ldst;
  reg         rob_uop_2_31_ldst_val;
  reg  [1:0]  rob_uop_2_31_dst_rtype;
  reg         rob_uop_2_31_fp_val;
  reg         rob_predicated_2_0;
  reg         rob_predicated_2_1;
  reg         rob_predicated_2_2;
  reg         rob_predicated_2_3;
  reg         rob_predicated_2_4;
  reg         rob_predicated_2_5;
  reg         rob_predicated_2_6;
  reg         rob_predicated_2_7;
  reg         rob_predicated_2_8;
  reg         rob_predicated_2_9;
  reg         rob_predicated_2_10;
  reg         rob_predicated_2_11;
  reg         rob_predicated_2_12;
  reg         rob_predicated_2_13;
  reg         rob_predicated_2_14;
  reg         rob_predicated_2_15;
  reg         rob_predicated_2_16;
  reg         rob_predicated_2_17;
  reg         rob_predicated_2_18;
  reg         rob_predicated_2_19;
  reg         rob_predicated_2_20;
  reg         rob_predicated_2_21;
  reg         rob_predicated_2_22;
  reg         rob_predicated_2_23;
  reg         rob_predicated_2_24;
  reg         rob_predicated_2_25;
  reg         rob_predicated_2_26;
  reg         rob_predicated_2_27;
  reg         rob_predicated_2_28;
  reg         rob_predicated_2_29;
  reg         rob_predicated_2_30;
  reg         rob_predicated_2_31;
  wire        _GEN_1360 = io_enq_valids_2 & _GEN_2;
  wire        _GEN_1361 = io_enq_valids_2 & _GEN_3;
  wire        _GEN_1362 = io_enq_valids_2 & _GEN_4;
  wire        _GEN_1363 = io_enq_valids_2 & _GEN_5;
  wire        _GEN_1364 = io_enq_valids_2 & _GEN_6;
  wire        _GEN_1365 = io_enq_valids_2 & _GEN_7;
  wire        _GEN_1366 = io_enq_valids_2 & _GEN_8;
  wire        _GEN_1367 = io_enq_valids_2 & _GEN_9;
  wire        _GEN_1368 = io_enq_valids_2 & _GEN_10;
  wire        _GEN_1369 = io_enq_valids_2 & _GEN_11;
  wire        _GEN_1370 = io_enq_valids_2 & _GEN_12;
  wire        _GEN_1371 = io_enq_valids_2 & _GEN_13;
  wire        _GEN_1372 = io_enq_valids_2 & _GEN_14;
  wire        _GEN_1373 = io_enq_valids_2 & _GEN_15;
  wire        _GEN_1374 = io_enq_valids_2 & _GEN_16;
  wire        _GEN_1375 = io_enq_valids_2 & _GEN_17;
  wire        _GEN_1376 = io_enq_valids_2 & _GEN_18;
  wire        _GEN_1377 = io_enq_valids_2 & _GEN_19;
  wire        _GEN_1378 = io_enq_valids_2 & _GEN_20;
  wire        _GEN_1379 = io_enq_valids_2 & _GEN_21;
  wire        _GEN_1380 = io_enq_valids_2 & _GEN_22;
  wire        _GEN_1381 = io_enq_valids_2 & _GEN_23;
  wire        _GEN_1382 = io_enq_valids_2 & _GEN_24;
  wire        _GEN_1383 = io_enq_valids_2 & _GEN_25;
  wire        _GEN_1384 = io_enq_valids_2 & _GEN_26;
  wire        _GEN_1385 = io_enq_valids_2 & _GEN_27;
  wire        _GEN_1386 = io_enq_valids_2 & _GEN_28;
  wire        _GEN_1387 = io_enq_valids_2 & _GEN_29;
  wire        _GEN_1388 = io_enq_valids_2 & _GEN_30;
  wire        _GEN_1389 = io_enq_valids_2 & _GEN_31;
  wire        _GEN_1390 = io_enq_valids_2 & _GEN_32;
  wire        _GEN_1391 = io_enq_valids_2 & (&rob_tail);
  wire        _GEN_1392 = io_wb_resps_0_valid & io_wb_resps_0_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1393 = _GEN_1392 & _GEN_66;
  wire        _GEN_1394 = _GEN_1392 & _GEN_67;
  wire        _GEN_1395 = _GEN_1392 & _GEN_68;
  wire        _GEN_1396 = _GEN_1392 & _GEN_69;
  wire        _GEN_1397 = _GEN_1392 & _GEN_70;
  wire        _GEN_1398 = _GEN_1392 & _GEN_71;
  wire        _GEN_1399 = _GEN_1392 & _GEN_72;
  wire        _GEN_1400 = _GEN_1392 & _GEN_73;
  wire        _GEN_1401 = _GEN_1392 & _GEN_74;
  wire        _GEN_1402 = _GEN_1392 & _GEN_75;
  wire        _GEN_1403 = _GEN_1392 & _GEN_76;
  wire        _GEN_1404 = _GEN_1392 & _GEN_77;
  wire        _GEN_1405 = _GEN_1392 & _GEN_78;
  wire        _GEN_1406 = _GEN_1392 & _GEN_79;
  wire        _GEN_1407 = _GEN_1392 & _GEN_80;
  wire        _GEN_1408 = _GEN_1392 & _GEN_81;
  wire        _GEN_1409 = _GEN_1392 & _GEN_82;
  wire        _GEN_1410 = _GEN_1392 & _GEN_83;
  wire        _GEN_1411 = _GEN_1392 & _GEN_84;
  wire        _GEN_1412 = _GEN_1392 & _GEN_85;
  wire        _GEN_1413 = _GEN_1392 & _GEN_86;
  wire        _GEN_1414 = _GEN_1392 & _GEN_87;
  wire        _GEN_1415 = _GEN_1392 & _GEN_88;
  wire        _GEN_1416 = _GEN_1392 & _GEN_89;
  wire        _GEN_1417 = _GEN_1392 & _GEN_90;
  wire        _GEN_1418 = _GEN_1392 & _GEN_91;
  wire        _GEN_1419 = _GEN_1392 & _GEN_92;
  wire        _GEN_1420 = _GEN_1392 & _GEN_93;
  wire        _GEN_1421 = _GEN_1392 & _GEN_94;
  wire        _GEN_1422 = _GEN_1392 & _GEN_95;
  wire        _GEN_1423 = _GEN_1392 & _GEN_96;
  wire        _GEN_1424 = _GEN_1392 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_1425 = io_wb_resps_1_valid & io_wb_resps_1_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1426 = _GEN_130 | _GEN_1393;
  wire        _GEN_1427 = _GEN_132 | _GEN_1394;
  wire        _GEN_1428 = _GEN_134 | _GEN_1395;
  wire        _GEN_1429 = _GEN_136 | _GEN_1396;
  wire        _GEN_1430 = _GEN_138 | _GEN_1397;
  wire        _GEN_1431 = _GEN_140 | _GEN_1398;
  wire        _GEN_1432 = _GEN_142 | _GEN_1399;
  wire        _GEN_1433 = _GEN_144 | _GEN_1400;
  wire        _GEN_1434 = _GEN_146 | _GEN_1401;
  wire        _GEN_1435 = _GEN_148 | _GEN_1402;
  wire        _GEN_1436 = _GEN_150 | _GEN_1403;
  wire        _GEN_1437 = _GEN_152 | _GEN_1404;
  wire        _GEN_1438 = _GEN_154 | _GEN_1405;
  wire        _GEN_1439 = _GEN_156 | _GEN_1406;
  wire        _GEN_1440 = _GEN_158 | _GEN_1407;
  wire        _GEN_1441 = _GEN_160 | _GEN_1408;
  wire        _GEN_1442 = _GEN_162 | _GEN_1409;
  wire        _GEN_1443 = _GEN_164 | _GEN_1410;
  wire        _GEN_1444 = _GEN_166 | _GEN_1411;
  wire        _GEN_1445 = _GEN_168 | _GEN_1412;
  wire        _GEN_1446 = _GEN_170 | _GEN_1413;
  wire        _GEN_1447 = _GEN_172 | _GEN_1414;
  wire        _GEN_1448 = _GEN_174 | _GEN_1415;
  wire        _GEN_1449 = _GEN_176 | _GEN_1416;
  wire        _GEN_1450 = _GEN_178 | _GEN_1417;
  wire        _GEN_1451 = _GEN_180 | _GEN_1418;
  wire        _GEN_1452 = _GEN_182 | _GEN_1419;
  wire        _GEN_1453 = _GEN_184 | _GEN_1420;
  wire        _GEN_1454 = _GEN_186 | _GEN_1421;
  wire        _GEN_1455 = _GEN_188 | _GEN_1422;
  wire        _GEN_1456 = _GEN_190 | _GEN_1423;
  wire        _GEN_1457 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_1424;
  wire        _GEN_1458 = io_wb_resps_2_valid & io_wb_resps_2_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1459 = _GEN_1458 & _GEN_194;
  wire        _GEN_1460 = _GEN_1458 & _GEN_195;
  wire        _GEN_1461 = _GEN_1458 & _GEN_196;
  wire        _GEN_1462 = _GEN_1458 & _GEN_197;
  wire        _GEN_1463 = _GEN_1458 & _GEN_198;
  wire        _GEN_1464 = _GEN_1458 & _GEN_199;
  wire        _GEN_1465 = _GEN_1458 & _GEN_200;
  wire        _GEN_1466 = _GEN_1458 & _GEN_201;
  wire        _GEN_1467 = _GEN_1458 & _GEN_202;
  wire        _GEN_1468 = _GEN_1458 & _GEN_203;
  wire        _GEN_1469 = _GEN_1458 & _GEN_204;
  wire        _GEN_1470 = _GEN_1458 & _GEN_205;
  wire        _GEN_1471 = _GEN_1458 & _GEN_206;
  wire        _GEN_1472 = _GEN_1458 & _GEN_207;
  wire        _GEN_1473 = _GEN_1458 & _GEN_208;
  wire        _GEN_1474 = _GEN_1458 & _GEN_209;
  wire        _GEN_1475 = _GEN_1458 & _GEN_210;
  wire        _GEN_1476 = _GEN_1458 & _GEN_211;
  wire        _GEN_1477 = _GEN_1458 & _GEN_212;
  wire        _GEN_1478 = _GEN_1458 & _GEN_213;
  wire        _GEN_1479 = _GEN_1458 & _GEN_214;
  wire        _GEN_1480 = _GEN_1458 & _GEN_215;
  wire        _GEN_1481 = _GEN_1458 & _GEN_216;
  wire        _GEN_1482 = _GEN_1458 & _GEN_217;
  wire        _GEN_1483 = _GEN_1458 & _GEN_218;
  wire        _GEN_1484 = _GEN_1458 & _GEN_219;
  wire        _GEN_1485 = _GEN_1458 & _GEN_220;
  wire        _GEN_1486 = _GEN_1458 & _GEN_221;
  wire        _GEN_1487 = _GEN_1458 & _GEN_222;
  wire        _GEN_1488 = _GEN_1458 & _GEN_223;
  wire        _GEN_1489 = _GEN_1458 & _GEN_224;
  wire        _GEN_1490 = _GEN_1458 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_1491 = io_wb_resps_3_valid & io_wb_resps_3_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1492 = _GEN_258 | _GEN_1459;
  wire        _GEN_1493 = _GEN_260 | _GEN_1460;
  wire        _GEN_1494 = _GEN_262 | _GEN_1461;
  wire        _GEN_1495 = _GEN_264 | _GEN_1462;
  wire        _GEN_1496 = _GEN_266 | _GEN_1463;
  wire        _GEN_1497 = _GEN_268 | _GEN_1464;
  wire        _GEN_1498 = _GEN_270 | _GEN_1465;
  wire        _GEN_1499 = _GEN_272 | _GEN_1466;
  wire        _GEN_1500 = _GEN_274 | _GEN_1467;
  wire        _GEN_1501 = _GEN_276 | _GEN_1468;
  wire        _GEN_1502 = _GEN_278 | _GEN_1469;
  wire        _GEN_1503 = _GEN_280 | _GEN_1470;
  wire        _GEN_1504 = _GEN_282 | _GEN_1471;
  wire        _GEN_1505 = _GEN_284 | _GEN_1472;
  wire        _GEN_1506 = _GEN_286 | _GEN_1473;
  wire        _GEN_1507 = _GEN_288 | _GEN_1474;
  wire        _GEN_1508 = _GEN_290 | _GEN_1475;
  wire        _GEN_1509 = _GEN_292 | _GEN_1476;
  wire        _GEN_1510 = _GEN_294 | _GEN_1477;
  wire        _GEN_1511 = _GEN_296 | _GEN_1478;
  wire        _GEN_1512 = _GEN_298 | _GEN_1479;
  wire        _GEN_1513 = _GEN_300 | _GEN_1480;
  wire        _GEN_1514 = _GEN_302 | _GEN_1481;
  wire        _GEN_1515 = _GEN_304 | _GEN_1482;
  wire        _GEN_1516 = _GEN_306 | _GEN_1483;
  wire        _GEN_1517 = _GEN_308 | _GEN_1484;
  wire        _GEN_1518 = _GEN_310 | _GEN_1485;
  wire        _GEN_1519 = _GEN_312 | _GEN_1486;
  wire        _GEN_1520 = _GEN_314 | _GEN_1487;
  wire        _GEN_1521 = _GEN_316 | _GEN_1488;
  wire        _GEN_1522 = _GEN_318 | _GEN_1489;
  wire        _GEN_1523 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1490;
  wire        _GEN_1524 = io_wb_resps_4_valid & io_wb_resps_4_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1525 = _GEN_1524 & _GEN_322;
  wire        _GEN_1526 = _GEN_1524 & _GEN_323;
  wire        _GEN_1527 = _GEN_1524 & _GEN_324;
  wire        _GEN_1528 = _GEN_1524 & _GEN_325;
  wire        _GEN_1529 = _GEN_1524 & _GEN_326;
  wire        _GEN_1530 = _GEN_1524 & _GEN_327;
  wire        _GEN_1531 = _GEN_1524 & _GEN_328;
  wire        _GEN_1532 = _GEN_1524 & _GEN_329;
  wire        _GEN_1533 = _GEN_1524 & _GEN_330;
  wire        _GEN_1534 = _GEN_1524 & _GEN_331;
  wire        _GEN_1535 = _GEN_1524 & _GEN_332;
  wire        _GEN_1536 = _GEN_1524 & _GEN_333;
  wire        _GEN_1537 = _GEN_1524 & _GEN_334;
  wire        _GEN_1538 = _GEN_1524 & _GEN_335;
  wire        _GEN_1539 = _GEN_1524 & _GEN_336;
  wire        _GEN_1540 = _GEN_1524 & _GEN_337;
  wire        _GEN_1541 = _GEN_1524 & _GEN_338;
  wire        _GEN_1542 = _GEN_1524 & _GEN_339;
  wire        _GEN_1543 = _GEN_1524 & _GEN_340;
  wire        _GEN_1544 = _GEN_1524 & _GEN_341;
  wire        _GEN_1545 = _GEN_1524 & _GEN_342;
  wire        _GEN_1546 = _GEN_1524 & _GEN_343;
  wire        _GEN_1547 = _GEN_1524 & _GEN_344;
  wire        _GEN_1548 = _GEN_1524 & _GEN_345;
  wire        _GEN_1549 = _GEN_1524 & _GEN_346;
  wire        _GEN_1550 = _GEN_1524 & _GEN_347;
  wire        _GEN_1551 = _GEN_1524 & _GEN_348;
  wire        _GEN_1552 = _GEN_1524 & _GEN_349;
  wire        _GEN_1553 = _GEN_1524 & _GEN_350;
  wire        _GEN_1554 = _GEN_1524 & _GEN_351;
  wire        _GEN_1555 = _GEN_1524 & _GEN_352;
  wire        _GEN_1556 = _GEN_1524 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_1557 = io_wb_resps_5_valid & io_wb_resps_5_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1558 = _GEN_386 | _GEN_1525;
  wire        _GEN_1559 = _GEN_388 | _GEN_1526;
  wire        _GEN_1560 = _GEN_390 | _GEN_1527;
  wire        _GEN_1561 = _GEN_392 | _GEN_1528;
  wire        _GEN_1562 = _GEN_394 | _GEN_1529;
  wire        _GEN_1563 = _GEN_396 | _GEN_1530;
  wire        _GEN_1564 = _GEN_398 | _GEN_1531;
  wire        _GEN_1565 = _GEN_400 | _GEN_1532;
  wire        _GEN_1566 = _GEN_402 | _GEN_1533;
  wire        _GEN_1567 = _GEN_404 | _GEN_1534;
  wire        _GEN_1568 = _GEN_406 | _GEN_1535;
  wire        _GEN_1569 = _GEN_408 | _GEN_1536;
  wire        _GEN_1570 = _GEN_410 | _GEN_1537;
  wire        _GEN_1571 = _GEN_412 | _GEN_1538;
  wire        _GEN_1572 = _GEN_414 | _GEN_1539;
  wire        _GEN_1573 = _GEN_416 | _GEN_1540;
  wire        _GEN_1574 = _GEN_418 | _GEN_1541;
  wire        _GEN_1575 = _GEN_420 | _GEN_1542;
  wire        _GEN_1576 = _GEN_422 | _GEN_1543;
  wire        _GEN_1577 = _GEN_424 | _GEN_1544;
  wire        _GEN_1578 = _GEN_426 | _GEN_1545;
  wire        _GEN_1579 = _GEN_428 | _GEN_1546;
  wire        _GEN_1580 = _GEN_430 | _GEN_1547;
  wire        _GEN_1581 = _GEN_432 | _GEN_1548;
  wire        _GEN_1582 = _GEN_434 | _GEN_1549;
  wire        _GEN_1583 = _GEN_436 | _GEN_1550;
  wire        _GEN_1584 = _GEN_438 | _GEN_1551;
  wire        _GEN_1585 = _GEN_440 | _GEN_1552;
  wire        _GEN_1586 = _GEN_442 | _GEN_1553;
  wire        _GEN_1587 = _GEN_444 | _GEN_1554;
  wire        _GEN_1588 = _GEN_446 | _GEN_1555;
  wire        _GEN_1589 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1556;
  wire        _GEN_1590 = io_wb_resps_6_valid & io_wb_resps_6_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1591 = _GEN_1590 & _GEN_450;
  wire        _GEN_1592 = _GEN_1590 & _GEN_451;
  wire        _GEN_1593 = _GEN_1590 & _GEN_452;
  wire        _GEN_1594 = _GEN_1590 & _GEN_453;
  wire        _GEN_1595 = _GEN_1590 & _GEN_454;
  wire        _GEN_1596 = _GEN_1590 & _GEN_455;
  wire        _GEN_1597 = _GEN_1590 & _GEN_456;
  wire        _GEN_1598 = _GEN_1590 & _GEN_457;
  wire        _GEN_1599 = _GEN_1590 & _GEN_458;
  wire        _GEN_1600 = _GEN_1590 & _GEN_459;
  wire        _GEN_1601 = _GEN_1590 & _GEN_460;
  wire        _GEN_1602 = _GEN_1590 & _GEN_461;
  wire        _GEN_1603 = _GEN_1590 & _GEN_462;
  wire        _GEN_1604 = _GEN_1590 & _GEN_463;
  wire        _GEN_1605 = _GEN_1590 & _GEN_464;
  wire        _GEN_1606 = _GEN_1590 & _GEN_465;
  wire        _GEN_1607 = _GEN_1590 & _GEN_466;
  wire        _GEN_1608 = _GEN_1590 & _GEN_467;
  wire        _GEN_1609 = _GEN_1590 & _GEN_468;
  wire        _GEN_1610 = _GEN_1590 & _GEN_469;
  wire        _GEN_1611 = _GEN_1590 & _GEN_470;
  wire        _GEN_1612 = _GEN_1590 & _GEN_471;
  wire        _GEN_1613 = _GEN_1590 & _GEN_472;
  wire        _GEN_1614 = _GEN_1590 & _GEN_473;
  wire        _GEN_1615 = _GEN_1590 & _GEN_474;
  wire        _GEN_1616 = _GEN_1590 & _GEN_475;
  wire        _GEN_1617 = _GEN_1590 & _GEN_476;
  wire        _GEN_1618 = _GEN_1590 & _GEN_477;
  wire        _GEN_1619 = _GEN_1590 & _GEN_478;
  wire        _GEN_1620 = _GEN_1590 & _GEN_479;
  wire        _GEN_1621 = _GEN_1590 & _GEN_480;
  wire        _GEN_1622 = _GEN_1590 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_1623 = io_wb_resps_7_valid & io_wb_resps_7_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1624 = _GEN_514 | _GEN_1591;
  wire        _GEN_1625 = _GEN_516 | _GEN_1592;
  wire        _GEN_1626 = _GEN_518 | _GEN_1593;
  wire        _GEN_1627 = _GEN_520 | _GEN_1594;
  wire        _GEN_1628 = _GEN_522 | _GEN_1595;
  wire        _GEN_1629 = _GEN_524 | _GEN_1596;
  wire        _GEN_1630 = _GEN_526 | _GEN_1597;
  wire        _GEN_1631 = _GEN_528 | _GEN_1598;
  wire        _GEN_1632 = _GEN_530 | _GEN_1599;
  wire        _GEN_1633 = _GEN_532 | _GEN_1600;
  wire        _GEN_1634 = _GEN_534 | _GEN_1601;
  wire        _GEN_1635 = _GEN_536 | _GEN_1602;
  wire        _GEN_1636 = _GEN_538 | _GEN_1603;
  wire        _GEN_1637 = _GEN_540 | _GEN_1604;
  wire        _GEN_1638 = _GEN_542 | _GEN_1605;
  wire        _GEN_1639 = _GEN_544 | _GEN_1606;
  wire        _GEN_1640 = _GEN_546 | _GEN_1607;
  wire        _GEN_1641 = _GEN_548 | _GEN_1608;
  wire        _GEN_1642 = _GEN_550 | _GEN_1609;
  wire        _GEN_1643 = _GEN_552 | _GEN_1610;
  wire        _GEN_1644 = _GEN_554 | _GEN_1611;
  wire        _GEN_1645 = _GEN_556 | _GEN_1612;
  wire        _GEN_1646 = _GEN_558 | _GEN_1613;
  wire        _GEN_1647 = _GEN_560 | _GEN_1614;
  wire        _GEN_1648 = _GEN_562 | _GEN_1615;
  wire        _GEN_1649 = _GEN_564 | _GEN_1616;
  wire        _GEN_1650 = _GEN_566 | _GEN_1617;
  wire        _GEN_1651 = _GEN_568 | _GEN_1618;
  wire        _GEN_1652 = _GEN_570 | _GEN_1619;
  wire        _GEN_1653 = _GEN_572 | _GEN_1620;
  wire        _GEN_1654 = _GEN_574 | _GEN_1621;
  wire        _GEN_1655 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_1622;
  wire        _GEN_1656 = io_wb_resps_8_valid & io_wb_resps_8_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1657 = _GEN_1656 & _GEN_578;
  wire        _GEN_1658 = _GEN_1656 & _GEN_579;
  wire        _GEN_1659 = _GEN_1656 & _GEN_580;
  wire        _GEN_1660 = _GEN_1656 & _GEN_581;
  wire        _GEN_1661 = _GEN_1656 & _GEN_582;
  wire        _GEN_1662 = _GEN_1656 & _GEN_583;
  wire        _GEN_1663 = _GEN_1656 & _GEN_584;
  wire        _GEN_1664 = _GEN_1656 & _GEN_585;
  wire        _GEN_1665 = _GEN_1656 & _GEN_586;
  wire        _GEN_1666 = _GEN_1656 & _GEN_587;
  wire        _GEN_1667 = _GEN_1656 & _GEN_588;
  wire        _GEN_1668 = _GEN_1656 & _GEN_589;
  wire        _GEN_1669 = _GEN_1656 & _GEN_590;
  wire        _GEN_1670 = _GEN_1656 & _GEN_591;
  wire        _GEN_1671 = _GEN_1656 & _GEN_592;
  wire        _GEN_1672 = _GEN_1656 & _GEN_593;
  wire        _GEN_1673 = _GEN_1656 & _GEN_594;
  wire        _GEN_1674 = _GEN_1656 & _GEN_595;
  wire        _GEN_1675 = _GEN_1656 & _GEN_596;
  wire        _GEN_1676 = _GEN_1656 & _GEN_597;
  wire        _GEN_1677 = _GEN_1656 & _GEN_598;
  wire        _GEN_1678 = _GEN_1656 & _GEN_599;
  wire        _GEN_1679 = _GEN_1656 & _GEN_600;
  wire        _GEN_1680 = _GEN_1656 & _GEN_601;
  wire        _GEN_1681 = _GEN_1656 & _GEN_602;
  wire        _GEN_1682 = _GEN_1656 & _GEN_603;
  wire        _GEN_1683 = _GEN_1656 & _GEN_604;
  wire        _GEN_1684 = _GEN_1656 & _GEN_605;
  wire        _GEN_1685 = _GEN_1656 & _GEN_606;
  wire        _GEN_1686 = _GEN_1656 & _GEN_607;
  wire        _GEN_1687 = _GEN_1656 & _GEN_608;
  wire        _GEN_1688 = _GEN_1656 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_1689 = io_wb_resps_9_valid & io_wb_resps_9_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_1690 = _GEN_642 | _GEN_1657;
  wire        _GEN_1691 = _GEN_644 | _GEN_1658;
  wire        _GEN_1692 = _GEN_646 | _GEN_1659;
  wire        _GEN_1693 = _GEN_648 | _GEN_1660;
  wire        _GEN_1694 = _GEN_650 | _GEN_1661;
  wire        _GEN_1695 = _GEN_652 | _GEN_1662;
  wire        _GEN_1696 = _GEN_654 | _GEN_1663;
  wire        _GEN_1697 = _GEN_656 | _GEN_1664;
  wire        _GEN_1698 = _GEN_658 | _GEN_1665;
  wire        _GEN_1699 = _GEN_660 | _GEN_1666;
  wire        _GEN_1700 = _GEN_662 | _GEN_1667;
  wire        _GEN_1701 = _GEN_664 | _GEN_1668;
  wire        _GEN_1702 = _GEN_666 | _GEN_1669;
  wire        _GEN_1703 = _GEN_668 | _GEN_1670;
  wire        _GEN_1704 = _GEN_670 | _GEN_1671;
  wire        _GEN_1705 = _GEN_672 | _GEN_1672;
  wire        _GEN_1706 = _GEN_674 | _GEN_1673;
  wire        _GEN_1707 = _GEN_676 | _GEN_1674;
  wire        _GEN_1708 = _GEN_678 | _GEN_1675;
  wire        _GEN_1709 = _GEN_680 | _GEN_1676;
  wire        _GEN_1710 = _GEN_682 | _GEN_1677;
  wire        _GEN_1711 = _GEN_684 | _GEN_1678;
  wire        _GEN_1712 = _GEN_686 | _GEN_1679;
  wire        _GEN_1713 = _GEN_688 | _GEN_1680;
  wire        _GEN_1714 = _GEN_690 | _GEN_1681;
  wire        _GEN_1715 = _GEN_692 | _GEN_1682;
  wire        _GEN_1716 = _GEN_694 | _GEN_1683;
  wire        _GEN_1717 = _GEN_696 | _GEN_1684;
  wire        _GEN_1718 = _GEN_698 | _GEN_1685;
  wire        _GEN_1719 = _GEN_700 | _GEN_1686;
  wire        _GEN_1720 = _GEN_702 | _GEN_1687;
  wire        _GEN_1721 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1688;
  wire        _GEN_1722 = io_lsu_clr_bsy_0_valid & io_lsu_clr_bsy_0_bits[1:0] == 2'h2;
  wire        _GEN_1723 = _GEN_1722 & _GEN_706;
  wire        _GEN_1724 = _GEN_1722 & _GEN_707;
  wire        _GEN_1725 = _GEN_1722 & _GEN_708;
  wire        _GEN_1726 = _GEN_1722 & _GEN_709;
  wire        _GEN_1727 = _GEN_1722 & _GEN_710;
  wire        _GEN_1728 = _GEN_1722 & _GEN_711;
  wire        _GEN_1729 = _GEN_1722 & _GEN_712;
  wire        _GEN_1730 = _GEN_1722 & _GEN_713;
  wire        _GEN_1731 = _GEN_1722 & _GEN_714;
  wire        _GEN_1732 = _GEN_1722 & _GEN_715;
  wire        _GEN_1733 = _GEN_1722 & _GEN_716;
  wire        _GEN_1734 = _GEN_1722 & _GEN_717;
  wire        _GEN_1735 = _GEN_1722 & _GEN_718;
  wire        _GEN_1736 = _GEN_1722 & _GEN_719;
  wire        _GEN_1737 = _GEN_1722 & _GEN_720;
  wire        _GEN_1738 = _GEN_1722 & _GEN_721;
  wire        _GEN_1739 = _GEN_1722 & _GEN_722;
  wire        _GEN_1740 = _GEN_1722 & _GEN_723;
  wire        _GEN_1741 = _GEN_1722 & _GEN_724;
  wire        _GEN_1742 = _GEN_1722 & _GEN_725;
  wire        _GEN_1743 = _GEN_1722 & _GEN_726;
  wire        _GEN_1744 = _GEN_1722 & _GEN_727;
  wire        _GEN_1745 = _GEN_1722 & _GEN_728;
  wire        _GEN_1746 = _GEN_1722 & _GEN_729;
  wire        _GEN_1747 = _GEN_1722 & _GEN_730;
  wire        _GEN_1748 = _GEN_1722 & _GEN_731;
  wire        _GEN_1749 = _GEN_1722 & _GEN_732;
  wire        _GEN_1750 = _GEN_1722 & _GEN_733;
  wire        _GEN_1751 = _GEN_1722 & _GEN_734;
  wire        _GEN_1752 = _GEN_1722 & _GEN_735;
  wire        _GEN_1753 = _GEN_1722 & _GEN_736;
  wire        _GEN_1754 = _GEN_1722 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_1755 = io_lsu_clr_bsy_1_valid & io_lsu_clr_bsy_1_bits[1:0] == 2'h2;
  wire        _GEN_1756 = _GEN_770 | _GEN_1723;
  wire        _GEN_1757 = _GEN_772 | _GEN_1724;
  wire        _GEN_1758 = _GEN_774 | _GEN_1725;
  wire        _GEN_1759 = _GEN_776 | _GEN_1726;
  wire        _GEN_1760 = _GEN_778 | _GEN_1727;
  wire        _GEN_1761 = _GEN_780 | _GEN_1728;
  wire        _GEN_1762 = _GEN_782 | _GEN_1729;
  wire        _GEN_1763 = _GEN_784 | _GEN_1730;
  wire        _GEN_1764 = _GEN_786 | _GEN_1731;
  wire        _GEN_1765 = _GEN_788 | _GEN_1732;
  wire        _GEN_1766 = _GEN_790 | _GEN_1733;
  wire        _GEN_1767 = _GEN_792 | _GEN_1734;
  wire        _GEN_1768 = _GEN_794 | _GEN_1735;
  wire        _GEN_1769 = _GEN_796 | _GEN_1736;
  wire        _GEN_1770 = _GEN_798 | _GEN_1737;
  wire        _GEN_1771 = _GEN_800 | _GEN_1738;
  wire        _GEN_1772 = _GEN_802 | _GEN_1739;
  wire        _GEN_1773 = _GEN_804 | _GEN_1740;
  wire        _GEN_1774 = _GEN_806 | _GEN_1741;
  wire        _GEN_1775 = _GEN_808 | _GEN_1742;
  wire        _GEN_1776 = _GEN_810 | _GEN_1743;
  wire        _GEN_1777 = _GEN_812 | _GEN_1744;
  wire        _GEN_1778 = _GEN_814 | _GEN_1745;
  wire        _GEN_1779 = _GEN_816 | _GEN_1746;
  wire        _GEN_1780 = _GEN_818 | _GEN_1747;
  wire        _GEN_1781 = _GEN_820 | _GEN_1748;
  wire        _GEN_1782 = _GEN_822 | _GEN_1749;
  wire        _GEN_1783 = _GEN_824 | _GEN_1750;
  wire        _GEN_1784 = _GEN_826 | _GEN_1751;
  wire        _GEN_1785 = _GEN_828 | _GEN_1752;
  wire        _GEN_1786 = _GEN_830 | _GEN_1753;
  wire        _GEN_1787 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_1754;
  wire        _GEN_1788 = io_lsu_clr_bsy_2_valid & io_lsu_clr_bsy_2_bits[1:0] == 2'h2;
  wire        _GEN_1789 = _GEN_1788 & _GEN_834;
  wire        _GEN_1790 = _GEN_1788 & _GEN_835;
  wire        _GEN_1791 = _GEN_1788 & _GEN_836;
  wire        _GEN_1792 = _GEN_1788 & _GEN_837;
  wire        _GEN_1793 = _GEN_1788 & _GEN_838;
  wire        _GEN_1794 = _GEN_1788 & _GEN_839;
  wire        _GEN_1795 = _GEN_1788 & _GEN_840;
  wire        _GEN_1796 = _GEN_1788 & _GEN_841;
  wire        _GEN_1797 = _GEN_1788 & _GEN_842;
  wire        _GEN_1798 = _GEN_1788 & _GEN_843;
  wire        _GEN_1799 = _GEN_1788 & _GEN_844;
  wire        _GEN_1800 = _GEN_1788 & _GEN_845;
  wire        _GEN_1801 = _GEN_1788 & _GEN_846;
  wire        _GEN_1802 = _GEN_1788 & _GEN_847;
  wire        _GEN_1803 = _GEN_1788 & _GEN_848;
  wire        _GEN_1804 = _GEN_1788 & _GEN_849;
  wire        _GEN_1805 = _GEN_1788 & _GEN_850;
  wire        _GEN_1806 = _GEN_1788 & _GEN_851;
  wire        _GEN_1807 = _GEN_1788 & _GEN_852;
  wire        _GEN_1808 = _GEN_1788 & _GEN_853;
  wire        _GEN_1809 = _GEN_1788 & _GEN_854;
  wire        _GEN_1810 = _GEN_1788 & _GEN_855;
  wire        _GEN_1811 = _GEN_1788 & _GEN_856;
  wire        _GEN_1812 = _GEN_1788 & _GEN_857;
  wire        _GEN_1813 = _GEN_1788 & _GEN_858;
  wire        _GEN_1814 = _GEN_1788 & _GEN_859;
  wire        _GEN_1815 = _GEN_1788 & _GEN_860;
  wire        _GEN_1816 = _GEN_1788 & _GEN_861;
  wire        _GEN_1817 = _GEN_1788 & _GEN_862;
  wire        _GEN_1818 = _GEN_1788 & _GEN_863;
  wire        _GEN_1819 = _GEN_1788 & _GEN_864;
  wire        _GEN_1820 = _GEN_1788 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_1821 = io_lxcpt_valid & io_lxcpt_bits_uop_rob_idx[1:0] == 2'h2;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_51 = rob_predicated_2_0;
      5'b00001:
        casez_tmp_51 = rob_predicated_2_1;
      5'b00010:
        casez_tmp_51 = rob_predicated_2_2;
      5'b00011:
        casez_tmp_51 = rob_predicated_2_3;
      5'b00100:
        casez_tmp_51 = rob_predicated_2_4;
      5'b00101:
        casez_tmp_51 = rob_predicated_2_5;
      5'b00110:
        casez_tmp_51 = rob_predicated_2_6;
      5'b00111:
        casez_tmp_51 = rob_predicated_2_7;
      5'b01000:
        casez_tmp_51 = rob_predicated_2_8;
      5'b01001:
        casez_tmp_51 = rob_predicated_2_9;
      5'b01010:
        casez_tmp_51 = rob_predicated_2_10;
      5'b01011:
        casez_tmp_51 = rob_predicated_2_11;
      5'b01100:
        casez_tmp_51 = rob_predicated_2_12;
      5'b01101:
        casez_tmp_51 = rob_predicated_2_13;
      5'b01110:
        casez_tmp_51 = rob_predicated_2_14;
      5'b01111:
        casez_tmp_51 = rob_predicated_2_15;
      5'b10000:
        casez_tmp_51 = rob_predicated_2_16;
      5'b10001:
        casez_tmp_51 = rob_predicated_2_17;
      5'b10010:
        casez_tmp_51 = rob_predicated_2_18;
      5'b10011:
        casez_tmp_51 = rob_predicated_2_19;
      5'b10100:
        casez_tmp_51 = rob_predicated_2_20;
      5'b10101:
        casez_tmp_51 = rob_predicated_2_21;
      5'b10110:
        casez_tmp_51 = rob_predicated_2_22;
      5'b10111:
        casez_tmp_51 = rob_predicated_2_23;
      5'b11000:
        casez_tmp_51 = rob_predicated_2_24;
      5'b11001:
        casez_tmp_51 = rob_predicated_2_25;
      5'b11010:
        casez_tmp_51 = rob_predicated_2_26;
      5'b11011:
        casez_tmp_51 = rob_predicated_2_27;
      5'b11100:
        casez_tmp_51 = rob_predicated_2_28;
      5'b11101:
        casez_tmp_51 = rob_predicated_2_29;
      5'b11110:
        casez_tmp_51 = rob_predicated_2_30;
      default:
        casez_tmp_51 = rob_predicated_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_52 = rob_uop_2_0_uopc;
      5'b00001:
        casez_tmp_52 = rob_uop_2_1_uopc;
      5'b00010:
        casez_tmp_52 = rob_uop_2_2_uopc;
      5'b00011:
        casez_tmp_52 = rob_uop_2_3_uopc;
      5'b00100:
        casez_tmp_52 = rob_uop_2_4_uopc;
      5'b00101:
        casez_tmp_52 = rob_uop_2_5_uopc;
      5'b00110:
        casez_tmp_52 = rob_uop_2_6_uopc;
      5'b00111:
        casez_tmp_52 = rob_uop_2_7_uopc;
      5'b01000:
        casez_tmp_52 = rob_uop_2_8_uopc;
      5'b01001:
        casez_tmp_52 = rob_uop_2_9_uopc;
      5'b01010:
        casez_tmp_52 = rob_uop_2_10_uopc;
      5'b01011:
        casez_tmp_52 = rob_uop_2_11_uopc;
      5'b01100:
        casez_tmp_52 = rob_uop_2_12_uopc;
      5'b01101:
        casez_tmp_52 = rob_uop_2_13_uopc;
      5'b01110:
        casez_tmp_52 = rob_uop_2_14_uopc;
      5'b01111:
        casez_tmp_52 = rob_uop_2_15_uopc;
      5'b10000:
        casez_tmp_52 = rob_uop_2_16_uopc;
      5'b10001:
        casez_tmp_52 = rob_uop_2_17_uopc;
      5'b10010:
        casez_tmp_52 = rob_uop_2_18_uopc;
      5'b10011:
        casez_tmp_52 = rob_uop_2_19_uopc;
      5'b10100:
        casez_tmp_52 = rob_uop_2_20_uopc;
      5'b10101:
        casez_tmp_52 = rob_uop_2_21_uopc;
      5'b10110:
        casez_tmp_52 = rob_uop_2_22_uopc;
      5'b10111:
        casez_tmp_52 = rob_uop_2_23_uopc;
      5'b11000:
        casez_tmp_52 = rob_uop_2_24_uopc;
      5'b11001:
        casez_tmp_52 = rob_uop_2_25_uopc;
      5'b11010:
        casez_tmp_52 = rob_uop_2_26_uopc;
      5'b11011:
        casez_tmp_52 = rob_uop_2_27_uopc;
      5'b11100:
        casez_tmp_52 = rob_uop_2_28_uopc;
      5'b11101:
        casez_tmp_52 = rob_uop_2_29_uopc;
      5'b11110:
        casez_tmp_52 = rob_uop_2_30_uopc;
      default:
        casez_tmp_52 = rob_uop_2_31_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_53 = rob_uop_2_0_is_rvc;
      5'b00001:
        casez_tmp_53 = rob_uop_2_1_is_rvc;
      5'b00010:
        casez_tmp_53 = rob_uop_2_2_is_rvc;
      5'b00011:
        casez_tmp_53 = rob_uop_2_3_is_rvc;
      5'b00100:
        casez_tmp_53 = rob_uop_2_4_is_rvc;
      5'b00101:
        casez_tmp_53 = rob_uop_2_5_is_rvc;
      5'b00110:
        casez_tmp_53 = rob_uop_2_6_is_rvc;
      5'b00111:
        casez_tmp_53 = rob_uop_2_7_is_rvc;
      5'b01000:
        casez_tmp_53 = rob_uop_2_8_is_rvc;
      5'b01001:
        casez_tmp_53 = rob_uop_2_9_is_rvc;
      5'b01010:
        casez_tmp_53 = rob_uop_2_10_is_rvc;
      5'b01011:
        casez_tmp_53 = rob_uop_2_11_is_rvc;
      5'b01100:
        casez_tmp_53 = rob_uop_2_12_is_rvc;
      5'b01101:
        casez_tmp_53 = rob_uop_2_13_is_rvc;
      5'b01110:
        casez_tmp_53 = rob_uop_2_14_is_rvc;
      5'b01111:
        casez_tmp_53 = rob_uop_2_15_is_rvc;
      5'b10000:
        casez_tmp_53 = rob_uop_2_16_is_rvc;
      5'b10001:
        casez_tmp_53 = rob_uop_2_17_is_rvc;
      5'b10010:
        casez_tmp_53 = rob_uop_2_18_is_rvc;
      5'b10011:
        casez_tmp_53 = rob_uop_2_19_is_rvc;
      5'b10100:
        casez_tmp_53 = rob_uop_2_20_is_rvc;
      5'b10101:
        casez_tmp_53 = rob_uop_2_21_is_rvc;
      5'b10110:
        casez_tmp_53 = rob_uop_2_22_is_rvc;
      5'b10111:
        casez_tmp_53 = rob_uop_2_23_is_rvc;
      5'b11000:
        casez_tmp_53 = rob_uop_2_24_is_rvc;
      5'b11001:
        casez_tmp_53 = rob_uop_2_25_is_rvc;
      5'b11010:
        casez_tmp_53 = rob_uop_2_26_is_rvc;
      5'b11011:
        casez_tmp_53 = rob_uop_2_27_is_rvc;
      5'b11100:
        casez_tmp_53 = rob_uop_2_28_is_rvc;
      5'b11101:
        casez_tmp_53 = rob_uop_2_29_is_rvc;
      5'b11110:
        casez_tmp_53 = rob_uop_2_30_is_rvc;
      default:
        casez_tmp_53 = rob_uop_2_31_is_rvc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_54 = rob_uop_2_0_ftq_idx;
      5'b00001:
        casez_tmp_54 = rob_uop_2_1_ftq_idx;
      5'b00010:
        casez_tmp_54 = rob_uop_2_2_ftq_idx;
      5'b00011:
        casez_tmp_54 = rob_uop_2_3_ftq_idx;
      5'b00100:
        casez_tmp_54 = rob_uop_2_4_ftq_idx;
      5'b00101:
        casez_tmp_54 = rob_uop_2_5_ftq_idx;
      5'b00110:
        casez_tmp_54 = rob_uop_2_6_ftq_idx;
      5'b00111:
        casez_tmp_54 = rob_uop_2_7_ftq_idx;
      5'b01000:
        casez_tmp_54 = rob_uop_2_8_ftq_idx;
      5'b01001:
        casez_tmp_54 = rob_uop_2_9_ftq_idx;
      5'b01010:
        casez_tmp_54 = rob_uop_2_10_ftq_idx;
      5'b01011:
        casez_tmp_54 = rob_uop_2_11_ftq_idx;
      5'b01100:
        casez_tmp_54 = rob_uop_2_12_ftq_idx;
      5'b01101:
        casez_tmp_54 = rob_uop_2_13_ftq_idx;
      5'b01110:
        casez_tmp_54 = rob_uop_2_14_ftq_idx;
      5'b01111:
        casez_tmp_54 = rob_uop_2_15_ftq_idx;
      5'b10000:
        casez_tmp_54 = rob_uop_2_16_ftq_idx;
      5'b10001:
        casez_tmp_54 = rob_uop_2_17_ftq_idx;
      5'b10010:
        casez_tmp_54 = rob_uop_2_18_ftq_idx;
      5'b10011:
        casez_tmp_54 = rob_uop_2_19_ftq_idx;
      5'b10100:
        casez_tmp_54 = rob_uop_2_20_ftq_idx;
      5'b10101:
        casez_tmp_54 = rob_uop_2_21_ftq_idx;
      5'b10110:
        casez_tmp_54 = rob_uop_2_22_ftq_idx;
      5'b10111:
        casez_tmp_54 = rob_uop_2_23_ftq_idx;
      5'b11000:
        casez_tmp_54 = rob_uop_2_24_ftq_idx;
      5'b11001:
        casez_tmp_54 = rob_uop_2_25_ftq_idx;
      5'b11010:
        casez_tmp_54 = rob_uop_2_26_ftq_idx;
      5'b11011:
        casez_tmp_54 = rob_uop_2_27_ftq_idx;
      5'b11100:
        casez_tmp_54 = rob_uop_2_28_ftq_idx;
      5'b11101:
        casez_tmp_54 = rob_uop_2_29_ftq_idx;
      5'b11110:
        casez_tmp_54 = rob_uop_2_30_ftq_idx;
      default:
        casez_tmp_54 = rob_uop_2_31_ftq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_55 = rob_uop_2_0_edge_inst;
      5'b00001:
        casez_tmp_55 = rob_uop_2_1_edge_inst;
      5'b00010:
        casez_tmp_55 = rob_uop_2_2_edge_inst;
      5'b00011:
        casez_tmp_55 = rob_uop_2_3_edge_inst;
      5'b00100:
        casez_tmp_55 = rob_uop_2_4_edge_inst;
      5'b00101:
        casez_tmp_55 = rob_uop_2_5_edge_inst;
      5'b00110:
        casez_tmp_55 = rob_uop_2_6_edge_inst;
      5'b00111:
        casez_tmp_55 = rob_uop_2_7_edge_inst;
      5'b01000:
        casez_tmp_55 = rob_uop_2_8_edge_inst;
      5'b01001:
        casez_tmp_55 = rob_uop_2_9_edge_inst;
      5'b01010:
        casez_tmp_55 = rob_uop_2_10_edge_inst;
      5'b01011:
        casez_tmp_55 = rob_uop_2_11_edge_inst;
      5'b01100:
        casez_tmp_55 = rob_uop_2_12_edge_inst;
      5'b01101:
        casez_tmp_55 = rob_uop_2_13_edge_inst;
      5'b01110:
        casez_tmp_55 = rob_uop_2_14_edge_inst;
      5'b01111:
        casez_tmp_55 = rob_uop_2_15_edge_inst;
      5'b10000:
        casez_tmp_55 = rob_uop_2_16_edge_inst;
      5'b10001:
        casez_tmp_55 = rob_uop_2_17_edge_inst;
      5'b10010:
        casez_tmp_55 = rob_uop_2_18_edge_inst;
      5'b10011:
        casez_tmp_55 = rob_uop_2_19_edge_inst;
      5'b10100:
        casez_tmp_55 = rob_uop_2_20_edge_inst;
      5'b10101:
        casez_tmp_55 = rob_uop_2_21_edge_inst;
      5'b10110:
        casez_tmp_55 = rob_uop_2_22_edge_inst;
      5'b10111:
        casez_tmp_55 = rob_uop_2_23_edge_inst;
      5'b11000:
        casez_tmp_55 = rob_uop_2_24_edge_inst;
      5'b11001:
        casez_tmp_55 = rob_uop_2_25_edge_inst;
      5'b11010:
        casez_tmp_55 = rob_uop_2_26_edge_inst;
      5'b11011:
        casez_tmp_55 = rob_uop_2_27_edge_inst;
      5'b11100:
        casez_tmp_55 = rob_uop_2_28_edge_inst;
      5'b11101:
        casez_tmp_55 = rob_uop_2_29_edge_inst;
      5'b11110:
        casez_tmp_55 = rob_uop_2_30_edge_inst;
      default:
        casez_tmp_55 = rob_uop_2_31_edge_inst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_56 = rob_uop_2_0_pc_lob;
      5'b00001:
        casez_tmp_56 = rob_uop_2_1_pc_lob;
      5'b00010:
        casez_tmp_56 = rob_uop_2_2_pc_lob;
      5'b00011:
        casez_tmp_56 = rob_uop_2_3_pc_lob;
      5'b00100:
        casez_tmp_56 = rob_uop_2_4_pc_lob;
      5'b00101:
        casez_tmp_56 = rob_uop_2_5_pc_lob;
      5'b00110:
        casez_tmp_56 = rob_uop_2_6_pc_lob;
      5'b00111:
        casez_tmp_56 = rob_uop_2_7_pc_lob;
      5'b01000:
        casez_tmp_56 = rob_uop_2_8_pc_lob;
      5'b01001:
        casez_tmp_56 = rob_uop_2_9_pc_lob;
      5'b01010:
        casez_tmp_56 = rob_uop_2_10_pc_lob;
      5'b01011:
        casez_tmp_56 = rob_uop_2_11_pc_lob;
      5'b01100:
        casez_tmp_56 = rob_uop_2_12_pc_lob;
      5'b01101:
        casez_tmp_56 = rob_uop_2_13_pc_lob;
      5'b01110:
        casez_tmp_56 = rob_uop_2_14_pc_lob;
      5'b01111:
        casez_tmp_56 = rob_uop_2_15_pc_lob;
      5'b10000:
        casez_tmp_56 = rob_uop_2_16_pc_lob;
      5'b10001:
        casez_tmp_56 = rob_uop_2_17_pc_lob;
      5'b10010:
        casez_tmp_56 = rob_uop_2_18_pc_lob;
      5'b10011:
        casez_tmp_56 = rob_uop_2_19_pc_lob;
      5'b10100:
        casez_tmp_56 = rob_uop_2_20_pc_lob;
      5'b10101:
        casez_tmp_56 = rob_uop_2_21_pc_lob;
      5'b10110:
        casez_tmp_56 = rob_uop_2_22_pc_lob;
      5'b10111:
        casez_tmp_56 = rob_uop_2_23_pc_lob;
      5'b11000:
        casez_tmp_56 = rob_uop_2_24_pc_lob;
      5'b11001:
        casez_tmp_56 = rob_uop_2_25_pc_lob;
      5'b11010:
        casez_tmp_56 = rob_uop_2_26_pc_lob;
      5'b11011:
        casez_tmp_56 = rob_uop_2_27_pc_lob;
      5'b11100:
        casez_tmp_56 = rob_uop_2_28_pc_lob;
      5'b11101:
        casez_tmp_56 = rob_uop_2_29_pc_lob;
      5'b11110:
        casez_tmp_56 = rob_uop_2_30_pc_lob;
      default:
        casez_tmp_56 = rob_uop_2_31_pc_lob;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_57 = rob_uop_2_0_pdst;
      5'b00001:
        casez_tmp_57 = rob_uop_2_1_pdst;
      5'b00010:
        casez_tmp_57 = rob_uop_2_2_pdst;
      5'b00011:
        casez_tmp_57 = rob_uop_2_3_pdst;
      5'b00100:
        casez_tmp_57 = rob_uop_2_4_pdst;
      5'b00101:
        casez_tmp_57 = rob_uop_2_5_pdst;
      5'b00110:
        casez_tmp_57 = rob_uop_2_6_pdst;
      5'b00111:
        casez_tmp_57 = rob_uop_2_7_pdst;
      5'b01000:
        casez_tmp_57 = rob_uop_2_8_pdst;
      5'b01001:
        casez_tmp_57 = rob_uop_2_9_pdst;
      5'b01010:
        casez_tmp_57 = rob_uop_2_10_pdst;
      5'b01011:
        casez_tmp_57 = rob_uop_2_11_pdst;
      5'b01100:
        casez_tmp_57 = rob_uop_2_12_pdst;
      5'b01101:
        casez_tmp_57 = rob_uop_2_13_pdst;
      5'b01110:
        casez_tmp_57 = rob_uop_2_14_pdst;
      5'b01111:
        casez_tmp_57 = rob_uop_2_15_pdst;
      5'b10000:
        casez_tmp_57 = rob_uop_2_16_pdst;
      5'b10001:
        casez_tmp_57 = rob_uop_2_17_pdst;
      5'b10010:
        casez_tmp_57 = rob_uop_2_18_pdst;
      5'b10011:
        casez_tmp_57 = rob_uop_2_19_pdst;
      5'b10100:
        casez_tmp_57 = rob_uop_2_20_pdst;
      5'b10101:
        casez_tmp_57 = rob_uop_2_21_pdst;
      5'b10110:
        casez_tmp_57 = rob_uop_2_22_pdst;
      5'b10111:
        casez_tmp_57 = rob_uop_2_23_pdst;
      5'b11000:
        casez_tmp_57 = rob_uop_2_24_pdst;
      5'b11001:
        casez_tmp_57 = rob_uop_2_25_pdst;
      5'b11010:
        casez_tmp_57 = rob_uop_2_26_pdst;
      5'b11011:
        casez_tmp_57 = rob_uop_2_27_pdst;
      5'b11100:
        casez_tmp_57 = rob_uop_2_28_pdst;
      5'b11101:
        casez_tmp_57 = rob_uop_2_29_pdst;
      5'b11110:
        casez_tmp_57 = rob_uop_2_30_pdst;
      default:
        casez_tmp_57 = rob_uop_2_31_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_58 = rob_uop_2_0_stale_pdst;
      5'b00001:
        casez_tmp_58 = rob_uop_2_1_stale_pdst;
      5'b00010:
        casez_tmp_58 = rob_uop_2_2_stale_pdst;
      5'b00011:
        casez_tmp_58 = rob_uop_2_3_stale_pdst;
      5'b00100:
        casez_tmp_58 = rob_uop_2_4_stale_pdst;
      5'b00101:
        casez_tmp_58 = rob_uop_2_5_stale_pdst;
      5'b00110:
        casez_tmp_58 = rob_uop_2_6_stale_pdst;
      5'b00111:
        casez_tmp_58 = rob_uop_2_7_stale_pdst;
      5'b01000:
        casez_tmp_58 = rob_uop_2_8_stale_pdst;
      5'b01001:
        casez_tmp_58 = rob_uop_2_9_stale_pdst;
      5'b01010:
        casez_tmp_58 = rob_uop_2_10_stale_pdst;
      5'b01011:
        casez_tmp_58 = rob_uop_2_11_stale_pdst;
      5'b01100:
        casez_tmp_58 = rob_uop_2_12_stale_pdst;
      5'b01101:
        casez_tmp_58 = rob_uop_2_13_stale_pdst;
      5'b01110:
        casez_tmp_58 = rob_uop_2_14_stale_pdst;
      5'b01111:
        casez_tmp_58 = rob_uop_2_15_stale_pdst;
      5'b10000:
        casez_tmp_58 = rob_uop_2_16_stale_pdst;
      5'b10001:
        casez_tmp_58 = rob_uop_2_17_stale_pdst;
      5'b10010:
        casez_tmp_58 = rob_uop_2_18_stale_pdst;
      5'b10011:
        casez_tmp_58 = rob_uop_2_19_stale_pdst;
      5'b10100:
        casez_tmp_58 = rob_uop_2_20_stale_pdst;
      5'b10101:
        casez_tmp_58 = rob_uop_2_21_stale_pdst;
      5'b10110:
        casez_tmp_58 = rob_uop_2_22_stale_pdst;
      5'b10111:
        casez_tmp_58 = rob_uop_2_23_stale_pdst;
      5'b11000:
        casez_tmp_58 = rob_uop_2_24_stale_pdst;
      5'b11001:
        casez_tmp_58 = rob_uop_2_25_stale_pdst;
      5'b11010:
        casez_tmp_58 = rob_uop_2_26_stale_pdst;
      5'b11011:
        casez_tmp_58 = rob_uop_2_27_stale_pdst;
      5'b11100:
        casez_tmp_58 = rob_uop_2_28_stale_pdst;
      5'b11101:
        casez_tmp_58 = rob_uop_2_29_stale_pdst;
      5'b11110:
        casez_tmp_58 = rob_uop_2_30_stale_pdst;
      default:
        casez_tmp_58 = rob_uop_2_31_stale_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_59 = rob_uop_2_0_is_fencei;
      5'b00001:
        casez_tmp_59 = rob_uop_2_1_is_fencei;
      5'b00010:
        casez_tmp_59 = rob_uop_2_2_is_fencei;
      5'b00011:
        casez_tmp_59 = rob_uop_2_3_is_fencei;
      5'b00100:
        casez_tmp_59 = rob_uop_2_4_is_fencei;
      5'b00101:
        casez_tmp_59 = rob_uop_2_5_is_fencei;
      5'b00110:
        casez_tmp_59 = rob_uop_2_6_is_fencei;
      5'b00111:
        casez_tmp_59 = rob_uop_2_7_is_fencei;
      5'b01000:
        casez_tmp_59 = rob_uop_2_8_is_fencei;
      5'b01001:
        casez_tmp_59 = rob_uop_2_9_is_fencei;
      5'b01010:
        casez_tmp_59 = rob_uop_2_10_is_fencei;
      5'b01011:
        casez_tmp_59 = rob_uop_2_11_is_fencei;
      5'b01100:
        casez_tmp_59 = rob_uop_2_12_is_fencei;
      5'b01101:
        casez_tmp_59 = rob_uop_2_13_is_fencei;
      5'b01110:
        casez_tmp_59 = rob_uop_2_14_is_fencei;
      5'b01111:
        casez_tmp_59 = rob_uop_2_15_is_fencei;
      5'b10000:
        casez_tmp_59 = rob_uop_2_16_is_fencei;
      5'b10001:
        casez_tmp_59 = rob_uop_2_17_is_fencei;
      5'b10010:
        casez_tmp_59 = rob_uop_2_18_is_fencei;
      5'b10011:
        casez_tmp_59 = rob_uop_2_19_is_fencei;
      5'b10100:
        casez_tmp_59 = rob_uop_2_20_is_fencei;
      5'b10101:
        casez_tmp_59 = rob_uop_2_21_is_fencei;
      5'b10110:
        casez_tmp_59 = rob_uop_2_22_is_fencei;
      5'b10111:
        casez_tmp_59 = rob_uop_2_23_is_fencei;
      5'b11000:
        casez_tmp_59 = rob_uop_2_24_is_fencei;
      5'b11001:
        casez_tmp_59 = rob_uop_2_25_is_fencei;
      5'b11010:
        casez_tmp_59 = rob_uop_2_26_is_fencei;
      5'b11011:
        casez_tmp_59 = rob_uop_2_27_is_fencei;
      5'b11100:
        casez_tmp_59 = rob_uop_2_28_is_fencei;
      5'b11101:
        casez_tmp_59 = rob_uop_2_29_is_fencei;
      5'b11110:
        casez_tmp_59 = rob_uop_2_30_is_fencei;
      default:
        casez_tmp_59 = rob_uop_2_31_is_fencei;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_60 = rob_uop_2_0_uses_ldq;
      5'b00001:
        casez_tmp_60 = rob_uop_2_1_uses_ldq;
      5'b00010:
        casez_tmp_60 = rob_uop_2_2_uses_ldq;
      5'b00011:
        casez_tmp_60 = rob_uop_2_3_uses_ldq;
      5'b00100:
        casez_tmp_60 = rob_uop_2_4_uses_ldq;
      5'b00101:
        casez_tmp_60 = rob_uop_2_5_uses_ldq;
      5'b00110:
        casez_tmp_60 = rob_uop_2_6_uses_ldq;
      5'b00111:
        casez_tmp_60 = rob_uop_2_7_uses_ldq;
      5'b01000:
        casez_tmp_60 = rob_uop_2_8_uses_ldq;
      5'b01001:
        casez_tmp_60 = rob_uop_2_9_uses_ldq;
      5'b01010:
        casez_tmp_60 = rob_uop_2_10_uses_ldq;
      5'b01011:
        casez_tmp_60 = rob_uop_2_11_uses_ldq;
      5'b01100:
        casez_tmp_60 = rob_uop_2_12_uses_ldq;
      5'b01101:
        casez_tmp_60 = rob_uop_2_13_uses_ldq;
      5'b01110:
        casez_tmp_60 = rob_uop_2_14_uses_ldq;
      5'b01111:
        casez_tmp_60 = rob_uop_2_15_uses_ldq;
      5'b10000:
        casez_tmp_60 = rob_uop_2_16_uses_ldq;
      5'b10001:
        casez_tmp_60 = rob_uop_2_17_uses_ldq;
      5'b10010:
        casez_tmp_60 = rob_uop_2_18_uses_ldq;
      5'b10011:
        casez_tmp_60 = rob_uop_2_19_uses_ldq;
      5'b10100:
        casez_tmp_60 = rob_uop_2_20_uses_ldq;
      5'b10101:
        casez_tmp_60 = rob_uop_2_21_uses_ldq;
      5'b10110:
        casez_tmp_60 = rob_uop_2_22_uses_ldq;
      5'b10111:
        casez_tmp_60 = rob_uop_2_23_uses_ldq;
      5'b11000:
        casez_tmp_60 = rob_uop_2_24_uses_ldq;
      5'b11001:
        casez_tmp_60 = rob_uop_2_25_uses_ldq;
      5'b11010:
        casez_tmp_60 = rob_uop_2_26_uses_ldq;
      5'b11011:
        casez_tmp_60 = rob_uop_2_27_uses_ldq;
      5'b11100:
        casez_tmp_60 = rob_uop_2_28_uses_ldq;
      5'b11101:
        casez_tmp_60 = rob_uop_2_29_uses_ldq;
      5'b11110:
        casez_tmp_60 = rob_uop_2_30_uses_ldq;
      default:
        casez_tmp_60 = rob_uop_2_31_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_61 = rob_uop_2_0_uses_stq;
      5'b00001:
        casez_tmp_61 = rob_uop_2_1_uses_stq;
      5'b00010:
        casez_tmp_61 = rob_uop_2_2_uses_stq;
      5'b00011:
        casez_tmp_61 = rob_uop_2_3_uses_stq;
      5'b00100:
        casez_tmp_61 = rob_uop_2_4_uses_stq;
      5'b00101:
        casez_tmp_61 = rob_uop_2_5_uses_stq;
      5'b00110:
        casez_tmp_61 = rob_uop_2_6_uses_stq;
      5'b00111:
        casez_tmp_61 = rob_uop_2_7_uses_stq;
      5'b01000:
        casez_tmp_61 = rob_uop_2_8_uses_stq;
      5'b01001:
        casez_tmp_61 = rob_uop_2_9_uses_stq;
      5'b01010:
        casez_tmp_61 = rob_uop_2_10_uses_stq;
      5'b01011:
        casez_tmp_61 = rob_uop_2_11_uses_stq;
      5'b01100:
        casez_tmp_61 = rob_uop_2_12_uses_stq;
      5'b01101:
        casez_tmp_61 = rob_uop_2_13_uses_stq;
      5'b01110:
        casez_tmp_61 = rob_uop_2_14_uses_stq;
      5'b01111:
        casez_tmp_61 = rob_uop_2_15_uses_stq;
      5'b10000:
        casez_tmp_61 = rob_uop_2_16_uses_stq;
      5'b10001:
        casez_tmp_61 = rob_uop_2_17_uses_stq;
      5'b10010:
        casez_tmp_61 = rob_uop_2_18_uses_stq;
      5'b10011:
        casez_tmp_61 = rob_uop_2_19_uses_stq;
      5'b10100:
        casez_tmp_61 = rob_uop_2_20_uses_stq;
      5'b10101:
        casez_tmp_61 = rob_uop_2_21_uses_stq;
      5'b10110:
        casez_tmp_61 = rob_uop_2_22_uses_stq;
      5'b10111:
        casez_tmp_61 = rob_uop_2_23_uses_stq;
      5'b11000:
        casez_tmp_61 = rob_uop_2_24_uses_stq;
      5'b11001:
        casez_tmp_61 = rob_uop_2_25_uses_stq;
      5'b11010:
        casez_tmp_61 = rob_uop_2_26_uses_stq;
      5'b11011:
        casez_tmp_61 = rob_uop_2_27_uses_stq;
      5'b11100:
        casez_tmp_61 = rob_uop_2_28_uses_stq;
      5'b11101:
        casez_tmp_61 = rob_uop_2_29_uses_stq;
      5'b11110:
        casez_tmp_61 = rob_uop_2_30_uses_stq;
      default:
        casez_tmp_61 = rob_uop_2_31_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_62 = rob_uop_2_0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_62 = rob_uop_2_1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_62 = rob_uop_2_2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_62 = rob_uop_2_3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_62 = rob_uop_2_4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_62 = rob_uop_2_5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_62 = rob_uop_2_6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_62 = rob_uop_2_7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_62 = rob_uop_2_8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_62 = rob_uop_2_9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_62 = rob_uop_2_10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_62 = rob_uop_2_11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_62 = rob_uop_2_12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_62 = rob_uop_2_13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_62 = rob_uop_2_14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_62 = rob_uop_2_15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_62 = rob_uop_2_16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_62 = rob_uop_2_17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_62 = rob_uop_2_18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_62 = rob_uop_2_19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_62 = rob_uop_2_20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_62 = rob_uop_2_21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_62 = rob_uop_2_22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_62 = rob_uop_2_23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_62 = rob_uop_2_24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_62 = rob_uop_2_25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_62 = rob_uop_2_26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_62 = rob_uop_2_27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_62 = rob_uop_2_28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_62 = rob_uop_2_29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_62 = rob_uop_2_30_is_sys_pc2epc;
      default:
        casez_tmp_62 = rob_uop_2_31_is_sys_pc2epc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_63 = rob_uop_2_0_flush_on_commit;
      5'b00001:
        casez_tmp_63 = rob_uop_2_1_flush_on_commit;
      5'b00010:
        casez_tmp_63 = rob_uop_2_2_flush_on_commit;
      5'b00011:
        casez_tmp_63 = rob_uop_2_3_flush_on_commit;
      5'b00100:
        casez_tmp_63 = rob_uop_2_4_flush_on_commit;
      5'b00101:
        casez_tmp_63 = rob_uop_2_5_flush_on_commit;
      5'b00110:
        casez_tmp_63 = rob_uop_2_6_flush_on_commit;
      5'b00111:
        casez_tmp_63 = rob_uop_2_7_flush_on_commit;
      5'b01000:
        casez_tmp_63 = rob_uop_2_8_flush_on_commit;
      5'b01001:
        casez_tmp_63 = rob_uop_2_9_flush_on_commit;
      5'b01010:
        casez_tmp_63 = rob_uop_2_10_flush_on_commit;
      5'b01011:
        casez_tmp_63 = rob_uop_2_11_flush_on_commit;
      5'b01100:
        casez_tmp_63 = rob_uop_2_12_flush_on_commit;
      5'b01101:
        casez_tmp_63 = rob_uop_2_13_flush_on_commit;
      5'b01110:
        casez_tmp_63 = rob_uop_2_14_flush_on_commit;
      5'b01111:
        casez_tmp_63 = rob_uop_2_15_flush_on_commit;
      5'b10000:
        casez_tmp_63 = rob_uop_2_16_flush_on_commit;
      5'b10001:
        casez_tmp_63 = rob_uop_2_17_flush_on_commit;
      5'b10010:
        casez_tmp_63 = rob_uop_2_18_flush_on_commit;
      5'b10011:
        casez_tmp_63 = rob_uop_2_19_flush_on_commit;
      5'b10100:
        casez_tmp_63 = rob_uop_2_20_flush_on_commit;
      5'b10101:
        casez_tmp_63 = rob_uop_2_21_flush_on_commit;
      5'b10110:
        casez_tmp_63 = rob_uop_2_22_flush_on_commit;
      5'b10111:
        casez_tmp_63 = rob_uop_2_23_flush_on_commit;
      5'b11000:
        casez_tmp_63 = rob_uop_2_24_flush_on_commit;
      5'b11001:
        casez_tmp_63 = rob_uop_2_25_flush_on_commit;
      5'b11010:
        casez_tmp_63 = rob_uop_2_26_flush_on_commit;
      5'b11011:
        casez_tmp_63 = rob_uop_2_27_flush_on_commit;
      5'b11100:
        casez_tmp_63 = rob_uop_2_28_flush_on_commit;
      5'b11101:
        casez_tmp_63 = rob_uop_2_29_flush_on_commit;
      5'b11110:
        casez_tmp_63 = rob_uop_2_30_flush_on_commit;
      default:
        casez_tmp_63 = rob_uop_2_31_flush_on_commit;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_64 = rob_uop_2_0_ldst;
      5'b00001:
        casez_tmp_64 = rob_uop_2_1_ldst;
      5'b00010:
        casez_tmp_64 = rob_uop_2_2_ldst;
      5'b00011:
        casez_tmp_64 = rob_uop_2_3_ldst;
      5'b00100:
        casez_tmp_64 = rob_uop_2_4_ldst;
      5'b00101:
        casez_tmp_64 = rob_uop_2_5_ldst;
      5'b00110:
        casez_tmp_64 = rob_uop_2_6_ldst;
      5'b00111:
        casez_tmp_64 = rob_uop_2_7_ldst;
      5'b01000:
        casez_tmp_64 = rob_uop_2_8_ldst;
      5'b01001:
        casez_tmp_64 = rob_uop_2_9_ldst;
      5'b01010:
        casez_tmp_64 = rob_uop_2_10_ldst;
      5'b01011:
        casez_tmp_64 = rob_uop_2_11_ldst;
      5'b01100:
        casez_tmp_64 = rob_uop_2_12_ldst;
      5'b01101:
        casez_tmp_64 = rob_uop_2_13_ldst;
      5'b01110:
        casez_tmp_64 = rob_uop_2_14_ldst;
      5'b01111:
        casez_tmp_64 = rob_uop_2_15_ldst;
      5'b10000:
        casez_tmp_64 = rob_uop_2_16_ldst;
      5'b10001:
        casez_tmp_64 = rob_uop_2_17_ldst;
      5'b10010:
        casez_tmp_64 = rob_uop_2_18_ldst;
      5'b10011:
        casez_tmp_64 = rob_uop_2_19_ldst;
      5'b10100:
        casez_tmp_64 = rob_uop_2_20_ldst;
      5'b10101:
        casez_tmp_64 = rob_uop_2_21_ldst;
      5'b10110:
        casez_tmp_64 = rob_uop_2_22_ldst;
      5'b10111:
        casez_tmp_64 = rob_uop_2_23_ldst;
      5'b11000:
        casez_tmp_64 = rob_uop_2_24_ldst;
      5'b11001:
        casez_tmp_64 = rob_uop_2_25_ldst;
      5'b11010:
        casez_tmp_64 = rob_uop_2_26_ldst;
      5'b11011:
        casez_tmp_64 = rob_uop_2_27_ldst;
      5'b11100:
        casez_tmp_64 = rob_uop_2_28_ldst;
      5'b11101:
        casez_tmp_64 = rob_uop_2_29_ldst;
      5'b11110:
        casez_tmp_64 = rob_uop_2_30_ldst;
      default:
        casez_tmp_64 = rob_uop_2_31_ldst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_65 = rob_uop_2_0_ldst_val;
      5'b00001:
        casez_tmp_65 = rob_uop_2_1_ldst_val;
      5'b00010:
        casez_tmp_65 = rob_uop_2_2_ldst_val;
      5'b00011:
        casez_tmp_65 = rob_uop_2_3_ldst_val;
      5'b00100:
        casez_tmp_65 = rob_uop_2_4_ldst_val;
      5'b00101:
        casez_tmp_65 = rob_uop_2_5_ldst_val;
      5'b00110:
        casez_tmp_65 = rob_uop_2_6_ldst_val;
      5'b00111:
        casez_tmp_65 = rob_uop_2_7_ldst_val;
      5'b01000:
        casez_tmp_65 = rob_uop_2_8_ldst_val;
      5'b01001:
        casez_tmp_65 = rob_uop_2_9_ldst_val;
      5'b01010:
        casez_tmp_65 = rob_uop_2_10_ldst_val;
      5'b01011:
        casez_tmp_65 = rob_uop_2_11_ldst_val;
      5'b01100:
        casez_tmp_65 = rob_uop_2_12_ldst_val;
      5'b01101:
        casez_tmp_65 = rob_uop_2_13_ldst_val;
      5'b01110:
        casez_tmp_65 = rob_uop_2_14_ldst_val;
      5'b01111:
        casez_tmp_65 = rob_uop_2_15_ldst_val;
      5'b10000:
        casez_tmp_65 = rob_uop_2_16_ldst_val;
      5'b10001:
        casez_tmp_65 = rob_uop_2_17_ldst_val;
      5'b10010:
        casez_tmp_65 = rob_uop_2_18_ldst_val;
      5'b10011:
        casez_tmp_65 = rob_uop_2_19_ldst_val;
      5'b10100:
        casez_tmp_65 = rob_uop_2_20_ldst_val;
      5'b10101:
        casez_tmp_65 = rob_uop_2_21_ldst_val;
      5'b10110:
        casez_tmp_65 = rob_uop_2_22_ldst_val;
      5'b10111:
        casez_tmp_65 = rob_uop_2_23_ldst_val;
      5'b11000:
        casez_tmp_65 = rob_uop_2_24_ldst_val;
      5'b11001:
        casez_tmp_65 = rob_uop_2_25_ldst_val;
      5'b11010:
        casez_tmp_65 = rob_uop_2_26_ldst_val;
      5'b11011:
        casez_tmp_65 = rob_uop_2_27_ldst_val;
      5'b11100:
        casez_tmp_65 = rob_uop_2_28_ldst_val;
      5'b11101:
        casez_tmp_65 = rob_uop_2_29_ldst_val;
      5'b11110:
        casez_tmp_65 = rob_uop_2_30_ldst_val;
      default:
        casez_tmp_65 = rob_uop_2_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_66 = rob_uop_2_0_dst_rtype;
      5'b00001:
        casez_tmp_66 = rob_uop_2_1_dst_rtype;
      5'b00010:
        casez_tmp_66 = rob_uop_2_2_dst_rtype;
      5'b00011:
        casez_tmp_66 = rob_uop_2_3_dst_rtype;
      5'b00100:
        casez_tmp_66 = rob_uop_2_4_dst_rtype;
      5'b00101:
        casez_tmp_66 = rob_uop_2_5_dst_rtype;
      5'b00110:
        casez_tmp_66 = rob_uop_2_6_dst_rtype;
      5'b00111:
        casez_tmp_66 = rob_uop_2_7_dst_rtype;
      5'b01000:
        casez_tmp_66 = rob_uop_2_8_dst_rtype;
      5'b01001:
        casez_tmp_66 = rob_uop_2_9_dst_rtype;
      5'b01010:
        casez_tmp_66 = rob_uop_2_10_dst_rtype;
      5'b01011:
        casez_tmp_66 = rob_uop_2_11_dst_rtype;
      5'b01100:
        casez_tmp_66 = rob_uop_2_12_dst_rtype;
      5'b01101:
        casez_tmp_66 = rob_uop_2_13_dst_rtype;
      5'b01110:
        casez_tmp_66 = rob_uop_2_14_dst_rtype;
      5'b01111:
        casez_tmp_66 = rob_uop_2_15_dst_rtype;
      5'b10000:
        casez_tmp_66 = rob_uop_2_16_dst_rtype;
      5'b10001:
        casez_tmp_66 = rob_uop_2_17_dst_rtype;
      5'b10010:
        casez_tmp_66 = rob_uop_2_18_dst_rtype;
      5'b10011:
        casez_tmp_66 = rob_uop_2_19_dst_rtype;
      5'b10100:
        casez_tmp_66 = rob_uop_2_20_dst_rtype;
      5'b10101:
        casez_tmp_66 = rob_uop_2_21_dst_rtype;
      5'b10110:
        casez_tmp_66 = rob_uop_2_22_dst_rtype;
      5'b10111:
        casez_tmp_66 = rob_uop_2_23_dst_rtype;
      5'b11000:
        casez_tmp_66 = rob_uop_2_24_dst_rtype;
      5'b11001:
        casez_tmp_66 = rob_uop_2_25_dst_rtype;
      5'b11010:
        casez_tmp_66 = rob_uop_2_26_dst_rtype;
      5'b11011:
        casez_tmp_66 = rob_uop_2_27_dst_rtype;
      5'b11100:
        casez_tmp_66 = rob_uop_2_28_dst_rtype;
      5'b11101:
        casez_tmp_66 = rob_uop_2_29_dst_rtype;
      5'b11110:
        casez_tmp_66 = rob_uop_2_30_dst_rtype;
      default:
        casez_tmp_66 = rob_uop_2_31_dst_rtype;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_67 = rob_uop_2_0_fp_val;
      5'b00001:
        casez_tmp_67 = rob_uop_2_1_fp_val;
      5'b00010:
        casez_tmp_67 = rob_uop_2_2_fp_val;
      5'b00011:
        casez_tmp_67 = rob_uop_2_3_fp_val;
      5'b00100:
        casez_tmp_67 = rob_uop_2_4_fp_val;
      5'b00101:
        casez_tmp_67 = rob_uop_2_5_fp_val;
      5'b00110:
        casez_tmp_67 = rob_uop_2_6_fp_val;
      5'b00111:
        casez_tmp_67 = rob_uop_2_7_fp_val;
      5'b01000:
        casez_tmp_67 = rob_uop_2_8_fp_val;
      5'b01001:
        casez_tmp_67 = rob_uop_2_9_fp_val;
      5'b01010:
        casez_tmp_67 = rob_uop_2_10_fp_val;
      5'b01011:
        casez_tmp_67 = rob_uop_2_11_fp_val;
      5'b01100:
        casez_tmp_67 = rob_uop_2_12_fp_val;
      5'b01101:
        casez_tmp_67 = rob_uop_2_13_fp_val;
      5'b01110:
        casez_tmp_67 = rob_uop_2_14_fp_val;
      5'b01111:
        casez_tmp_67 = rob_uop_2_15_fp_val;
      5'b10000:
        casez_tmp_67 = rob_uop_2_16_fp_val;
      5'b10001:
        casez_tmp_67 = rob_uop_2_17_fp_val;
      5'b10010:
        casez_tmp_67 = rob_uop_2_18_fp_val;
      5'b10011:
        casez_tmp_67 = rob_uop_2_19_fp_val;
      5'b10100:
        casez_tmp_67 = rob_uop_2_20_fp_val;
      5'b10101:
        casez_tmp_67 = rob_uop_2_21_fp_val;
      5'b10110:
        casez_tmp_67 = rob_uop_2_22_fp_val;
      5'b10111:
        casez_tmp_67 = rob_uop_2_23_fp_val;
      5'b11000:
        casez_tmp_67 = rob_uop_2_24_fp_val;
      5'b11001:
        casez_tmp_67 = rob_uop_2_25_fp_val;
      5'b11010:
        casez_tmp_67 = rob_uop_2_26_fp_val;
      5'b11011:
        casez_tmp_67 = rob_uop_2_27_fp_val;
      5'b11100:
        casez_tmp_67 = rob_uop_2_28_fp_val;
      5'b11101:
        casez_tmp_67 = rob_uop_2_29_fp_val;
      5'b11110:
        casez_tmp_67 = rob_uop_2_30_fp_val;
      default:
        casez_tmp_67 = rob_uop_2_31_fp_val;
    endcase
  end // always @(*)
  wire        rbk_row_2 = _io_commit_rollback_T_3 & ~full;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_68 = rob_val_2_0;
      5'b00001:
        casez_tmp_68 = rob_val_2_1;
      5'b00010:
        casez_tmp_68 = rob_val_2_2;
      5'b00011:
        casez_tmp_68 = rob_val_2_3;
      5'b00100:
        casez_tmp_68 = rob_val_2_4;
      5'b00101:
        casez_tmp_68 = rob_val_2_5;
      5'b00110:
        casez_tmp_68 = rob_val_2_6;
      5'b00111:
        casez_tmp_68 = rob_val_2_7;
      5'b01000:
        casez_tmp_68 = rob_val_2_8;
      5'b01001:
        casez_tmp_68 = rob_val_2_9;
      5'b01010:
        casez_tmp_68 = rob_val_2_10;
      5'b01011:
        casez_tmp_68 = rob_val_2_11;
      5'b01100:
        casez_tmp_68 = rob_val_2_12;
      5'b01101:
        casez_tmp_68 = rob_val_2_13;
      5'b01110:
        casez_tmp_68 = rob_val_2_14;
      5'b01111:
        casez_tmp_68 = rob_val_2_15;
      5'b10000:
        casez_tmp_68 = rob_val_2_16;
      5'b10001:
        casez_tmp_68 = rob_val_2_17;
      5'b10010:
        casez_tmp_68 = rob_val_2_18;
      5'b10011:
        casez_tmp_68 = rob_val_2_19;
      5'b10100:
        casez_tmp_68 = rob_val_2_20;
      5'b10101:
        casez_tmp_68 = rob_val_2_21;
      5'b10110:
        casez_tmp_68 = rob_val_2_22;
      5'b10111:
        casez_tmp_68 = rob_val_2_23;
      5'b11000:
        casez_tmp_68 = rob_val_2_24;
      5'b11001:
        casez_tmp_68 = rob_val_2_25;
      5'b11010:
        casez_tmp_68 = rob_val_2_26;
      5'b11011:
        casez_tmp_68 = rob_val_2_27;
      5'b11100:
        casez_tmp_68 = rob_val_2_28;
      5'b11101:
        casez_tmp_68 = rob_val_2_29;
      5'b11110:
        casez_tmp_68 = rob_val_2_30;
      default:
        casez_tmp_68 = rob_val_2_31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_2_output = rbk_row_2 & casez_tmp_68;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_69 = rob_fflags_2_0;
      5'b00001:
        casez_tmp_69 = rob_fflags_2_1;
      5'b00010:
        casez_tmp_69 = rob_fflags_2_2;
      5'b00011:
        casez_tmp_69 = rob_fflags_2_3;
      5'b00100:
        casez_tmp_69 = rob_fflags_2_4;
      5'b00101:
        casez_tmp_69 = rob_fflags_2_5;
      5'b00110:
        casez_tmp_69 = rob_fflags_2_6;
      5'b00111:
        casez_tmp_69 = rob_fflags_2_7;
      5'b01000:
        casez_tmp_69 = rob_fflags_2_8;
      5'b01001:
        casez_tmp_69 = rob_fflags_2_9;
      5'b01010:
        casez_tmp_69 = rob_fflags_2_10;
      5'b01011:
        casez_tmp_69 = rob_fflags_2_11;
      5'b01100:
        casez_tmp_69 = rob_fflags_2_12;
      5'b01101:
        casez_tmp_69 = rob_fflags_2_13;
      5'b01110:
        casez_tmp_69 = rob_fflags_2_14;
      5'b01111:
        casez_tmp_69 = rob_fflags_2_15;
      5'b10000:
        casez_tmp_69 = rob_fflags_2_16;
      5'b10001:
        casez_tmp_69 = rob_fflags_2_17;
      5'b10010:
        casez_tmp_69 = rob_fflags_2_18;
      5'b10011:
        casez_tmp_69 = rob_fflags_2_19;
      5'b10100:
        casez_tmp_69 = rob_fflags_2_20;
      5'b10101:
        casez_tmp_69 = rob_fflags_2_21;
      5'b10110:
        casez_tmp_69 = rob_fflags_2_22;
      5'b10111:
        casez_tmp_69 = rob_fflags_2_23;
      5'b11000:
        casez_tmp_69 = rob_fflags_2_24;
      5'b11001:
        casez_tmp_69 = rob_fflags_2_25;
      5'b11010:
        casez_tmp_69 = rob_fflags_2_26;
      5'b11011:
        casez_tmp_69 = rob_fflags_2_27;
      5'b11100:
        casez_tmp_69 = rob_fflags_2_28;
      5'b11101:
        casez_tmp_69 = rob_fflags_2_29;
      5'b11110:
        casez_tmp_69 = rob_fflags_2_30;
      default:
        casez_tmp_69 = rob_fflags_2_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_70 = rob_uop_2_0_uses_ldq;
      5'b00001:
        casez_tmp_70 = rob_uop_2_1_uses_ldq;
      5'b00010:
        casez_tmp_70 = rob_uop_2_2_uses_ldq;
      5'b00011:
        casez_tmp_70 = rob_uop_2_3_uses_ldq;
      5'b00100:
        casez_tmp_70 = rob_uop_2_4_uses_ldq;
      5'b00101:
        casez_tmp_70 = rob_uop_2_5_uses_ldq;
      5'b00110:
        casez_tmp_70 = rob_uop_2_6_uses_ldq;
      5'b00111:
        casez_tmp_70 = rob_uop_2_7_uses_ldq;
      5'b01000:
        casez_tmp_70 = rob_uop_2_8_uses_ldq;
      5'b01001:
        casez_tmp_70 = rob_uop_2_9_uses_ldq;
      5'b01010:
        casez_tmp_70 = rob_uop_2_10_uses_ldq;
      5'b01011:
        casez_tmp_70 = rob_uop_2_11_uses_ldq;
      5'b01100:
        casez_tmp_70 = rob_uop_2_12_uses_ldq;
      5'b01101:
        casez_tmp_70 = rob_uop_2_13_uses_ldq;
      5'b01110:
        casez_tmp_70 = rob_uop_2_14_uses_ldq;
      5'b01111:
        casez_tmp_70 = rob_uop_2_15_uses_ldq;
      5'b10000:
        casez_tmp_70 = rob_uop_2_16_uses_ldq;
      5'b10001:
        casez_tmp_70 = rob_uop_2_17_uses_ldq;
      5'b10010:
        casez_tmp_70 = rob_uop_2_18_uses_ldq;
      5'b10011:
        casez_tmp_70 = rob_uop_2_19_uses_ldq;
      5'b10100:
        casez_tmp_70 = rob_uop_2_20_uses_ldq;
      5'b10101:
        casez_tmp_70 = rob_uop_2_21_uses_ldq;
      5'b10110:
        casez_tmp_70 = rob_uop_2_22_uses_ldq;
      5'b10111:
        casez_tmp_70 = rob_uop_2_23_uses_ldq;
      5'b11000:
        casez_tmp_70 = rob_uop_2_24_uses_ldq;
      5'b11001:
        casez_tmp_70 = rob_uop_2_25_uses_ldq;
      5'b11010:
        casez_tmp_70 = rob_uop_2_26_uses_ldq;
      5'b11011:
        casez_tmp_70 = rob_uop_2_27_uses_ldq;
      5'b11100:
        casez_tmp_70 = rob_uop_2_28_uses_ldq;
      5'b11101:
        casez_tmp_70 = rob_uop_2_29_uses_ldq;
      5'b11110:
        casez_tmp_70 = rob_uop_2_30_uses_ldq;
      default:
        casez_tmp_70 = rob_uop_2_31_uses_ldq;
    endcase
  end // always @(*)
  reg  [6:0]  rob_uop_3_0_uopc;
  reg         rob_uop_3_0_is_rvc;
  reg  [19:0] rob_uop_3_0_br_mask;
  reg  [5:0]  rob_uop_3_0_ftq_idx;
  reg         rob_uop_3_0_edge_inst;
  reg  [5:0]  rob_uop_3_0_pc_lob;
  reg  [6:0]  rob_uop_3_0_pdst;
  reg  [6:0]  rob_uop_3_0_stale_pdst;
  reg         rob_uop_3_0_is_fencei;
  reg         rob_uop_3_0_uses_ldq;
  reg         rob_uop_3_0_uses_stq;
  reg         rob_uop_3_0_is_sys_pc2epc;
  reg         rob_uop_3_0_flush_on_commit;
  reg  [5:0]  rob_uop_3_0_ldst;
  reg         rob_uop_3_0_ldst_val;
  reg  [1:0]  rob_uop_3_0_dst_rtype;
  reg         rob_uop_3_0_fp_val;
  reg  [6:0]  rob_uop_3_1_uopc;
  reg         rob_uop_3_1_is_rvc;
  reg  [19:0] rob_uop_3_1_br_mask;
  reg  [5:0]  rob_uop_3_1_ftq_idx;
  reg         rob_uop_3_1_edge_inst;
  reg  [5:0]  rob_uop_3_1_pc_lob;
  reg  [6:0]  rob_uop_3_1_pdst;
  reg  [6:0]  rob_uop_3_1_stale_pdst;
  reg         rob_uop_3_1_is_fencei;
  reg         rob_uop_3_1_uses_ldq;
  reg         rob_uop_3_1_uses_stq;
  reg         rob_uop_3_1_is_sys_pc2epc;
  reg         rob_uop_3_1_flush_on_commit;
  reg  [5:0]  rob_uop_3_1_ldst;
  reg         rob_uop_3_1_ldst_val;
  reg  [1:0]  rob_uop_3_1_dst_rtype;
  reg         rob_uop_3_1_fp_val;
  reg  [6:0]  rob_uop_3_2_uopc;
  reg         rob_uop_3_2_is_rvc;
  reg  [19:0] rob_uop_3_2_br_mask;
  reg  [5:0]  rob_uop_3_2_ftq_idx;
  reg         rob_uop_3_2_edge_inst;
  reg  [5:0]  rob_uop_3_2_pc_lob;
  reg  [6:0]  rob_uop_3_2_pdst;
  reg  [6:0]  rob_uop_3_2_stale_pdst;
  reg         rob_uop_3_2_is_fencei;
  reg         rob_uop_3_2_uses_ldq;
  reg         rob_uop_3_2_uses_stq;
  reg         rob_uop_3_2_is_sys_pc2epc;
  reg         rob_uop_3_2_flush_on_commit;
  reg  [5:0]  rob_uop_3_2_ldst;
  reg         rob_uop_3_2_ldst_val;
  reg  [1:0]  rob_uop_3_2_dst_rtype;
  reg         rob_uop_3_2_fp_val;
  reg  [6:0]  rob_uop_3_3_uopc;
  reg         rob_uop_3_3_is_rvc;
  reg  [19:0] rob_uop_3_3_br_mask;
  reg  [5:0]  rob_uop_3_3_ftq_idx;
  reg         rob_uop_3_3_edge_inst;
  reg  [5:0]  rob_uop_3_3_pc_lob;
  reg  [6:0]  rob_uop_3_3_pdst;
  reg  [6:0]  rob_uop_3_3_stale_pdst;
  reg         rob_uop_3_3_is_fencei;
  reg         rob_uop_3_3_uses_ldq;
  reg         rob_uop_3_3_uses_stq;
  reg         rob_uop_3_3_is_sys_pc2epc;
  reg         rob_uop_3_3_flush_on_commit;
  reg  [5:0]  rob_uop_3_3_ldst;
  reg         rob_uop_3_3_ldst_val;
  reg  [1:0]  rob_uop_3_3_dst_rtype;
  reg         rob_uop_3_3_fp_val;
  reg  [6:0]  rob_uop_3_4_uopc;
  reg         rob_uop_3_4_is_rvc;
  reg  [19:0] rob_uop_3_4_br_mask;
  reg  [5:0]  rob_uop_3_4_ftq_idx;
  reg         rob_uop_3_4_edge_inst;
  reg  [5:0]  rob_uop_3_4_pc_lob;
  reg  [6:0]  rob_uop_3_4_pdst;
  reg  [6:0]  rob_uop_3_4_stale_pdst;
  reg         rob_uop_3_4_is_fencei;
  reg         rob_uop_3_4_uses_ldq;
  reg         rob_uop_3_4_uses_stq;
  reg         rob_uop_3_4_is_sys_pc2epc;
  reg         rob_uop_3_4_flush_on_commit;
  reg  [5:0]  rob_uop_3_4_ldst;
  reg         rob_uop_3_4_ldst_val;
  reg  [1:0]  rob_uop_3_4_dst_rtype;
  reg         rob_uop_3_4_fp_val;
  reg  [6:0]  rob_uop_3_5_uopc;
  reg         rob_uop_3_5_is_rvc;
  reg  [19:0] rob_uop_3_5_br_mask;
  reg  [5:0]  rob_uop_3_5_ftq_idx;
  reg         rob_uop_3_5_edge_inst;
  reg  [5:0]  rob_uop_3_5_pc_lob;
  reg  [6:0]  rob_uop_3_5_pdst;
  reg  [6:0]  rob_uop_3_5_stale_pdst;
  reg         rob_uop_3_5_is_fencei;
  reg         rob_uop_3_5_uses_ldq;
  reg         rob_uop_3_5_uses_stq;
  reg         rob_uop_3_5_is_sys_pc2epc;
  reg         rob_uop_3_5_flush_on_commit;
  reg  [5:0]  rob_uop_3_5_ldst;
  reg         rob_uop_3_5_ldst_val;
  reg  [1:0]  rob_uop_3_5_dst_rtype;
  reg         rob_uop_3_5_fp_val;
  reg  [6:0]  rob_uop_3_6_uopc;
  reg         rob_uop_3_6_is_rvc;
  reg  [19:0] rob_uop_3_6_br_mask;
  reg  [5:0]  rob_uop_3_6_ftq_idx;
  reg         rob_uop_3_6_edge_inst;
  reg  [5:0]  rob_uop_3_6_pc_lob;
  reg  [6:0]  rob_uop_3_6_pdst;
  reg  [6:0]  rob_uop_3_6_stale_pdst;
  reg         rob_uop_3_6_is_fencei;
  reg         rob_uop_3_6_uses_ldq;
  reg         rob_uop_3_6_uses_stq;
  reg         rob_uop_3_6_is_sys_pc2epc;
  reg         rob_uop_3_6_flush_on_commit;
  reg  [5:0]  rob_uop_3_6_ldst;
  reg         rob_uop_3_6_ldst_val;
  reg  [1:0]  rob_uop_3_6_dst_rtype;
  reg         rob_uop_3_6_fp_val;
  reg  [6:0]  rob_uop_3_7_uopc;
  reg         rob_uop_3_7_is_rvc;
  reg  [19:0] rob_uop_3_7_br_mask;
  reg  [5:0]  rob_uop_3_7_ftq_idx;
  reg         rob_uop_3_7_edge_inst;
  reg  [5:0]  rob_uop_3_7_pc_lob;
  reg  [6:0]  rob_uop_3_7_pdst;
  reg  [6:0]  rob_uop_3_7_stale_pdst;
  reg         rob_uop_3_7_is_fencei;
  reg         rob_uop_3_7_uses_ldq;
  reg         rob_uop_3_7_uses_stq;
  reg         rob_uop_3_7_is_sys_pc2epc;
  reg         rob_uop_3_7_flush_on_commit;
  reg  [5:0]  rob_uop_3_7_ldst;
  reg         rob_uop_3_7_ldst_val;
  reg  [1:0]  rob_uop_3_7_dst_rtype;
  reg         rob_uop_3_7_fp_val;
  reg  [6:0]  rob_uop_3_8_uopc;
  reg         rob_uop_3_8_is_rvc;
  reg  [19:0] rob_uop_3_8_br_mask;
  reg  [5:0]  rob_uop_3_8_ftq_idx;
  reg         rob_uop_3_8_edge_inst;
  reg  [5:0]  rob_uop_3_8_pc_lob;
  reg  [6:0]  rob_uop_3_8_pdst;
  reg  [6:0]  rob_uop_3_8_stale_pdst;
  reg         rob_uop_3_8_is_fencei;
  reg         rob_uop_3_8_uses_ldq;
  reg         rob_uop_3_8_uses_stq;
  reg         rob_uop_3_8_is_sys_pc2epc;
  reg         rob_uop_3_8_flush_on_commit;
  reg  [5:0]  rob_uop_3_8_ldst;
  reg         rob_uop_3_8_ldst_val;
  reg  [1:0]  rob_uop_3_8_dst_rtype;
  reg         rob_uop_3_8_fp_val;
  reg  [6:0]  rob_uop_3_9_uopc;
  reg         rob_uop_3_9_is_rvc;
  reg  [19:0] rob_uop_3_9_br_mask;
  reg  [5:0]  rob_uop_3_9_ftq_idx;
  reg         rob_uop_3_9_edge_inst;
  reg  [5:0]  rob_uop_3_9_pc_lob;
  reg  [6:0]  rob_uop_3_9_pdst;
  reg  [6:0]  rob_uop_3_9_stale_pdst;
  reg         rob_uop_3_9_is_fencei;
  reg         rob_uop_3_9_uses_ldq;
  reg         rob_uop_3_9_uses_stq;
  reg         rob_uop_3_9_is_sys_pc2epc;
  reg         rob_uop_3_9_flush_on_commit;
  reg  [5:0]  rob_uop_3_9_ldst;
  reg         rob_uop_3_9_ldst_val;
  reg  [1:0]  rob_uop_3_9_dst_rtype;
  reg         rob_uop_3_9_fp_val;
  reg  [6:0]  rob_uop_3_10_uopc;
  reg         rob_uop_3_10_is_rvc;
  reg  [19:0] rob_uop_3_10_br_mask;
  reg  [5:0]  rob_uop_3_10_ftq_idx;
  reg         rob_uop_3_10_edge_inst;
  reg  [5:0]  rob_uop_3_10_pc_lob;
  reg  [6:0]  rob_uop_3_10_pdst;
  reg  [6:0]  rob_uop_3_10_stale_pdst;
  reg         rob_uop_3_10_is_fencei;
  reg         rob_uop_3_10_uses_ldq;
  reg         rob_uop_3_10_uses_stq;
  reg         rob_uop_3_10_is_sys_pc2epc;
  reg         rob_uop_3_10_flush_on_commit;
  reg  [5:0]  rob_uop_3_10_ldst;
  reg         rob_uop_3_10_ldst_val;
  reg  [1:0]  rob_uop_3_10_dst_rtype;
  reg         rob_uop_3_10_fp_val;
  reg  [6:0]  rob_uop_3_11_uopc;
  reg         rob_uop_3_11_is_rvc;
  reg  [19:0] rob_uop_3_11_br_mask;
  reg  [5:0]  rob_uop_3_11_ftq_idx;
  reg         rob_uop_3_11_edge_inst;
  reg  [5:0]  rob_uop_3_11_pc_lob;
  reg  [6:0]  rob_uop_3_11_pdst;
  reg  [6:0]  rob_uop_3_11_stale_pdst;
  reg         rob_uop_3_11_is_fencei;
  reg         rob_uop_3_11_uses_ldq;
  reg         rob_uop_3_11_uses_stq;
  reg         rob_uop_3_11_is_sys_pc2epc;
  reg         rob_uop_3_11_flush_on_commit;
  reg  [5:0]  rob_uop_3_11_ldst;
  reg         rob_uop_3_11_ldst_val;
  reg  [1:0]  rob_uop_3_11_dst_rtype;
  reg         rob_uop_3_11_fp_val;
  reg  [6:0]  rob_uop_3_12_uopc;
  reg         rob_uop_3_12_is_rvc;
  reg  [19:0] rob_uop_3_12_br_mask;
  reg  [5:0]  rob_uop_3_12_ftq_idx;
  reg         rob_uop_3_12_edge_inst;
  reg  [5:0]  rob_uop_3_12_pc_lob;
  reg  [6:0]  rob_uop_3_12_pdst;
  reg  [6:0]  rob_uop_3_12_stale_pdst;
  reg         rob_uop_3_12_is_fencei;
  reg         rob_uop_3_12_uses_ldq;
  reg         rob_uop_3_12_uses_stq;
  reg         rob_uop_3_12_is_sys_pc2epc;
  reg         rob_uop_3_12_flush_on_commit;
  reg  [5:0]  rob_uop_3_12_ldst;
  reg         rob_uop_3_12_ldst_val;
  reg  [1:0]  rob_uop_3_12_dst_rtype;
  reg         rob_uop_3_12_fp_val;
  reg  [6:0]  rob_uop_3_13_uopc;
  reg         rob_uop_3_13_is_rvc;
  reg  [19:0] rob_uop_3_13_br_mask;
  reg  [5:0]  rob_uop_3_13_ftq_idx;
  reg         rob_uop_3_13_edge_inst;
  reg  [5:0]  rob_uop_3_13_pc_lob;
  reg  [6:0]  rob_uop_3_13_pdst;
  reg  [6:0]  rob_uop_3_13_stale_pdst;
  reg         rob_uop_3_13_is_fencei;
  reg         rob_uop_3_13_uses_ldq;
  reg         rob_uop_3_13_uses_stq;
  reg         rob_uop_3_13_is_sys_pc2epc;
  reg         rob_uop_3_13_flush_on_commit;
  reg  [5:0]  rob_uop_3_13_ldst;
  reg         rob_uop_3_13_ldst_val;
  reg  [1:0]  rob_uop_3_13_dst_rtype;
  reg         rob_uop_3_13_fp_val;
  reg  [6:0]  rob_uop_3_14_uopc;
  reg         rob_uop_3_14_is_rvc;
  reg  [19:0] rob_uop_3_14_br_mask;
  reg  [5:0]  rob_uop_3_14_ftq_idx;
  reg         rob_uop_3_14_edge_inst;
  reg  [5:0]  rob_uop_3_14_pc_lob;
  reg  [6:0]  rob_uop_3_14_pdst;
  reg  [6:0]  rob_uop_3_14_stale_pdst;
  reg         rob_uop_3_14_is_fencei;
  reg         rob_uop_3_14_uses_ldq;
  reg         rob_uop_3_14_uses_stq;
  reg         rob_uop_3_14_is_sys_pc2epc;
  reg         rob_uop_3_14_flush_on_commit;
  reg  [5:0]  rob_uop_3_14_ldst;
  reg         rob_uop_3_14_ldst_val;
  reg  [1:0]  rob_uop_3_14_dst_rtype;
  reg         rob_uop_3_14_fp_val;
  reg  [6:0]  rob_uop_3_15_uopc;
  reg         rob_uop_3_15_is_rvc;
  reg  [19:0] rob_uop_3_15_br_mask;
  reg  [5:0]  rob_uop_3_15_ftq_idx;
  reg         rob_uop_3_15_edge_inst;
  reg  [5:0]  rob_uop_3_15_pc_lob;
  reg  [6:0]  rob_uop_3_15_pdst;
  reg  [6:0]  rob_uop_3_15_stale_pdst;
  reg         rob_uop_3_15_is_fencei;
  reg         rob_uop_3_15_uses_ldq;
  reg         rob_uop_3_15_uses_stq;
  reg         rob_uop_3_15_is_sys_pc2epc;
  reg         rob_uop_3_15_flush_on_commit;
  reg  [5:0]  rob_uop_3_15_ldst;
  reg         rob_uop_3_15_ldst_val;
  reg  [1:0]  rob_uop_3_15_dst_rtype;
  reg         rob_uop_3_15_fp_val;
  reg  [6:0]  rob_uop_3_16_uopc;
  reg         rob_uop_3_16_is_rvc;
  reg  [19:0] rob_uop_3_16_br_mask;
  reg  [5:0]  rob_uop_3_16_ftq_idx;
  reg         rob_uop_3_16_edge_inst;
  reg  [5:0]  rob_uop_3_16_pc_lob;
  reg  [6:0]  rob_uop_3_16_pdst;
  reg  [6:0]  rob_uop_3_16_stale_pdst;
  reg         rob_uop_3_16_is_fencei;
  reg         rob_uop_3_16_uses_ldq;
  reg         rob_uop_3_16_uses_stq;
  reg         rob_uop_3_16_is_sys_pc2epc;
  reg         rob_uop_3_16_flush_on_commit;
  reg  [5:0]  rob_uop_3_16_ldst;
  reg         rob_uop_3_16_ldst_val;
  reg  [1:0]  rob_uop_3_16_dst_rtype;
  reg         rob_uop_3_16_fp_val;
  reg  [6:0]  rob_uop_3_17_uopc;
  reg         rob_uop_3_17_is_rvc;
  reg  [19:0] rob_uop_3_17_br_mask;
  reg  [5:0]  rob_uop_3_17_ftq_idx;
  reg         rob_uop_3_17_edge_inst;
  reg  [5:0]  rob_uop_3_17_pc_lob;
  reg  [6:0]  rob_uop_3_17_pdst;
  reg  [6:0]  rob_uop_3_17_stale_pdst;
  reg         rob_uop_3_17_is_fencei;
  reg         rob_uop_3_17_uses_ldq;
  reg         rob_uop_3_17_uses_stq;
  reg         rob_uop_3_17_is_sys_pc2epc;
  reg         rob_uop_3_17_flush_on_commit;
  reg  [5:0]  rob_uop_3_17_ldst;
  reg         rob_uop_3_17_ldst_val;
  reg  [1:0]  rob_uop_3_17_dst_rtype;
  reg         rob_uop_3_17_fp_val;
  reg  [6:0]  rob_uop_3_18_uopc;
  reg         rob_uop_3_18_is_rvc;
  reg  [19:0] rob_uop_3_18_br_mask;
  reg  [5:0]  rob_uop_3_18_ftq_idx;
  reg         rob_uop_3_18_edge_inst;
  reg  [5:0]  rob_uop_3_18_pc_lob;
  reg  [6:0]  rob_uop_3_18_pdst;
  reg  [6:0]  rob_uop_3_18_stale_pdst;
  reg         rob_uop_3_18_is_fencei;
  reg         rob_uop_3_18_uses_ldq;
  reg         rob_uop_3_18_uses_stq;
  reg         rob_uop_3_18_is_sys_pc2epc;
  reg         rob_uop_3_18_flush_on_commit;
  reg  [5:0]  rob_uop_3_18_ldst;
  reg         rob_uop_3_18_ldst_val;
  reg  [1:0]  rob_uop_3_18_dst_rtype;
  reg         rob_uop_3_18_fp_val;
  reg  [6:0]  rob_uop_3_19_uopc;
  reg         rob_uop_3_19_is_rvc;
  reg  [19:0] rob_uop_3_19_br_mask;
  reg  [5:0]  rob_uop_3_19_ftq_idx;
  reg         rob_uop_3_19_edge_inst;
  reg  [5:0]  rob_uop_3_19_pc_lob;
  reg  [6:0]  rob_uop_3_19_pdst;
  reg  [6:0]  rob_uop_3_19_stale_pdst;
  reg         rob_uop_3_19_is_fencei;
  reg         rob_uop_3_19_uses_ldq;
  reg         rob_uop_3_19_uses_stq;
  reg         rob_uop_3_19_is_sys_pc2epc;
  reg         rob_uop_3_19_flush_on_commit;
  reg  [5:0]  rob_uop_3_19_ldst;
  reg         rob_uop_3_19_ldst_val;
  reg  [1:0]  rob_uop_3_19_dst_rtype;
  reg         rob_uop_3_19_fp_val;
  reg  [6:0]  rob_uop_3_20_uopc;
  reg         rob_uop_3_20_is_rvc;
  reg  [19:0] rob_uop_3_20_br_mask;
  reg  [5:0]  rob_uop_3_20_ftq_idx;
  reg         rob_uop_3_20_edge_inst;
  reg  [5:0]  rob_uop_3_20_pc_lob;
  reg  [6:0]  rob_uop_3_20_pdst;
  reg  [6:0]  rob_uop_3_20_stale_pdst;
  reg         rob_uop_3_20_is_fencei;
  reg         rob_uop_3_20_uses_ldq;
  reg         rob_uop_3_20_uses_stq;
  reg         rob_uop_3_20_is_sys_pc2epc;
  reg         rob_uop_3_20_flush_on_commit;
  reg  [5:0]  rob_uop_3_20_ldst;
  reg         rob_uop_3_20_ldst_val;
  reg  [1:0]  rob_uop_3_20_dst_rtype;
  reg         rob_uop_3_20_fp_val;
  reg  [6:0]  rob_uop_3_21_uopc;
  reg         rob_uop_3_21_is_rvc;
  reg  [19:0] rob_uop_3_21_br_mask;
  reg  [5:0]  rob_uop_3_21_ftq_idx;
  reg         rob_uop_3_21_edge_inst;
  reg  [5:0]  rob_uop_3_21_pc_lob;
  reg  [6:0]  rob_uop_3_21_pdst;
  reg  [6:0]  rob_uop_3_21_stale_pdst;
  reg         rob_uop_3_21_is_fencei;
  reg         rob_uop_3_21_uses_ldq;
  reg         rob_uop_3_21_uses_stq;
  reg         rob_uop_3_21_is_sys_pc2epc;
  reg         rob_uop_3_21_flush_on_commit;
  reg  [5:0]  rob_uop_3_21_ldst;
  reg         rob_uop_3_21_ldst_val;
  reg  [1:0]  rob_uop_3_21_dst_rtype;
  reg         rob_uop_3_21_fp_val;
  reg  [6:0]  rob_uop_3_22_uopc;
  reg         rob_uop_3_22_is_rvc;
  reg  [19:0] rob_uop_3_22_br_mask;
  reg  [5:0]  rob_uop_3_22_ftq_idx;
  reg         rob_uop_3_22_edge_inst;
  reg  [5:0]  rob_uop_3_22_pc_lob;
  reg  [6:0]  rob_uop_3_22_pdst;
  reg  [6:0]  rob_uop_3_22_stale_pdst;
  reg         rob_uop_3_22_is_fencei;
  reg         rob_uop_3_22_uses_ldq;
  reg         rob_uop_3_22_uses_stq;
  reg         rob_uop_3_22_is_sys_pc2epc;
  reg         rob_uop_3_22_flush_on_commit;
  reg  [5:0]  rob_uop_3_22_ldst;
  reg         rob_uop_3_22_ldst_val;
  reg  [1:0]  rob_uop_3_22_dst_rtype;
  reg         rob_uop_3_22_fp_val;
  reg  [6:0]  rob_uop_3_23_uopc;
  reg         rob_uop_3_23_is_rvc;
  reg  [19:0] rob_uop_3_23_br_mask;
  reg  [5:0]  rob_uop_3_23_ftq_idx;
  reg         rob_uop_3_23_edge_inst;
  reg  [5:0]  rob_uop_3_23_pc_lob;
  reg  [6:0]  rob_uop_3_23_pdst;
  reg  [6:0]  rob_uop_3_23_stale_pdst;
  reg         rob_uop_3_23_is_fencei;
  reg         rob_uop_3_23_uses_ldq;
  reg         rob_uop_3_23_uses_stq;
  reg         rob_uop_3_23_is_sys_pc2epc;
  reg         rob_uop_3_23_flush_on_commit;
  reg  [5:0]  rob_uop_3_23_ldst;
  reg         rob_uop_3_23_ldst_val;
  reg  [1:0]  rob_uop_3_23_dst_rtype;
  reg         rob_uop_3_23_fp_val;
  reg  [6:0]  rob_uop_3_24_uopc;
  reg         rob_uop_3_24_is_rvc;
  reg  [19:0] rob_uop_3_24_br_mask;
  reg  [5:0]  rob_uop_3_24_ftq_idx;
  reg         rob_uop_3_24_edge_inst;
  reg  [5:0]  rob_uop_3_24_pc_lob;
  reg  [6:0]  rob_uop_3_24_pdst;
  reg  [6:0]  rob_uop_3_24_stale_pdst;
  reg         rob_uop_3_24_is_fencei;
  reg         rob_uop_3_24_uses_ldq;
  reg         rob_uop_3_24_uses_stq;
  reg         rob_uop_3_24_is_sys_pc2epc;
  reg         rob_uop_3_24_flush_on_commit;
  reg  [5:0]  rob_uop_3_24_ldst;
  reg         rob_uop_3_24_ldst_val;
  reg  [1:0]  rob_uop_3_24_dst_rtype;
  reg         rob_uop_3_24_fp_val;
  reg  [6:0]  rob_uop_3_25_uopc;
  reg         rob_uop_3_25_is_rvc;
  reg  [19:0] rob_uop_3_25_br_mask;
  reg  [5:0]  rob_uop_3_25_ftq_idx;
  reg         rob_uop_3_25_edge_inst;
  reg  [5:0]  rob_uop_3_25_pc_lob;
  reg  [6:0]  rob_uop_3_25_pdst;
  reg  [6:0]  rob_uop_3_25_stale_pdst;
  reg         rob_uop_3_25_is_fencei;
  reg         rob_uop_3_25_uses_ldq;
  reg         rob_uop_3_25_uses_stq;
  reg         rob_uop_3_25_is_sys_pc2epc;
  reg         rob_uop_3_25_flush_on_commit;
  reg  [5:0]  rob_uop_3_25_ldst;
  reg         rob_uop_3_25_ldst_val;
  reg  [1:0]  rob_uop_3_25_dst_rtype;
  reg         rob_uop_3_25_fp_val;
  reg  [6:0]  rob_uop_3_26_uopc;
  reg         rob_uop_3_26_is_rvc;
  reg  [19:0] rob_uop_3_26_br_mask;
  reg  [5:0]  rob_uop_3_26_ftq_idx;
  reg         rob_uop_3_26_edge_inst;
  reg  [5:0]  rob_uop_3_26_pc_lob;
  reg  [6:0]  rob_uop_3_26_pdst;
  reg  [6:0]  rob_uop_3_26_stale_pdst;
  reg         rob_uop_3_26_is_fencei;
  reg         rob_uop_3_26_uses_ldq;
  reg         rob_uop_3_26_uses_stq;
  reg         rob_uop_3_26_is_sys_pc2epc;
  reg         rob_uop_3_26_flush_on_commit;
  reg  [5:0]  rob_uop_3_26_ldst;
  reg         rob_uop_3_26_ldst_val;
  reg  [1:0]  rob_uop_3_26_dst_rtype;
  reg         rob_uop_3_26_fp_val;
  reg  [6:0]  rob_uop_3_27_uopc;
  reg         rob_uop_3_27_is_rvc;
  reg  [19:0] rob_uop_3_27_br_mask;
  reg  [5:0]  rob_uop_3_27_ftq_idx;
  reg         rob_uop_3_27_edge_inst;
  reg  [5:0]  rob_uop_3_27_pc_lob;
  reg  [6:0]  rob_uop_3_27_pdst;
  reg  [6:0]  rob_uop_3_27_stale_pdst;
  reg         rob_uop_3_27_is_fencei;
  reg         rob_uop_3_27_uses_ldq;
  reg         rob_uop_3_27_uses_stq;
  reg         rob_uop_3_27_is_sys_pc2epc;
  reg         rob_uop_3_27_flush_on_commit;
  reg  [5:0]  rob_uop_3_27_ldst;
  reg         rob_uop_3_27_ldst_val;
  reg  [1:0]  rob_uop_3_27_dst_rtype;
  reg         rob_uop_3_27_fp_val;
  reg  [6:0]  rob_uop_3_28_uopc;
  reg         rob_uop_3_28_is_rvc;
  reg  [19:0] rob_uop_3_28_br_mask;
  reg  [5:0]  rob_uop_3_28_ftq_idx;
  reg         rob_uop_3_28_edge_inst;
  reg  [5:0]  rob_uop_3_28_pc_lob;
  reg  [6:0]  rob_uop_3_28_pdst;
  reg  [6:0]  rob_uop_3_28_stale_pdst;
  reg         rob_uop_3_28_is_fencei;
  reg         rob_uop_3_28_uses_ldq;
  reg         rob_uop_3_28_uses_stq;
  reg         rob_uop_3_28_is_sys_pc2epc;
  reg         rob_uop_3_28_flush_on_commit;
  reg  [5:0]  rob_uop_3_28_ldst;
  reg         rob_uop_3_28_ldst_val;
  reg  [1:0]  rob_uop_3_28_dst_rtype;
  reg         rob_uop_3_28_fp_val;
  reg  [6:0]  rob_uop_3_29_uopc;
  reg         rob_uop_3_29_is_rvc;
  reg  [19:0] rob_uop_3_29_br_mask;
  reg  [5:0]  rob_uop_3_29_ftq_idx;
  reg         rob_uop_3_29_edge_inst;
  reg  [5:0]  rob_uop_3_29_pc_lob;
  reg  [6:0]  rob_uop_3_29_pdst;
  reg  [6:0]  rob_uop_3_29_stale_pdst;
  reg         rob_uop_3_29_is_fencei;
  reg         rob_uop_3_29_uses_ldq;
  reg         rob_uop_3_29_uses_stq;
  reg         rob_uop_3_29_is_sys_pc2epc;
  reg         rob_uop_3_29_flush_on_commit;
  reg  [5:0]  rob_uop_3_29_ldst;
  reg         rob_uop_3_29_ldst_val;
  reg  [1:0]  rob_uop_3_29_dst_rtype;
  reg         rob_uop_3_29_fp_val;
  reg  [6:0]  rob_uop_3_30_uopc;
  reg         rob_uop_3_30_is_rvc;
  reg  [19:0] rob_uop_3_30_br_mask;
  reg  [5:0]  rob_uop_3_30_ftq_idx;
  reg         rob_uop_3_30_edge_inst;
  reg  [5:0]  rob_uop_3_30_pc_lob;
  reg  [6:0]  rob_uop_3_30_pdst;
  reg  [6:0]  rob_uop_3_30_stale_pdst;
  reg         rob_uop_3_30_is_fencei;
  reg         rob_uop_3_30_uses_ldq;
  reg         rob_uop_3_30_uses_stq;
  reg         rob_uop_3_30_is_sys_pc2epc;
  reg         rob_uop_3_30_flush_on_commit;
  reg  [5:0]  rob_uop_3_30_ldst;
  reg         rob_uop_3_30_ldst_val;
  reg  [1:0]  rob_uop_3_30_dst_rtype;
  reg         rob_uop_3_30_fp_val;
  reg  [6:0]  rob_uop_3_31_uopc;
  reg         rob_uop_3_31_is_rvc;
  reg  [19:0] rob_uop_3_31_br_mask;
  reg  [5:0]  rob_uop_3_31_ftq_idx;
  reg         rob_uop_3_31_edge_inst;
  reg  [5:0]  rob_uop_3_31_pc_lob;
  reg  [6:0]  rob_uop_3_31_pdst;
  reg  [6:0]  rob_uop_3_31_stale_pdst;
  reg         rob_uop_3_31_is_fencei;
  reg         rob_uop_3_31_uses_ldq;
  reg         rob_uop_3_31_uses_stq;
  reg         rob_uop_3_31_is_sys_pc2epc;
  reg         rob_uop_3_31_flush_on_commit;
  reg  [5:0]  rob_uop_3_31_ldst;
  reg         rob_uop_3_31_ldst_val;
  reg  [1:0]  rob_uop_3_31_dst_rtype;
  reg         rob_uop_3_31_fp_val;
  reg         rob_predicated_3_0;
  reg         rob_predicated_3_1;
  reg         rob_predicated_3_2;
  reg         rob_predicated_3_3;
  reg         rob_predicated_3_4;
  reg         rob_predicated_3_5;
  reg         rob_predicated_3_6;
  reg         rob_predicated_3_7;
  reg         rob_predicated_3_8;
  reg         rob_predicated_3_9;
  reg         rob_predicated_3_10;
  reg         rob_predicated_3_11;
  reg         rob_predicated_3_12;
  reg         rob_predicated_3_13;
  reg         rob_predicated_3_14;
  reg         rob_predicated_3_15;
  reg         rob_predicated_3_16;
  reg         rob_predicated_3_17;
  reg         rob_predicated_3_18;
  reg         rob_predicated_3_19;
  reg         rob_predicated_3_20;
  reg         rob_predicated_3_21;
  reg         rob_predicated_3_22;
  reg         rob_predicated_3_23;
  reg         rob_predicated_3_24;
  reg         rob_predicated_3_25;
  reg         rob_predicated_3_26;
  reg         rob_predicated_3_27;
  reg         rob_predicated_3_28;
  reg         rob_predicated_3_29;
  reg         rob_predicated_3_30;
  reg         rob_predicated_3_31;
  wire        _GEN_1822 = io_enq_valids_3 & _GEN_2;
  wire        _GEN_1823 = io_enq_valids_3 & _GEN_3;
  wire        _GEN_1824 = io_enq_valids_3 & _GEN_4;
  wire        _GEN_1825 = io_enq_valids_3 & _GEN_5;
  wire        _GEN_1826 = io_enq_valids_3 & _GEN_6;
  wire        _GEN_1827 = io_enq_valids_3 & _GEN_7;
  wire        _GEN_1828 = io_enq_valids_3 & _GEN_8;
  wire        _GEN_1829 = io_enq_valids_3 & _GEN_9;
  wire        _GEN_1830 = io_enq_valids_3 & _GEN_10;
  wire        _GEN_1831 = io_enq_valids_3 & _GEN_11;
  wire        _GEN_1832 = io_enq_valids_3 & _GEN_12;
  wire        _GEN_1833 = io_enq_valids_3 & _GEN_13;
  wire        _GEN_1834 = io_enq_valids_3 & _GEN_14;
  wire        _GEN_1835 = io_enq_valids_3 & _GEN_15;
  wire        _GEN_1836 = io_enq_valids_3 & _GEN_16;
  wire        _GEN_1837 = io_enq_valids_3 & _GEN_17;
  wire        _GEN_1838 = io_enq_valids_3 & _GEN_18;
  wire        _GEN_1839 = io_enq_valids_3 & _GEN_19;
  wire        _GEN_1840 = io_enq_valids_3 & _GEN_20;
  wire        _GEN_1841 = io_enq_valids_3 & _GEN_21;
  wire        _GEN_1842 = io_enq_valids_3 & _GEN_22;
  wire        _GEN_1843 = io_enq_valids_3 & _GEN_23;
  wire        _GEN_1844 = io_enq_valids_3 & _GEN_24;
  wire        _GEN_1845 = io_enq_valids_3 & _GEN_25;
  wire        _GEN_1846 = io_enq_valids_3 & _GEN_26;
  wire        _GEN_1847 = io_enq_valids_3 & _GEN_27;
  wire        _GEN_1848 = io_enq_valids_3 & _GEN_28;
  wire        _GEN_1849 = io_enq_valids_3 & _GEN_29;
  wire        _GEN_1850 = io_enq_valids_3 & _GEN_30;
  wire        _GEN_1851 = io_enq_valids_3 & _GEN_31;
  wire        _GEN_1852 = io_enq_valids_3 & _GEN_32;
  wire        _GEN_1853 = io_enq_valids_3 & (&rob_tail);
  wire        _GEN_1854 = io_wb_resps_0_valid & (&(io_wb_resps_0_bits_uop_rob_idx[1:0]));
  wire        _GEN_1855 = _GEN_1854 & _GEN_66;
  wire        _GEN_1856 = _GEN_1854 & _GEN_67;
  wire        _GEN_1857 = _GEN_1854 & _GEN_68;
  wire        _GEN_1858 = _GEN_1854 & _GEN_69;
  wire        _GEN_1859 = _GEN_1854 & _GEN_70;
  wire        _GEN_1860 = _GEN_1854 & _GEN_71;
  wire        _GEN_1861 = _GEN_1854 & _GEN_72;
  wire        _GEN_1862 = _GEN_1854 & _GEN_73;
  wire        _GEN_1863 = _GEN_1854 & _GEN_74;
  wire        _GEN_1864 = _GEN_1854 & _GEN_75;
  wire        _GEN_1865 = _GEN_1854 & _GEN_76;
  wire        _GEN_1866 = _GEN_1854 & _GEN_77;
  wire        _GEN_1867 = _GEN_1854 & _GEN_78;
  wire        _GEN_1868 = _GEN_1854 & _GEN_79;
  wire        _GEN_1869 = _GEN_1854 & _GEN_80;
  wire        _GEN_1870 = _GEN_1854 & _GEN_81;
  wire        _GEN_1871 = _GEN_1854 & _GEN_82;
  wire        _GEN_1872 = _GEN_1854 & _GEN_83;
  wire        _GEN_1873 = _GEN_1854 & _GEN_84;
  wire        _GEN_1874 = _GEN_1854 & _GEN_85;
  wire        _GEN_1875 = _GEN_1854 & _GEN_86;
  wire        _GEN_1876 = _GEN_1854 & _GEN_87;
  wire        _GEN_1877 = _GEN_1854 & _GEN_88;
  wire        _GEN_1878 = _GEN_1854 & _GEN_89;
  wire        _GEN_1879 = _GEN_1854 & _GEN_90;
  wire        _GEN_1880 = _GEN_1854 & _GEN_91;
  wire        _GEN_1881 = _GEN_1854 & _GEN_92;
  wire        _GEN_1882 = _GEN_1854 & _GEN_93;
  wire        _GEN_1883 = _GEN_1854 & _GEN_94;
  wire        _GEN_1884 = _GEN_1854 & _GEN_95;
  wire        _GEN_1885 = _GEN_1854 & _GEN_96;
  wire        _GEN_1886 = _GEN_1854 & (&(io_wb_resps_0_bits_uop_rob_idx[6:2]));
  wire        _GEN_1887 = io_wb_resps_1_valid & (&(io_wb_resps_1_bits_uop_rob_idx[1:0]));
  wire        _GEN_1888 = _GEN_130 | _GEN_1855;
  wire        _GEN_1889 = _GEN_132 | _GEN_1856;
  wire        _GEN_1890 = _GEN_134 | _GEN_1857;
  wire        _GEN_1891 = _GEN_136 | _GEN_1858;
  wire        _GEN_1892 = _GEN_138 | _GEN_1859;
  wire        _GEN_1893 = _GEN_140 | _GEN_1860;
  wire        _GEN_1894 = _GEN_142 | _GEN_1861;
  wire        _GEN_1895 = _GEN_144 | _GEN_1862;
  wire        _GEN_1896 = _GEN_146 | _GEN_1863;
  wire        _GEN_1897 = _GEN_148 | _GEN_1864;
  wire        _GEN_1898 = _GEN_150 | _GEN_1865;
  wire        _GEN_1899 = _GEN_152 | _GEN_1866;
  wire        _GEN_1900 = _GEN_154 | _GEN_1867;
  wire        _GEN_1901 = _GEN_156 | _GEN_1868;
  wire        _GEN_1902 = _GEN_158 | _GEN_1869;
  wire        _GEN_1903 = _GEN_160 | _GEN_1870;
  wire        _GEN_1904 = _GEN_162 | _GEN_1871;
  wire        _GEN_1905 = _GEN_164 | _GEN_1872;
  wire        _GEN_1906 = _GEN_166 | _GEN_1873;
  wire        _GEN_1907 = _GEN_168 | _GEN_1874;
  wire        _GEN_1908 = _GEN_170 | _GEN_1875;
  wire        _GEN_1909 = _GEN_172 | _GEN_1876;
  wire        _GEN_1910 = _GEN_174 | _GEN_1877;
  wire        _GEN_1911 = _GEN_176 | _GEN_1878;
  wire        _GEN_1912 = _GEN_178 | _GEN_1879;
  wire        _GEN_1913 = _GEN_180 | _GEN_1880;
  wire        _GEN_1914 = _GEN_182 | _GEN_1881;
  wire        _GEN_1915 = _GEN_184 | _GEN_1882;
  wire        _GEN_1916 = _GEN_186 | _GEN_1883;
  wire        _GEN_1917 = _GEN_188 | _GEN_1884;
  wire        _GEN_1918 = _GEN_190 | _GEN_1885;
  wire        _GEN_1919 = (&(io_wb_resps_1_bits_uop_rob_idx[6:2])) | _GEN_1886;
  wire        _GEN_1920 = io_wb_resps_2_valid & (&(io_wb_resps_2_bits_uop_rob_idx[1:0]));
  wire        _GEN_1921 = _GEN_1920 & _GEN_194;
  wire        _GEN_1922 = _GEN_1920 & _GEN_195;
  wire        _GEN_1923 = _GEN_1920 & _GEN_196;
  wire        _GEN_1924 = _GEN_1920 & _GEN_197;
  wire        _GEN_1925 = _GEN_1920 & _GEN_198;
  wire        _GEN_1926 = _GEN_1920 & _GEN_199;
  wire        _GEN_1927 = _GEN_1920 & _GEN_200;
  wire        _GEN_1928 = _GEN_1920 & _GEN_201;
  wire        _GEN_1929 = _GEN_1920 & _GEN_202;
  wire        _GEN_1930 = _GEN_1920 & _GEN_203;
  wire        _GEN_1931 = _GEN_1920 & _GEN_204;
  wire        _GEN_1932 = _GEN_1920 & _GEN_205;
  wire        _GEN_1933 = _GEN_1920 & _GEN_206;
  wire        _GEN_1934 = _GEN_1920 & _GEN_207;
  wire        _GEN_1935 = _GEN_1920 & _GEN_208;
  wire        _GEN_1936 = _GEN_1920 & _GEN_209;
  wire        _GEN_1937 = _GEN_1920 & _GEN_210;
  wire        _GEN_1938 = _GEN_1920 & _GEN_211;
  wire        _GEN_1939 = _GEN_1920 & _GEN_212;
  wire        _GEN_1940 = _GEN_1920 & _GEN_213;
  wire        _GEN_1941 = _GEN_1920 & _GEN_214;
  wire        _GEN_1942 = _GEN_1920 & _GEN_215;
  wire        _GEN_1943 = _GEN_1920 & _GEN_216;
  wire        _GEN_1944 = _GEN_1920 & _GEN_217;
  wire        _GEN_1945 = _GEN_1920 & _GEN_218;
  wire        _GEN_1946 = _GEN_1920 & _GEN_219;
  wire        _GEN_1947 = _GEN_1920 & _GEN_220;
  wire        _GEN_1948 = _GEN_1920 & _GEN_221;
  wire        _GEN_1949 = _GEN_1920 & _GEN_222;
  wire        _GEN_1950 = _GEN_1920 & _GEN_223;
  wire        _GEN_1951 = _GEN_1920 & _GEN_224;
  wire        _GEN_1952 = _GEN_1920 & (&(io_wb_resps_2_bits_uop_rob_idx[6:2]));
  wire        _GEN_1953 = io_wb_resps_3_valid & (&(io_wb_resps_3_bits_uop_rob_idx[1:0]));
  wire        _GEN_1954 = _GEN_258 | _GEN_1921;
  wire        _GEN_1955 = _GEN_260 | _GEN_1922;
  wire        _GEN_1956 = _GEN_262 | _GEN_1923;
  wire        _GEN_1957 = _GEN_264 | _GEN_1924;
  wire        _GEN_1958 = _GEN_266 | _GEN_1925;
  wire        _GEN_1959 = _GEN_268 | _GEN_1926;
  wire        _GEN_1960 = _GEN_270 | _GEN_1927;
  wire        _GEN_1961 = _GEN_272 | _GEN_1928;
  wire        _GEN_1962 = _GEN_274 | _GEN_1929;
  wire        _GEN_1963 = _GEN_276 | _GEN_1930;
  wire        _GEN_1964 = _GEN_278 | _GEN_1931;
  wire        _GEN_1965 = _GEN_280 | _GEN_1932;
  wire        _GEN_1966 = _GEN_282 | _GEN_1933;
  wire        _GEN_1967 = _GEN_284 | _GEN_1934;
  wire        _GEN_1968 = _GEN_286 | _GEN_1935;
  wire        _GEN_1969 = _GEN_288 | _GEN_1936;
  wire        _GEN_1970 = _GEN_290 | _GEN_1937;
  wire        _GEN_1971 = _GEN_292 | _GEN_1938;
  wire        _GEN_1972 = _GEN_294 | _GEN_1939;
  wire        _GEN_1973 = _GEN_296 | _GEN_1940;
  wire        _GEN_1974 = _GEN_298 | _GEN_1941;
  wire        _GEN_1975 = _GEN_300 | _GEN_1942;
  wire        _GEN_1976 = _GEN_302 | _GEN_1943;
  wire        _GEN_1977 = _GEN_304 | _GEN_1944;
  wire        _GEN_1978 = _GEN_306 | _GEN_1945;
  wire        _GEN_1979 = _GEN_308 | _GEN_1946;
  wire        _GEN_1980 = _GEN_310 | _GEN_1947;
  wire        _GEN_1981 = _GEN_312 | _GEN_1948;
  wire        _GEN_1982 = _GEN_314 | _GEN_1949;
  wire        _GEN_1983 = _GEN_316 | _GEN_1950;
  wire        _GEN_1984 = _GEN_318 | _GEN_1951;
  wire        _GEN_1985 = (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1952;
  wire        _GEN_1986 = io_wb_resps_4_valid & (&(io_wb_resps_4_bits_uop_rob_idx[1:0]));
  wire        _GEN_1987 = _GEN_1986 & _GEN_322;
  wire        _GEN_1988 = _GEN_1986 & _GEN_323;
  wire        _GEN_1989 = _GEN_1986 & _GEN_324;
  wire        _GEN_1990 = _GEN_1986 & _GEN_325;
  wire        _GEN_1991 = _GEN_1986 & _GEN_326;
  wire        _GEN_1992 = _GEN_1986 & _GEN_327;
  wire        _GEN_1993 = _GEN_1986 & _GEN_328;
  wire        _GEN_1994 = _GEN_1986 & _GEN_329;
  wire        _GEN_1995 = _GEN_1986 & _GEN_330;
  wire        _GEN_1996 = _GEN_1986 & _GEN_331;
  wire        _GEN_1997 = _GEN_1986 & _GEN_332;
  wire        _GEN_1998 = _GEN_1986 & _GEN_333;
  wire        _GEN_1999 = _GEN_1986 & _GEN_334;
  wire        _GEN_2000 = _GEN_1986 & _GEN_335;
  wire        _GEN_2001 = _GEN_1986 & _GEN_336;
  wire        _GEN_2002 = _GEN_1986 & _GEN_337;
  wire        _GEN_2003 = _GEN_1986 & _GEN_338;
  wire        _GEN_2004 = _GEN_1986 & _GEN_339;
  wire        _GEN_2005 = _GEN_1986 & _GEN_340;
  wire        _GEN_2006 = _GEN_1986 & _GEN_341;
  wire        _GEN_2007 = _GEN_1986 & _GEN_342;
  wire        _GEN_2008 = _GEN_1986 & _GEN_343;
  wire        _GEN_2009 = _GEN_1986 & _GEN_344;
  wire        _GEN_2010 = _GEN_1986 & _GEN_345;
  wire        _GEN_2011 = _GEN_1986 & _GEN_346;
  wire        _GEN_2012 = _GEN_1986 & _GEN_347;
  wire        _GEN_2013 = _GEN_1986 & _GEN_348;
  wire        _GEN_2014 = _GEN_1986 & _GEN_349;
  wire        _GEN_2015 = _GEN_1986 & _GEN_350;
  wire        _GEN_2016 = _GEN_1986 & _GEN_351;
  wire        _GEN_2017 = _GEN_1986 & _GEN_352;
  wire        _GEN_2018 = _GEN_1986 & (&(io_wb_resps_4_bits_uop_rob_idx[6:2]));
  wire        _GEN_2019 = io_wb_resps_5_valid & (&(io_wb_resps_5_bits_uop_rob_idx[1:0]));
  wire        _GEN_2020 = _GEN_386 | _GEN_1987;
  wire        _GEN_2021 = _GEN_388 | _GEN_1988;
  wire        _GEN_2022 = _GEN_390 | _GEN_1989;
  wire        _GEN_2023 = _GEN_392 | _GEN_1990;
  wire        _GEN_2024 = _GEN_394 | _GEN_1991;
  wire        _GEN_2025 = _GEN_396 | _GEN_1992;
  wire        _GEN_2026 = _GEN_398 | _GEN_1993;
  wire        _GEN_2027 = _GEN_400 | _GEN_1994;
  wire        _GEN_2028 = _GEN_402 | _GEN_1995;
  wire        _GEN_2029 = _GEN_404 | _GEN_1996;
  wire        _GEN_2030 = _GEN_406 | _GEN_1997;
  wire        _GEN_2031 = _GEN_408 | _GEN_1998;
  wire        _GEN_2032 = _GEN_410 | _GEN_1999;
  wire        _GEN_2033 = _GEN_412 | _GEN_2000;
  wire        _GEN_2034 = _GEN_414 | _GEN_2001;
  wire        _GEN_2035 = _GEN_416 | _GEN_2002;
  wire        _GEN_2036 = _GEN_418 | _GEN_2003;
  wire        _GEN_2037 = _GEN_420 | _GEN_2004;
  wire        _GEN_2038 = _GEN_422 | _GEN_2005;
  wire        _GEN_2039 = _GEN_424 | _GEN_2006;
  wire        _GEN_2040 = _GEN_426 | _GEN_2007;
  wire        _GEN_2041 = _GEN_428 | _GEN_2008;
  wire        _GEN_2042 = _GEN_430 | _GEN_2009;
  wire        _GEN_2043 = _GEN_432 | _GEN_2010;
  wire        _GEN_2044 = _GEN_434 | _GEN_2011;
  wire        _GEN_2045 = _GEN_436 | _GEN_2012;
  wire        _GEN_2046 = _GEN_438 | _GEN_2013;
  wire        _GEN_2047 = _GEN_440 | _GEN_2014;
  wire        _GEN_2048 = _GEN_442 | _GEN_2015;
  wire        _GEN_2049 = _GEN_444 | _GEN_2016;
  wire        _GEN_2050 = _GEN_446 | _GEN_2017;
  wire        _GEN_2051 = (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2018;
  wire        _GEN_2052 = io_wb_resps_6_valid & (&(io_wb_resps_6_bits_uop_rob_idx[1:0]));
  wire        _GEN_2053 = _GEN_2052 & _GEN_450;
  wire        _GEN_2054 = _GEN_2052 & _GEN_451;
  wire        _GEN_2055 = _GEN_2052 & _GEN_452;
  wire        _GEN_2056 = _GEN_2052 & _GEN_453;
  wire        _GEN_2057 = _GEN_2052 & _GEN_454;
  wire        _GEN_2058 = _GEN_2052 & _GEN_455;
  wire        _GEN_2059 = _GEN_2052 & _GEN_456;
  wire        _GEN_2060 = _GEN_2052 & _GEN_457;
  wire        _GEN_2061 = _GEN_2052 & _GEN_458;
  wire        _GEN_2062 = _GEN_2052 & _GEN_459;
  wire        _GEN_2063 = _GEN_2052 & _GEN_460;
  wire        _GEN_2064 = _GEN_2052 & _GEN_461;
  wire        _GEN_2065 = _GEN_2052 & _GEN_462;
  wire        _GEN_2066 = _GEN_2052 & _GEN_463;
  wire        _GEN_2067 = _GEN_2052 & _GEN_464;
  wire        _GEN_2068 = _GEN_2052 & _GEN_465;
  wire        _GEN_2069 = _GEN_2052 & _GEN_466;
  wire        _GEN_2070 = _GEN_2052 & _GEN_467;
  wire        _GEN_2071 = _GEN_2052 & _GEN_468;
  wire        _GEN_2072 = _GEN_2052 & _GEN_469;
  wire        _GEN_2073 = _GEN_2052 & _GEN_470;
  wire        _GEN_2074 = _GEN_2052 & _GEN_471;
  wire        _GEN_2075 = _GEN_2052 & _GEN_472;
  wire        _GEN_2076 = _GEN_2052 & _GEN_473;
  wire        _GEN_2077 = _GEN_2052 & _GEN_474;
  wire        _GEN_2078 = _GEN_2052 & _GEN_475;
  wire        _GEN_2079 = _GEN_2052 & _GEN_476;
  wire        _GEN_2080 = _GEN_2052 & _GEN_477;
  wire        _GEN_2081 = _GEN_2052 & _GEN_478;
  wire        _GEN_2082 = _GEN_2052 & _GEN_479;
  wire        _GEN_2083 = _GEN_2052 & _GEN_480;
  wire        _GEN_2084 = _GEN_2052 & (&(io_wb_resps_6_bits_uop_rob_idx[6:2]));
  wire        _GEN_2085 = io_wb_resps_7_valid & (&(io_wb_resps_7_bits_uop_rob_idx[1:0]));
  wire        _GEN_2086 = _GEN_514 | _GEN_2053;
  wire        _GEN_2087 = _GEN_516 | _GEN_2054;
  wire        _GEN_2088 = _GEN_518 | _GEN_2055;
  wire        _GEN_2089 = _GEN_520 | _GEN_2056;
  wire        _GEN_2090 = _GEN_522 | _GEN_2057;
  wire        _GEN_2091 = _GEN_524 | _GEN_2058;
  wire        _GEN_2092 = _GEN_526 | _GEN_2059;
  wire        _GEN_2093 = _GEN_528 | _GEN_2060;
  wire        _GEN_2094 = _GEN_530 | _GEN_2061;
  wire        _GEN_2095 = _GEN_532 | _GEN_2062;
  wire        _GEN_2096 = _GEN_534 | _GEN_2063;
  wire        _GEN_2097 = _GEN_536 | _GEN_2064;
  wire        _GEN_2098 = _GEN_538 | _GEN_2065;
  wire        _GEN_2099 = _GEN_540 | _GEN_2066;
  wire        _GEN_2100 = _GEN_542 | _GEN_2067;
  wire        _GEN_2101 = _GEN_544 | _GEN_2068;
  wire        _GEN_2102 = _GEN_546 | _GEN_2069;
  wire        _GEN_2103 = _GEN_548 | _GEN_2070;
  wire        _GEN_2104 = _GEN_550 | _GEN_2071;
  wire        _GEN_2105 = _GEN_552 | _GEN_2072;
  wire        _GEN_2106 = _GEN_554 | _GEN_2073;
  wire        _GEN_2107 = _GEN_556 | _GEN_2074;
  wire        _GEN_2108 = _GEN_558 | _GEN_2075;
  wire        _GEN_2109 = _GEN_560 | _GEN_2076;
  wire        _GEN_2110 = _GEN_562 | _GEN_2077;
  wire        _GEN_2111 = _GEN_564 | _GEN_2078;
  wire        _GEN_2112 = _GEN_566 | _GEN_2079;
  wire        _GEN_2113 = _GEN_568 | _GEN_2080;
  wire        _GEN_2114 = _GEN_570 | _GEN_2081;
  wire        _GEN_2115 = _GEN_572 | _GEN_2082;
  wire        _GEN_2116 = _GEN_574 | _GEN_2083;
  wire        _GEN_2117 = (&(io_wb_resps_7_bits_uop_rob_idx[6:2])) | _GEN_2084;
  wire        _GEN_2118 = io_wb_resps_8_valid & (&(io_wb_resps_8_bits_uop_rob_idx[1:0]));
  wire        _GEN_2119 = _GEN_2118 & _GEN_578;
  wire        _GEN_2120 = _GEN_2118 & _GEN_579;
  wire        _GEN_2121 = _GEN_2118 & _GEN_580;
  wire        _GEN_2122 = _GEN_2118 & _GEN_581;
  wire        _GEN_2123 = _GEN_2118 & _GEN_582;
  wire        _GEN_2124 = _GEN_2118 & _GEN_583;
  wire        _GEN_2125 = _GEN_2118 & _GEN_584;
  wire        _GEN_2126 = _GEN_2118 & _GEN_585;
  wire        _GEN_2127 = _GEN_2118 & _GEN_586;
  wire        _GEN_2128 = _GEN_2118 & _GEN_587;
  wire        _GEN_2129 = _GEN_2118 & _GEN_588;
  wire        _GEN_2130 = _GEN_2118 & _GEN_589;
  wire        _GEN_2131 = _GEN_2118 & _GEN_590;
  wire        _GEN_2132 = _GEN_2118 & _GEN_591;
  wire        _GEN_2133 = _GEN_2118 & _GEN_592;
  wire        _GEN_2134 = _GEN_2118 & _GEN_593;
  wire        _GEN_2135 = _GEN_2118 & _GEN_594;
  wire        _GEN_2136 = _GEN_2118 & _GEN_595;
  wire        _GEN_2137 = _GEN_2118 & _GEN_596;
  wire        _GEN_2138 = _GEN_2118 & _GEN_597;
  wire        _GEN_2139 = _GEN_2118 & _GEN_598;
  wire        _GEN_2140 = _GEN_2118 & _GEN_599;
  wire        _GEN_2141 = _GEN_2118 & _GEN_600;
  wire        _GEN_2142 = _GEN_2118 & _GEN_601;
  wire        _GEN_2143 = _GEN_2118 & _GEN_602;
  wire        _GEN_2144 = _GEN_2118 & _GEN_603;
  wire        _GEN_2145 = _GEN_2118 & _GEN_604;
  wire        _GEN_2146 = _GEN_2118 & _GEN_605;
  wire        _GEN_2147 = _GEN_2118 & _GEN_606;
  wire        _GEN_2148 = _GEN_2118 & _GEN_607;
  wire        _GEN_2149 = _GEN_2118 & _GEN_608;
  wire        _GEN_2150 = _GEN_2118 & (&(io_wb_resps_8_bits_uop_rob_idx[6:2]));
  wire        _GEN_2151 = io_wb_resps_9_valid & (&(io_wb_resps_9_bits_uop_rob_idx[1:0]));
  wire        _GEN_2152 = _GEN_642 | _GEN_2119;
  wire        _GEN_2153 = _GEN_644 | _GEN_2120;
  wire        _GEN_2154 = _GEN_646 | _GEN_2121;
  wire        _GEN_2155 = _GEN_648 | _GEN_2122;
  wire        _GEN_2156 = _GEN_650 | _GEN_2123;
  wire        _GEN_2157 = _GEN_652 | _GEN_2124;
  wire        _GEN_2158 = _GEN_654 | _GEN_2125;
  wire        _GEN_2159 = _GEN_656 | _GEN_2126;
  wire        _GEN_2160 = _GEN_658 | _GEN_2127;
  wire        _GEN_2161 = _GEN_660 | _GEN_2128;
  wire        _GEN_2162 = _GEN_662 | _GEN_2129;
  wire        _GEN_2163 = _GEN_664 | _GEN_2130;
  wire        _GEN_2164 = _GEN_666 | _GEN_2131;
  wire        _GEN_2165 = _GEN_668 | _GEN_2132;
  wire        _GEN_2166 = _GEN_670 | _GEN_2133;
  wire        _GEN_2167 = _GEN_672 | _GEN_2134;
  wire        _GEN_2168 = _GEN_674 | _GEN_2135;
  wire        _GEN_2169 = _GEN_676 | _GEN_2136;
  wire        _GEN_2170 = _GEN_678 | _GEN_2137;
  wire        _GEN_2171 = _GEN_680 | _GEN_2138;
  wire        _GEN_2172 = _GEN_682 | _GEN_2139;
  wire        _GEN_2173 = _GEN_684 | _GEN_2140;
  wire        _GEN_2174 = _GEN_686 | _GEN_2141;
  wire        _GEN_2175 = _GEN_688 | _GEN_2142;
  wire        _GEN_2176 = _GEN_690 | _GEN_2143;
  wire        _GEN_2177 = _GEN_692 | _GEN_2144;
  wire        _GEN_2178 = _GEN_694 | _GEN_2145;
  wire        _GEN_2179 = _GEN_696 | _GEN_2146;
  wire        _GEN_2180 = _GEN_698 | _GEN_2147;
  wire        _GEN_2181 = _GEN_700 | _GEN_2148;
  wire        _GEN_2182 = _GEN_702 | _GEN_2149;
  wire        _GEN_2183 = (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_2150;
  wire        _GEN_2184 = io_lsu_clr_bsy_0_valid & (&(io_lsu_clr_bsy_0_bits[1:0]));
  wire        _GEN_2185 = _GEN_2184 & _GEN_706;
  wire        _GEN_2186 = _GEN_2184 & _GEN_707;
  wire        _GEN_2187 = _GEN_2184 & _GEN_708;
  wire        _GEN_2188 = _GEN_2184 & _GEN_709;
  wire        _GEN_2189 = _GEN_2184 & _GEN_710;
  wire        _GEN_2190 = _GEN_2184 & _GEN_711;
  wire        _GEN_2191 = _GEN_2184 & _GEN_712;
  wire        _GEN_2192 = _GEN_2184 & _GEN_713;
  wire        _GEN_2193 = _GEN_2184 & _GEN_714;
  wire        _GEN_2194 = _GEN_2184 & _GEN_715;
  wire        _GEN_2195 = _GEN_2184 & _GEN_716;
  wire        _GEN_2196 = _GEN_2184 & _GEN_717;
  wire        _GEN_2197 = _GEN_2184 & _GEN_718;
  wire        _GEN_2198 = _GEN_2184 & _GEN_719;
  wire        _GEN_2199 = _GEN_2184 & _GEN_720;
  wire        _GEN_2200 = _GEN_2184 & _GEN_721;
  wire        _GEN_2201 = _GEN_2184 & _GEN_722;
  wire        _GEN_2202 = _GEN_2184 & _GEN_723;
  wire        _GEN_2203 = _GEN_2184 & _GEN_724;
  wire        _GEN_2204 = _GEN_2184 & _GEN_725;
  wire        _GEN_2205 = _GEN_2184 & _GEN_726;
  wire        _GEN_2206 = _GEN_2184 & _GEN_727;
  wire        _GEN_2207 = _GEN_2184 & _GEN_728;
  wire        _GEN_2208 = _GEN_2184 & _GEN_729;
  wire        _GEN_2209 = _GEN_2184 & _GEN_730;
  wire        _GEN_2210 = _GEN_2184 & _GEN_731;
  wire        _GEN_2211 = _GEN_2184 & _GEN_732;
  wire        _GEN_2212 = _GEN_2184 & _GEN_733;
  wire        _GEN_2213 = _GEN_2184 & _GEN_734;
  wire        _GEN_2214 = _GEN_2184 & _GEN_735;
  wire        _GEN_2215 = _GEN_2184 & _GEN_736;
  wire        _GEN_2216 = _GEN_2184 & (&(io_lsu_clr_bsy_0_bits[6:2]));
  wire        _GEN_2217 = io_lsu_clr_bsy_1_valid & (&(io_lsu_clr_bsy_1_bits[1:0]));
  wire        _GEN_2218 = _GEN_770 | _GEN_2185;
  wire        _GEN_2219 = _GEN_772 | _GEN_2186;
  wire        _GEN_2220 = _GEN_774 | _GEN_2187;
  wire        _GEN_2221 = _GEN_776 | _GEN_2188;
  wire        _GEN_2222 = _GEN_778 | _GEN_2189;
  wire        _GEN_2223 = _GEN_780 | _GEN_2190;
  wire        _GEN_2224 = _GEN_782 | _GEN_2191;
  wire        _GEN_2225 = _GEN_784 | _GEN_2192;
  wire        _GEN_2226 = _GEN_786 | _GEN_2193;
  wire        _GEN_2227 = _GEN_788 | _GEN_2194;
  wire        _GEN_2228 = _GEN_790 | _GEN_2195;
  wire        _GEN_2229 = _GEN_792 | _GEN_2196;
  wire        _GEN_2230 = _GEN_794 | _GEN_2197;
  wire        _GEN_2231 = _GEN_796 | _GEN_2198;
  wire        _GEN_2232 = _GEN_798 | _GEN_2199;
  wire        _GEN_2233 = _GEN_800 | _GEN_2200;
  wire        _GEN_2234 = _GEN_802 | _GEN_2201;
  wire        _GEN_2235 = _GEN_804 | _GEN_2202;
  wire        _GEN_2236 = _GEN_806 | _GEN_2203;
  wire        _GEN_2237 = _GEN_808 | _GEN_2204;
  wire        _GEN_2238 = _GEN_810 | _GEN_2205;
  wire        _GEN_2239 = _GEN_812 | _GEN_2206;
  wire        _GEN_2240 = _GEN_814 | _GEN_2207;
  wire        _GEN_2241 = _GEN_816 | _GEN_2208;
  wire        _GEN_2242 = _GEN_818 | _GEN_2209;
  wire        _GEN_2243 = _GEN_820 | _GEN_2210;
  wire        _GEN_2244 = _GEN_822 | _GEN_2211;
  wire        _GEN_2245 = _GEN_824 | _GEN_2212;
  wire        _GEN_2246 = _GEN_826 | _GEN_2213;
  wire        _GEN_2247 = _GEN_828 | _GEN_2214;
  wire        _GEN_2248 = _GEN_830 | _GEN_2215;
  wire        _GEN_2249 = (&(io_lsu_clr_bsy_1_bits[6:2])) | _GEN_2216;
  wire        _GEN_2250 = io_lsu_clr_bsy_2_valid & (&(io_lsu_clr_bsy_2_bits[1:0]));
  wire        _GEN_2251 = _GEN_2250 & _GEN_834;
  wire        _GEN_2252 = _GEN_2250 & _GEN_835;
  wire        _GEN_2253 = _GEN_2250 & _GEN_836;
  wire        _GEN_2254 = _GEN_2250 & _GEN_837;
  wire        _GEN_2255 = _GEN_2250 & _GEN_838;
  wire        _GEN_2256 = _GEN_2250 & _GEN_839;
  wire        _GEN_2257 = _GEN_2250 & _GEN_840;
  wire        _GEN_2258 = _GEN_2250 & _GEN_841;
  wire        _GEN_2259 = _GEN_2250 & _GEN_842;
  wire        _GEN_2260 = _GEN_2250 & _GEN_843;
  wire        _GEN_2261 = _GEN_2250 & _GEN_844;
  wire        _GEN_2262 = _GEN_2250 & _GEN_845;
  wire        _GEN_2263 = _GEN_2250 & _GEN_846;
  wire        _GEN_2264 = _GEN_2250 & _GEN_847;
  wire        _GEN_2265 = _GEN_2250 & _GEN_848;
  wire        _GEN_2266 = _GEN_2250 & _GEN_849;
  wire        _GEN_2267 = _GEN_2250 & _GEN_850;
  wire        _GEN_2268 = _GEN_2250 & _GEN_851;
  wire        _GEN_2269 = _GEN_2250 & _GEN_852;
  wire        _GEN_2270 = _GEN_2250 & _GEN_853;
  wire        _GEN_2271 = _GEN_2250 & _GEN_854;
  wire        _GEN_2272 = _GEN_2250 & _GEN_855;
  wire        _GEN_2273 = _GEN_2250 & _GEN_856;
  wire        _GEN_2274 = _GEN_2250 & _GEN_857;
  wire        _GEN_2275 = _GEN_2250 & _GEN_858;
  wire        _GEN_2276 = _GEN_2250 & _GEN_859;
  wire        _GEN_2277 = _GEN_2250 & _GEN_860;
  wire        _GEN_2278 = _GEN_2250 & _GEN_861;
  wire        _GEN_2279 = _GEN_2250 & _GEN_862;
  wire        _GEN_2280 = _GEN_2250 & _GEN_863;
  wire        _GEN_2281 = _GEN_2250 & _GEN_864;
  wire        _GEN_2282 = _GEN_2250 & (&(io_lsu_clr_bsy_2_bits[6:2]));
  wire        _GEN_2283 = io_lxcpt_valid & (&(io_lxcpt_bits_uop_rob_idx[1:0]));
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_71 = rob_predicated_3_0;
      5'b00001:
        casez_tmp_71 = rob_predicated_3_1;
      5'b00010:
        casez_tmp_71 = rob_predicated_3_2;
      5'b00011:
        casez_tmp_71 = rob_predicated_3_3;
      5'b00100:
        casez_tmp_71 = rob_predicated_3_4;
      5'b00101:
        casez_tmp_71 = rob_predicated_3_5;
      5'b00110:
        casez_tmp_71 = rob_predicated_3_6;
      5'b00111:
        casez_tmp_71 = rob_predicated_3_7;
      5'b01000:
        casez_tmp_71 = rob_predicated_3_8;
      5'b01001:
        casez_tmp_71 = rob_predicated_3_9;
      5'b01010:
        casez_tmp_71 = rob_predicated_3_10;
      5'b01011:
        casez_tmp_71 = rob_predicated_3_11;
      5'b01100:
        casez_tmp_71 = rob_predicated_3_12;
      5'b01101:
        casez_tmp_71 = rob_predicated_3_13;
      5'b01110:
        casez_tmp_71 = rob_predicated_3_14;
      5'b01111:
        casez_tmp_71 = rob_predicated_3_15;
      5'b10000:
        casez_tmp_71 = rob_predicated_3_16;
      5'b10001:
        casez_tmp_71 = rob_predicated_3_17;
      5'b10010:
        casez_tmp_71 = rob_predicated_3_18;
      5'b10011:
        casez_tmp_71 = rob_predicated_3_19;
      5'b10100:
        casez_tmp_71 = rob_predicated_3_20;
      5'b10101:
        casez_tmp_71 = rob_predicated_3_21;
      5'b10110:
        casez_tmp_71 = rob_predicated_3_22;
      5'b10111:
        casez_tmp_71 = rob_predicated_3_23;
      5'b11000:
        casez_tmp_71 = rob_predicated_3_24;
      5'b11001:
        casez_tmp_71 = rob_predicated_3_25;
      5'b11010:
        casez_tmp_71 = rob_predicated_3_26;
      5'b11011:
        casez_tmp_71 = rob_predicated_3_27;
      5'b11100:
        casez_tmp_71 = rob_predicated_3_28;
      5'b11101:
        casez_tmp_71 = rob_predicated_3_29;
      5'b11110:
        casez_tmp_71 = rob_predicated_3_30;
      default:
        casez_tmp_71 = rob_predicated_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_72 = rob_uop_3_0_uopc;
      5'b00001:
        casez_tmp_72 = rob_uop_3_1_uopc;
      5'b00010:
        casez_tmp_72 = rob_uop_3_2_uopc;
      5'b00011:
        casez_tmp_72 = rob_uop_3_3_uopc;
      5'b00100:
        casez_tmp_72 = rob_uop_3_4_uopc;
      5'b00101:
        casez_tmp_72 = rob_uop_3_5_uopc;
      5'b00110:
        casez_tmp_72 = rob_uop_3_6_uopc;
      5'b00111:
        casez_tmp_72 = rob_uop_3_7_uopc;
      5'b01000:
        casez_tmp_72 = rob_uop_3_8_uopc;
      5'b01001:
        casez_tmp_72 = rob_uop_3_9_uopc;
      5'b01010:
        casez_tmp_72 = rob_uop_3_10_uopc;
      5'b01011:
        casez_tmp_72 = rob_uop_3_11_uopc;
      5'b01100:
        casez_tmp_72 = rob_uop_3_12_uopc;
      5'b01101:
        casez_tmp_72 = rob_uop_3_13_uopc;
      5'b01110:
        casez_tmp_72 = rob_uop_3_14_uopc;
      5'b01111:
        casez_tmp_72 = rob_uop_3_15_uopc;
      5'b10000:
        casez_tmp_72 = rob_uop_3_16_uopc;
      5'b10001:
        casez_tmp_72 = rob_uop_3_17_uopc;
      5'b10010:
        casez_tmp_72 = rob_uop_3_18_uopc;
      5'b10011:
        casez_tmp_72 = rob_uop_3_19_uopc;
      5'b10100:
        casez_tmp_72 = rob_uop_3_20_uopc;
      5'b10101:
        casez_tmp_72 = rob_uop_3_21_uopc;
      5'b10110:
        casez_tmp_72 = rob_uop_3_22_uopc;
      5'b10111:
        casez_tmp_72 = rob_uop_3_23_uopc;
      5'b11000:
        casez_tmp_72 = rob_uop_3_24_uopc;
      5'b11001:
        casez_tmp_72 = rob_uop_3_25_uopc;
      5'b11010:
        casez_tmp_72 = rob_uop_3_26_uopc;
      5'b11011:
        casez_tmp_72 = rob_uop_3_27_uopc;
      5'b11100:
        casez_tmp_72 = rob_uop_3_28_uopc;
      5'b11101:
        casez_tmp_72 = rob_uop_3_29_uopc;
      5'b11110:
        casez_tmp_72 = rob_uop_3_30_uopc;
      default:
        casez_tmp_72 = rob_uop_3_31_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_73 = rob_uop_3_0_is_rvc;
      5'b00001:
        casez_tmp_73 = rob_uop_3_1_is_rvc;
      5'b00010:
        casez_tmp_73 = rob_uop_3_2_is_rvc;
      5'b00011:
        casez_tmp_73 = rob_uop_3_3_is_rvc;
      5'b00100:
        casez_tmp_73 = rob_uop_3_4_is_rvc;
      5'b00101:
        casez_tmp_73 = rob_uop_3_5_is_rvc;
      5'b00110:
        casez_tmp_73 = rob_uop_3_6_is_rvc;
      5'b00111:
        casez_tmp_73 = rob_uop_3_7_is_rvc;
      5'b01000:
        casez_tmp_73 = rob_uop_3_8_is_rvc;
      5'b01001:
        casez_tmp_73 = rob_uop_3_9_is_rvc;
      5'b01010:
        casez_tmp_73 = rob_uop_3_10_is_rvc;
      5'b01011:
        casez_tmp_73 = rob_uop_3_11_is_rvc;
      5'b01100:
        casez_tmp_73 = rob_uop_3_12_is_rvc;
      5'b01101:
        casez_tmp_73 = rob_uop_3_13_is_rvc;
      5'b01110:
        casez_tmp_73 = rob_uop_3_14_is_rvc;
      5'b01111:
        casez_tmp_73 = rob_uop_3_15_is_rvc;
      5'b10000:
        casez_tmp_73 = rob_uop_3_16_is_rvc;
      5'b10001:
        casez_tmp_73 = rob_uop_3_17_is_rvc;
      5'b10010:
        casez_tmp_73 = rob_uop_3_18_is_rvc;
      5'b10011:
        casez_tmp_73 = rob_uop_3_19_is_rvc;
      5'b10100:
        casez_tmp_73 = rob_uop_3_20_is_rvc;
      5'b10101:
        casez_tmp_73 = rob_uop_3_21_is_rvc;
      5'b10110:
        casez_tmp_73 = rob_uop_3_22_is_rvc;
      5'b10111:
        casez_tmp_73 = rob_uop_3_23_is_rvc;
      5'b11000:
        casez_tmp_73 = rob_uop_3_24_is_rvc;
      5'b11001:
        casez_tmp_73 = rob_uop_3_25_is_rvc;
      5'b11010:
        casez_tmp_73 = rob_uop_3_26_is_rvc;
      5'b11011:
        casez_tmp_73 = rob_uop_3_27_is_rvc;
      5'b11100:
        casez_tmp_73 = rob_uop_3_28_is_rvc;
      5'b11101:
        casez_tmp_73 = rob_uop_3_29_is_rvc;
      5'b11110:
        casez_tmp_73 = rob_uop_3_30_is_rvc;
      default:
        casez_tmp_73 = rob_uop_3_31_is_rvc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_74 = rob_uop_3_0_ftq_idx;
      5'b00001:
        casez_tmp_74 = rob_uop_3_1_ftq_idx;
      5'b00010:
        casez_tmp_74 = rob_uop_3_2_ftq_idx;
      5'b00011:
        casez_tmp_74 = rob_uop_3_3_ftq_idx;
      5'b00100:
        casez_tmp_74 = rob_uop_3_4_ftq_idx;
      5'b00101:
        casez_tmp_74 = rob_uop_3_5_ftq_idx;
      5'b00110:
        casez_tmp_74 = rob_uop_3_6_ftq_idx;
      5'b00111:
        casez_tmp_74 = rob_uop_3_7_ftq_idx;
      5'b01000:
        casez_tmp_74 = rob_uop_3_8_ftq_idx;
      5'b01001:
        casez_tmp_74 = rob_uop_3_9_ftq_idx;
      5'b01010:
        casez_tmp_74 = rob_uop_3_10_ftq_idx;
      5'b01011:
        casez_tmp_74 = rob_uop_3_11_ftq_idx;
      5'b01100:
        casez_tmp_74 = rob_uop_3_12_ftq_idx;
      5'b01101:
        casez_tmp_74 = rob_uop_3_13_ftq_idx;
      5'b01110:
        casez_tmp_74 = rob_uop_3_14_ftq_idx;
      5'b01111:
        casez_tmp_74 = rob_uop_3_15_ftq_idx;
      5'b10000:
        casez_tmp_74 = rob_uop_3_16_ftq_idx;
      5'b10001:
        casez_tmp_74 = rob_uop_3_17_ftq_idx;
      5'b10010:
        casez_tmp_74 = rob_uop_3_18_ftq_idx;
      5'b10011:
        casez_tmp_74 = rob_uop_3_19_ftq_idx;
      5'b10100:
        casez_tmp_74 = rob_uop_3_20_ftq_idx;
      5'b10101:
        casez_tmp_74 = rob_uop_3_21_ftq_idx;
      5'b10110:
        casez_tmp_74 = rob_uop_3_22_ftq_idx;
      5'b10111:
        casez_tmp_74 = rob_uop_3_23_ftq_idx;
      5'b11000:
        casez_tmp_74 = rob_uop_3_24_ftq_idx;
      5'b11001:
        casez_tmp_74 = rob_uop_3_25_ftq_idx;
      5'b11010:
        casez_tmp_74 = rob_uop_3_26_ftq_idx;
      5'b11011:
        casez_tmp_74 = rob_uop_3_27_ftq_idx;
      5'b11100:
        casez_tmp_74 = rob_uop_3_28_ftq_idx;
      5'b11101:
        casez_tmp_74 = rob_uop_3_29_ftq_idx;
      5'b11110:
        casez_tmp_74 = rob_uop_3_30_ftq_idx;
      default:
        casez_tmp_74 = rob_uop_3_31_ftq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_75 = rob_uop_3_0_edge_inst;
      5'b00001:
        casez_tmp_75 = rob_uop_3_1_edge_inst;
      5'b00010:
        casez_tmp_75 = rob_uop_3_2_edge_inst;
      5'b00011:
        casez_tmp_75 = rob_uop_3_3_edge_inst;
      5'b00100:
        casez_tmp_75 = rob_uop_3_4_edge_inst;
      5'b00101:
        casez_tmp_75 = rob_uop_3_5_edge_inst;
      5'b00110:
        casez_tmp_75 = rob_uop_3_6_edge_inst;
      5'b00111:
        casez_tmp_75 = rob_uop_3_7_edge_inst;
      5'b01000:
        casez_tmp_75 = rob_uop_3_8_edge_inst;
      5'b01001:
        casez_tmp_75 = rob_uop_3_9_edge_inst;
      5'b01010:
        casez_tmp_75 = rob_uop_3_10_edge_inst;
      5'b01011:
        casez_tmp_75 = rob_uop_3_11_edge_inst;
      5'b01100:
        casez_tmp_75 = rob_uop_3_12_edge_inst;
      5'b01101:
        casez_tmp_75 = rob_uop_3_13_edge_inst;
      5'b01110:
        casez_tmp_75 = rob_uop_3_14_edge_inst;
      5'b01111:
        casez_tmp_75 = rob_uop_3_15_edge_inst;
      5'b10000:
        casez_tmp_75 = rob_uop_3_16_edge_inst;
      5'b10001:
        casez_tmp_75 = rob_uop_3_17_edge_inst;
      5'b10010:
        casez_tmp_75 = rob_uop_3_18_edge_inst;
      5'b10011:
        casez_tmp_75 = rob_uop_3_19_edge_inst;
      5'b10100:
        casez_tmp_75 = rob_uop_3_20_edge_inst;
      5'b10101:
        casez_tmp_75 = rob_uop_3_21_edge_inst;
      5'b10110:
        casez_tmp_75 = rob_uop_3_22_edge_inst;
      5'b10111:
        casez_tmp_75 = rob_uop_3_23_edge_inst;
      5'b11000:
        casez_tmp_75 = rob_uop_3_24_edge_inst;
      5'b11001:
        casez_tmp_75 = rob_uop_3_25_edge_inst;
      5'b11010:
        casez_tmp_75 = rob_uop_3_26_edge_inst;
      5'b11011:
        casez_tmp_75 = rob_uop_3_27_edge_inst;
      5'b11100:
        casez_tmp_75 = rob_uop_3_28_edge_inst;
      5'b11101:
        casez_tmp_75 = rob_uop_3_29_edge_inst;
      5'b11110:
        casez_tmp_75 = rob_uop_3_30_edge_inst;
      default:
        casez_tmp_75 = rob_uop_3_31_edge_inst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_76 = rob_uop_3_0_pc_lob;
      5'b00001:
        casez_tmp_76 = rob_uop_3_1_pc_lob;
      5'b00010:
        casez_tmp_76 = rob_uop_3_2_pc_lob;
      5'b00011:
        casez_tmp_76 = rob_uop_3_3_pc_lob;
      5'b00100:
        casez_tmp_76 = rob_uop_3_4_pc_lob;
      5'b00101:
        casez_tmp_76 = rob_uop_3_5_pc_lob;
      5'b00110:
        casez_tmp_76 = rob_uop_3_6_pc_lob;
      5'b00111:
        casez_tmp_76 = rob_uop_3_7_pc_lob;
      5'b01000:
        casez_tmp_76 = rob_uop_3_8_pc_lob;
      5'b01001:
        casez_tmp_76 = rob_uop_3_9_pc_lob;
      5'b01010:
        casez_tmp_76 = rob_uop_3_10_pc_lob;
      5'b01011:
        casez_tmp_76 = rob_uop_3_11_pc_lob;
      5'b01100:
        casez_tmp_76 = rob_uop_3_12_pc_lob;
      5'b01101:
        casez_tmp_76 = rob_uop_3_13_pc_lob;
      5'b01110:
        casez_tmp_76 = rob_uop_3_14_pc_lob;
      5'b01111:
        casez_tmp_76 = rob_uop_3_15_pc_lob;
      5'b10000:
        casez_tmp_76 = rob_uop_3_16_pc_lob;
      5'b10001:
        casez_tmp_76 = rob_uop_3_17_pc_lob;
      5'b10010:
        casez_tmp_76 = rob_uop_3_18_pc_lob;
      5'b10011:
        casez_tmp_76 = rob_uop_3_19_pc_lob;
      5'b10100:
        casez_tmp_76 = rob_uop_3_20_pc_lob;
      5'b10101:
        casez_tmp_76 = rob_uop_3_21_pc_lob;
      5'b10110:
        casez_tmp_76 = rob_uop_3_22_pc_lob;
      5'b10111:
        casez_tmp_76 = rob_uop_3_23_pc_lob;
      5'b11000:
        casez_tmp_76 = rob_uop_3_24_pc_lob;
      5'b11001:
        casez_tmp_76 = rob_uop_3_25_pc_lob;
      5'b11010:
        casez_tmp_76 = rob_uop_3_26_pc_lob;
      5'b11011:
        casez_tmp_76 = rob_uop_3_27_pc_lob;
      5'b11100:
        casez_tmp_76 = rob_uop_3_28_pc_lob;
      5'b11101:
        casez_tmp_76 = rob_uop_3_29_pc_lob;
      5'b11110:
        casez_tmp_76 = rob_uop_3_30_pc_lob;
      default:
        casez_tmp_76 = rob_uop_3_31_pc_lob;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_77 = rob_uop_3_0_pdst;
      5'b00001:
        casez_tmp_77 = rob_uop_3_1_pdst;
      5'b00010:
        casez_tmp_77 = rob_uop_3_2_pdst;
      5'b00011:
        casez_tmp_77 = rob_uop_3_3_pdst;
      5'b00100:
        casez_tmp_77 = rob_uop_3_4_pdst;
      5'b00101:
        casez_tmp_77 = rob_uop_3_5_pdst;
      5'b00110:
        casez_tmp_77 = rob_uop_3_6_pdst;
      5'b00111:
        casez_tmp_77 = rob_uop_3_7_pdst;
      5'b01000:
        casez_tmp_77 = rob_uop_3_8_pdst;
      5'b01001:
        casez_tmp_77 = rob_uop_3_9_pdst;
      5'b01010:
        casez_tmp_77 = rob_uop_3_10_pdst;
      5'b01011:
        casez_tmp_77 = rob_uop_3_11_pdst;
      5'b01100:
        casez_tmp_77 = rob_uop_3_12_pdst;
      5'b01101:
        casez_tmp_77 = rob_uop_3_13_pdst;
      5'b01110:
        casez_tmp_77 = rob_uop_3_14_pdst;
      5'b01111:
        casez_tmp_77 = rob_uop_3_15_pdst;
      5'b10000:
        casez_tmp_77 = rob_uop_3_16_pdst;
      5'b10001:
        casez_tmp_77 = rob_uop_3_17_pdst;
      5'b10010:
        casez_tmp_77 = rob_uop_3_18_pdst;
      5'b10011:
        casez_tmp_77 = rob_uop_3_19_pdst;
      5'b10100:
        casez_tmp_77 = rob_uop_3_20_pdst;
      5'b10101:
        casez_tmp_77 = rob_uop_3_21_pdst;
      5'b10110:
        casez_tmp_77 = rob_uop_3_22_pdst;
      5'b10111:
        casez_tmp_77 = rob_uop_3_23_pdst;
      5'b11000:
        casez_tmp_77 = rob_uop_3_24_pdst;
      5'b11001:
        casez_tmp_77 = rob_uop_3_25_pdst;
      5'b11010:
        casez_tmp_77 = rob_uop_3_26_pdst;
      5'b11011:
        casez_tmp_77 = rob_uop_3_27_pdst;
      5'b11100:
        casez_tmp_77 = rob_uop_3_28_pdst;
      5'b11101:
        casez_tmp_77 = rob_uop_3_29_pdst;
      5'b11110:
        casez_tmp_77 = rob_uop_3_30_pdst;
      default:
        casez_tmp_77 = rob_uop_3_31_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_78 = rob_uop_3_0_stale_pdst;
      5'b00001:
        casez_tmp_78 = rob_uop_3_1_stale_pdst;
      5'b00010:
        casez_tmp_78 = rob_uop_3_2_stale_pdst;
      5'b00011:
        casez_tmp_78 = rob_uop_3_3_stale_pdst;
      5'b00100:
        casez_tmp_78 = rob_uop_3_4_stale_pdst;
      5'b00101:
        casez_tmp_78 = rob_uop_3_5_stale_pdst;
      5'b00110:
        casez_tmp_78 = rob_uop_3_6_stale_pdst;
      5'b00111:
        casez_tmp_78 = rob_uop_3_7_stale_pdst;
      5'b01000:
        casez_tmp_78 = rob_uop_3_8_stale_pdst;
      5'b01001:
        casez_tmp_78 = rob_uop_3_9_stale_pdst;
      5'b01010:
        casez_tmp_78 = rob_uop_3_10_stale_pdst;
      5'b01011:
        casez_tmp_78 = rob_uop_3_11_stale_pdst;
      5'b01100:
        casez_tmp_78 = rob_uop_3_12_stale_pdst;
      5'b01101:
        casez_tmp_78 = rob_uop_3_13_stale_pdst;
      5'b01110:
        casez_tmp_78 = rob_uop_3_14_stale_pdst;
      5'b01111:
        casez_tmp_78 = rob_uop_3_15_stale_pdst;
      5'b10000:
        casez_tmp_78 = rob_uop_3_16_stale_pdst;
      5'b10001:
        casez_tmp_78 = rob_uop_3_17_stale_pdst;
      5'b10010:
        casez_tmp_78 = rob_uop_3_18_stale_pdst;
      5'b10011:
        casez_tmp_78 = rob_uop_3_19_stale_pdst;
      5'b10100:
        casez_tmp_78 = rob_uop_3_20_stale_pdst;
      5'b10101:
        casez_tmp_78 = rob_uop_3_21_stale_pdst;
      5'b10110:
        casez_tmp_78 = rob_uop_3_22_stale_pdst;
      5'b10111:
        casez_tmp_78 = rob_uop_3_23_stale_pdst;
      5'b11000:
        casez_tmp_78 = rob_uop_3_24_stale_pdst;
      5'b11001:
        casez_tmp_78 = rob_uop_3_25_stale_pdst;
      5'b11010:
        casez_tmp_78 = rob_uop_3_26_stale_pdst;
      5'b11011:
        casez_tmp_78 = rob_uop_3_27_stale_pdst;
      5'b11100:
        casez_tmp_78 = rob_uop_3_28_stale_pdst;
      5'b11101:
        casez_tmp_78 = rob_uop_3_29_stale_pdst;
      5'b11110:
        casez_tmp_78 = rob_uop_3_30_stale_pdst;
      default:
        casez_tmp_78 = rob_uop_3_31_stale_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_79 = rob_uop_3_0_is_fencei;
      5'b00001:
        casez_tmp_79 = rob_uop_3_1_is_fencei;
      5'b00010:
        casez_tmp_79 = rob_uop_3_2_is_fencei;
      5'b00011:
        casez_tmp_79 = rob_uop_3_3_is_fencei;
      5'b00100:
        casez_tmp_79 = rob_uop_3_4_is_fencei;
      5'b00101:
        casez_tmp_79 = rob_uop_3_5_is_fencei;
      5'b00110:
        casez_tmp_79 = rob_uop_3_6_is_fencei;
      5'b00111:
        casez_tmp_79 = rob_uop_3_7_is_fencei;
      5'b01000:
        casez_tmp_79 = rob_uop_3_8_is_fencei;
      5'b01001:
        casez_tmp_79 = rob_uop_3_9_is_fencei;
      5'b01010:
        casez_tmp_79 = rob_uop_3_10_is_fencei;
      5'b01011:
        casez_tmp_79 = rob_uop_3_11_is_fencei;
      5'b01100:
        casez_tmp_79 = rob_uop_3_12_is_fencei;
      5'b01101:
        casez_tmp_79 = rob_uop_3_13_is_fencei;
      5'b01110:
        casez_tmp_79 = rob_uop_3_14_is_fencei;
      5'b01111:
        casez_tmp_79 = rob_uop_3_15_is_fencei;
      5'b10000:
        casez_tmp_79 = rob_uop_3_16_is_fencei;
      5'b10001:
        casez_tmp_79 = rob_uop_3_17_is_fencei;
      5'b10010:
        casez_tmp_79 = rob_uop_3_18_is_fencei;
      5'b10011:
        casez_tmp_79 = rob_uop_3_19_is_fencei;
      5'b10100:
        casez_tmp_79 = rob_uop_3_20_is_fencei;
      5'b10101:
        casez_tmp_79 = rob_uop_3_21_is_fencei;
      5'b10110:
        casez_tmp_79 = rob_uop_3_22_is_fencei;
      5'b10111:
        casez_tmp_79 = rob_uop_3_23_is_fencei;
      5'b11000:
        casez_tmp_79 = rob_uop_3_24_is_fencei;
      5'b11001:
        casez_tmp_79 = rob_uop_3_25_is_fencei;
      5'b11010:
        casez_tmp_79 = rob_uop_3_26_is_fencei;
      5'b11011:
        casez_tmp_79 = rob_uop_3_27_is_fencei;
      5'b11100:
        casez_tmp_79 = rob_uop_3_28_is_fencei;
      5'b11101:
        casez_tmp_79 = rob_uop_3_29_is_fencei;
      5'b11110:
        casez_tmp_79 = rob_uop_3_30_is_fencei;
      default:
        casez_tmp_79 = rob_uop_3_31_is_fencei;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_80 = rob_uop_3_0_uses_ldq;
      5'b00001:
        casez_tmp_80 = rob_uop_3_1_uses_ldq;
      5'b00010:
        casez_tmp_80 = rob_uop_3_2_uses_ldq;
      5'b00011:
        casez_tmp_80 = rob_uop_3_3_uses_ldq;
      5'b00100:
        casez_tmp_80 = rob_uop_3_4_uses_ldq;
      5'b00101:
        casez_tmp_80 = rob_uop_3_5_uses_ldq;
      5'b00110:
        casez_tmp_80 = rob_uop_3_6_uses_ldq;
      5'b00111:
        casez_tmp_80 = rob_uop_3_7_uses_ldq;
      5'b01000:
        casez_tmp_80 = rob_uop_3_8_uses_ldq;
      5'b01001:
        casez_tmp_80 = rob_uop_3_9_uses_ldq;
      5'b01010:
        casez_tmp_80 = rob_uop_3_10_uses_ldq;
      5'b01011:
        casez_tmp_80 = rob_uop_3_11_uses_ldq;
      5'b01100:
        casez_tmp_80 = rob_uop_3_12_uses_ldq;
      5'b01101:
        casez_tmp_80 = rob_uop_3_13_uses_ldq;
      5'b01110:
        casez_tmp_80 = rob_uop_3_14_uses_ldq;
      5'b01111:
        casez_tmp_80 = rob_uop_3_15_uses_ldq;
      5'b10000:
        casez_tmp_80 = rob_uop_3_16_uses_ldq;
      5'b10001:
        casez_tmp_80 = rob_uop_3_17_uses_ldq;
      5'b10010:
        casez_tmp_80 = rob_uop_3_18_uses_ldq;
      5'b10011:
        casez_tmp_80 = rob_uop_3_19_uses_ldq;
      5'b10100:
        casez_tmp_80 = rob_uop_3_20_uses_ldq;
      5'b10101:
        casez_tmp_80 = rob_uop_3_21_uses_ldq;
      5'b10110:
        casez_tmp_80 = rob_uop_3_22_uses_ldq;
      5'b10111:
        casez_tmp_80 = rob_uop_3_23_uses_ldq;
      5'b11000:
        casez_tmp_80 = rob_uop_3_24_uses_ldq;
      5'b11001:
        casez_tmp_80 = rob_uop_3_25_uses_ldq;
      5'b11010:
        casez_tmp_80 = rob_uop_3_26_uses_ldq;
      5'b11011:
        casez_tmp_80 = rob_uop_3_27_uses_ldq;
      5'b11100:
        casez_tmp_80 = rob_uop_3_28_uses_ldq;
      5'b11101:
        casez_tmp_80 = rob_uop_3_29_uses_ldq;
      5'b11110:
        casez_tmp_80 = rob_uop_3_30_uses_ldq;
      default:
        casez_tmp_80 = rob_uop_3_31_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_81 = rob_uop_3_0_uses_stq;
      5'b00001:
        casez_tmp_81 = rob_uop_3_1_uses_stq;
      5'b00010:
        casez_tmp_81 = rob_uop_3_2_uses_stq;
      5'b00011:
        casez_tmp_81 = rob_uop_3_3_uses_stq;
      5'b00100:
        casez_tmp_81 = rob_uop_3_4_uses_stq;
      5'b00101:
        casez_tmp_81 = rob_uop_3_5_uses_stq;
      5'b00110:
        casez_tmp_81 = rob_uop_3_6_uses_stq;
      5'b00111:
        casez_tmp_81 = rob_uop_3_7_uses_stq;
      5'b01000:
        casez_tmp_81 = rob_uop_3_8_uses_stq;
      5'b01001:
        casez_tmp_81 = rob_uop_3_9_uses_stq;
      5'b01010:
        casez_tmp_81 = rob_uop_3_10_uses_stq;
      5'b01011:
        casez_tmp_81 = rob_uop_3_11_uses_stq;
      5'b01100:
        casez_tmp_81 = rob_uop_3_12_uses_stq;
      5'b01101:
        casez_tmp_81 = rob_uop_3_13_uses_stq;
      5'b01110:
        casez_tmp_81 = rob_uop_3_14_uses_stq;
      5'b01111:
        casez_tmp_81 = rob_uop_3_15_uses_stq;
      5'b10000:
        casez_tmp_81 = rob_uop_3_16_uses_stq;
      5'b10001:
        casez_tmp_81 = rob_uop_3_17_uses_stq;
      5'b10010:
        casez_tmp_81 = rob_uop_3_18_uses_stq;
      5'b10011:
        casez_tmp_81 = rob_uop_3_19_uses_stq;
      5'b10100:
        casez_tmp_81 = rob_uop_3_20_uses_stq;
      5'b10101:
        casez_tmp_81 = rob_uop_3_21_uses_stq;
      5'b10110:
        casez_tmp_81 = rob_uop_3_22_uses_stq;
      5'b10111:
        casez_tmp_81 = rob_uop_3_23_uses_stq;
      5'b11000:
        casez_tmp_81 = rob_uop_3_24_uses_stq;
      5'b11001:
        casez_tmp_81 = rob_uop_3_25_uses_stq;
      5'b11010:
        casez_tmp_81 = rob_uop_3_26_uses_stq;
      5'b11011:
        casez_tmp_81 = rob_uop_3_27_uses_stq;
      5'b11100:
        casez_tmp_81 = rob_uop_3_28_uses_stq;
      5'b11101:
        casez_tmp_81 = rob_uop_3_29_uses_stq;
      5'b11110:
        casez_tmp_81 = rob_uop_3_30_uses_stq;
      default:
        casez_tmp_81 = rob_uop_3_31_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_82 = rob_uop_3_0_is_sys_pc2epc;
      5'b00001:
        casez_tmp_82 = rob_uop_3_1_is_sys_pc2epc;
      5'b00010:
        casez_tmp_82 = rob_uop_3_2_is_sys_pc2epc;
      5'b00011:
        casez_tmp_82 = rob_uop_3_3_is_sys_pc2epc;
      5'b00100:
        casez_tmp_82 = rob_uop_3_4_is_sys_pc2epc;
      5'b00101:
        casez_tmp_82 = rob_uop_3_5_is_sys_pc2epc;
      5'b00110:
        casez_tmp_82 = rob_uop_3_6_is_sys_pc2epc;
      5'b00111:
        casez_tmp_82 = rob_uop_3_7_is_sys_pc2epc;
      5'b01000:
        casez_tmp_82 = rob_uop_3_8_is_sys_pc2epc;
      5'b01001:
        casez_tmp_82 = rob_uop_3_9_is_sys_pc2epc;
      5'b01010:
        casez_tmp_82 = rob_uop_3_10_is_sys_pc2epc;
      5'b01011:
        casez_tmp_82 = rob_uop_3_11_is_sys_pc2epc;
      5'b01100:
        casez_tmp_82 = rob_uop_3_12_is_sys_pc2epc;
      5'b01101:
        casez_tmp_82 = rob_uop_3_13_is_sys_pc2epc;
      5'b01110:
        casez_tmp_82 = rob_uop_3_14_is_sys_pc2epc;
      5'b01111:
        casez_tmp_82 = rob_uop_3_15_is_sys_pc2epc;
      5'b10000:
        casez_tmp_82 = rob_uop_3_16_is_sys_pc2epc;
      5'b10001:
        casez_tmp_82 = rob_uop_3_17_is_sys_pc2epc;
      5'b10010:
        casez_tmp_82 = rob_uop_3_18_is_sys_pc2epc;
      5'b10011:
        casez_tmp_82 = rob_uop_3_19_is_sys_pc2epc;
      5'b10100:
        casez_tmp_82 = rob_uop_3_20_is_sys_pc2epc;
      5'b10101:
        casez_tmp_82 = rob_uop_3_21_is_sys_pc2epc;
      5'b10110:
        casez_tmp_82 = rob_uop_3_22_is_sys_pc2epc;
      5'b10111:
        casez_tmp_82 = rob_uop_3_23_is_sys_pc2epc;
      5'b11000:
        casez_tmp_82 = rob_uop_3_24_is_sys_pc2epc;
      5'b11001:
        casez_tmp_82 = rob_uop_3_25_is_sys_pc2epc;
      5'b11010:
        casez_tmp_82 = rob_uop_3_26_is_sys_pc2epc;
      5'b11011:
        casez_tmp_82 = rob_uop_3_27_is_sys_pc2epc;
      5'b11100:
        casez_tmp_82 = rob_uop_3_28_is_sys_pc2epc;
      5'b11101:
        casez_tmp_82 = rob_uop_3_29_is_sys_pc2epc;
      5'b11110:
        casez_tmp_82 = rob_uop_3_30_is_sys_pc2epc;
      default:
        casez_tmp_82 = rob_uop_3_31_is_sys_pc2epc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_83 = rob_uop_3_0_flush_on_commit;
      5'b00001:
        casez_tmp_83 = rob_uop_3_1_flush_on_commit;
      5'b00010:
        casez_tmp_83 = rob_uop_3_2_flush_on_commit;
      5'b00011:
        casez_tmp_83 = rob_uop_3_3_flush_on_commit;
      5'b00100:
        casez_tmp_83 = rob_uop_3_4_flush_on_commit;
      5'b00101:
        casez_tmp_83 = rob_uop_3_5_flush_on_commit;
      5'b00110:
        casez_tmp_83 = rob_uop_3_6_flush_on_commit;
      5'b00111:
        casez_tmp_83 = rob_uop_3_7_flush_on_commit;
      5'b01000:
        casez_tmp_83 = rob_uop_3_8_flush_on_commit;
      5'b01001:
        casez_tmp_83 = rob_uop_3_9_flush_on_commit;
      5'b01010:
        casez_tmp_83 = rob_uop_3_10_flush_on_commit;
      5'b01011:
        casez_tmp_83 = rob_uop_3_11_flush_on_commit;
      5'b01100:
        casez_tmp_83 = rob_uop_3_12_flush_on_commit;
      5'b01101:
        casez_tmp_83 = rob_uop_3_13_flush_on_commit;
      5'b01110:
        casez_tmp_83 = rob_uop_3_14_flush_on_commit;
      5'b01111:
        casez_tmp_83 = rob_uop_3_15_flush_on_commit;
      5'b10000:
        casez_tmp_83 = rob_uop_3_16_flush_on_commit;
      5'b10001:
        casez_tmp_83 = rob_uop_3_17_flush_on_commit;
      5'b10010:
        casez_tmp_83 = rob_uop_3_18_flush_on_commit;
      5'b10011:
        casez_tmp_83 = rob_uop_3_19_flush_on_commit;
      5'b10100:
        casez_tmp_83 = rob_uop_3_20_flush_on_commit;
      5'b10101:
        casez_tmp_83 = rob_uop_3_21_flush_on_commit;
      5'b10110:
        casez_tmp_83 = rob_uop_3_22_flush_on_commit;
      5'b10111:
        casez_tmp_83 = rob_uop_3_23_flush_on_commit;
      5'b11000:
        casez_tmp_83 = rob_uop_3_24_flush_on_commit;
      5'b11001:
        casez_tmp_83 = rob_uop_3_25_flush_on_commit;
      5'b11010:
        casez_tmp_83 = rob_uop_3_26_flush_on_commit;
      5'b11011:
        casez_tmp_83 = rob_uop_3_27_flush_on_commit;
      5'b11100:
        casez_tmp_83 = rob_uop_3_28_flush_on_commit;
      5'b11101:
        casez_tmp_83 = rob_uop_3_29_flush_on_commit;
      5'b11110:
        casez_tmp_83 = rob_uop_3_30_flush_on_commit;
      default:
        casez_tmp_83 = rob_uop_3_31_flush_on_commit;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_84 = rob_uop_3_0_ldst;
      5'b00001:
        casez_tmp_84 = rob_uop_3_1_ldst;
      5'b00010:
        casez_tmp_84 = rob_uop_3_2_ldst;
      5'b00011:
        casez_tmp_84 = rob_uop_3_3_ldst;
      5'b00100:
        casez_tmp_84 = rob_uop_3_4_ldst;
      5'b00101:
        casez_tmp_84 = rob_uop_3_5_ldst;
      5'b00110:
        casez_tmp_84 = rob_uop_3_6_ldst;
      5'b00111:
        casez_tmp_84 = rob_uop_3_7_ldst;
      5'b01000:
        casez_tmp_84 = rob_uop_3_8_ldst;
      5'b01001:
        casez_tmp_84 = rob_uop_3_9_ldst;
      5'b01010:
        casez_tmp_84 = rob_uop_3_10_ldst;
      5'b01011:
        casez_tmp_84 = rob_uop_3_11_ldst;
      5'b01100:
        casez_tmp_84 = rob_uop_3_12_ldst;
      5'b01101:
        casez_tmp_84 = rob_uop_3_13_ldst;
      5'b01110:
        casez_tmp_84 = rob_uop_3_14_ldst;
      5'b01111:
        casez_tmp_84 = rob_uop_3_15_ldst;
      5'b10000:
        casez_tmp_84 = rob_uop_3_16_ldst;
      5'b10001:
        casez_tmp_84 = rob_uop_3_17_ldst;
      5'b10010:
        casez_tmp_84 = rob_uop_3_18_ldst;
      5'b10011:
        casez_tmp_84 = rob_uop_3_19_ldst;
      5'b10100:
        casez_tmp_84 = rob_uop_3_20_ldst;
      5'b10101:
        casez_tmp_84 = rob_uop_3_21_ldst;
      5'b10110:
        casez_tmp_84 = rob_uop_3_22_ldst;
      5'b10111:
        casez_tmp_84 = rob_uop_3_23_ldst;
      5'b11000:
        casez_tmp_84 = rob_uop_3_24_ldst;
      5'b11001:
        casez_tmp_84 = rob_uop_3_25_ldst;
      5'b11010:
        casez_tmp_84 = rob_uop_3_26_ldst;
      5'b11011:
        casez_tmp_84 = rob_uop_3_27_ldst;
      5'b11100:
        casez_tmp_84 = rob_uop_3_28_ldst;
      5'b11101:
        casez_tmp_84 = rob_uop_3_29_ldst;
      5'b11110:
        casez_tmp_84 = rob_uop_3_30_ldst;
      default:
        casez_tmp_84 = rob_uop_3_31_ldst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_85 = rob_uop_3_0_ldst_val;
      5'b00001:
        casez_tmp_85 = rob_uop_3_1_ldst_val;
      5'b00010:
        casez_tmp_85 = rob_uop_3_2_ldst_val;
      5'b00011:
        casez_tmp_85 = rob_uop_3_3_ldst_val;
      5'b00100:
        casez_tmp_85 = rob_uop_3_4_ldst_val;
      5'b00101:
        casez_tmp_85 = rob_uop_3_5_ldst_val;
      5'b00110:
        casez_tmp_85 = rob_uop_3_6_ldst_val;
      5'b00111:
        casez_tmp_85 = rob_uop_3_7_ldst_val;
      5'b01000:
        casez_tmp_85 = rob_uop_3_8_ldst_val;
      5'b01001:
        casez_tmp_85 = rob_uop_3_9_ldst_val;
      5'b01010:
        casez_tmp_85 = rob_uop_3_10_ldst_val;
      5'b01011:
        casez_tmp_85 = rob_uop_3_11_ldst_val;
      5'b01100:
        casez_tmp_85 = rob_uop_3_12_ldst_val;
      5'b01101:
        casez_tmp_85 = rob_uop_3_13_ldst_val;
      5'b01110:
        casez_tmp_85 = rob_uop_3_14_ldst_val;
      5'b01111:
        casez_tmp_85 = rob_uop_3_15_ldst_val;
      5'b10000:
        casez_tmp_85 = rob_uop_3_16_ldst_val;
      5'b10001:
        casez_tmp_85 = rob_uop_3_17_ldst_val;
      5'b10010:
        casez_tmp_85 = rob_uop_3_18_ldst_val;
      5'b10011:
        casez_tmp_85 = rob_uop_3_19_ldst_val;
      5'b10100:
        casez_tmp_85 = rob_uop_3_20_ldst_val;
      5'b10101:
        casez_tmp_85 = rob_uop_3_21_ldst_val;
      5'b10110:
        casez_tmp_85 = rob_uop_3_22_ldst_val;
      5'b10111:
        casez_tmp_85 = rob_uop_3_23_ldst_val;
      5'b11000:
        casez_tmp_85 = rob_uop_3_24_ldst_val;
      5'b11001:
        casez_tmp_85 = rob_uop_3_25_ldst_val;
      5'b11010:
        casez_tmp_85 = rob_uop_3_26_ldst_val;
      5'b11011:
        casez_tmp_85 = rob_uop_3_27_ldst_val;
      5'b11100:
        casez_tmp_85 = rob_uop_3_28_ldst_val;
      5'b11101:
        casez_tmp_85 = rob_uop_3_29_ldst_val;
      5'b11110:
        casez_tmp_85 = rob_uop_3_30_ldst_val;
      default:
        casez_tmp_85 = rob_uop_3_31_ldst_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_86 = rob_uop_3_0_dst_rtype;
      5'b00001:
        casez_tmp_86 = rob_uop_3_1_dst_rtype;
      5'b00010:
        casez_tmp_86 = rob_uop_3_2_dst_rtype;
      5'b00011:
        casez_tmp_86 = rob_uop_3_3_dst_rtype;
      5'b00100:
        casez_tmp_86 = rob_uop_3_4_dst_rtype;
      5'b00101:
        casez_tmp_86 = rob_uop_3_5_dst_rtype;
      5'b00110:
        casez_tmp_86 = rob_uop_3_6_dst_rtype;
      5'b00111:
        casez_tmp_86 = rob_uop_3_7_dst_rtype;
      5'b01000:
        casez_tmp_86 = rob_uop_3_8_dst_rtype;
      5'b01001:
        casez_tmp_86 = rob_uop_3_9_dst_rtype;
      5'b01010:
        casez_tmp_86 = rob_uop_3_10_dst_rtype;
      5'b01011:
        casez_tmp_86 = rob_uop_3_11_dst_rtype;
      5'b01100:
        casez_tmp_86 = rob_uop_3_12_dst_rtype;
      5'b01101:
        casez_tmp_86 = rob_uop_3_13_dst_rtype;
      5'b01110:
        casez_tmp_86 = rob_uop_3_14_dst_rtype;
      5'b01111:
        casez_tmp_86 = rob_uop_3_15_dst_rtype;
      5'b10000:
        casez_tmp_86 = rob_uop_3_16_dst_rtype;
      5'b10001:
        casez_tmp_86 = rob_uop_3_17_dst_rtype;
      5'b10010:
        casez_tmp_86 = rob_uop_3_18_dst_rtype;
      5'b10011:
        casez_tmp_86 = rob_uop_3_19_dst_rtype;
      5'b10100:
        casez_tmp_86 = rob_uop_3_20_dst_rtype;
      5'b10101:
        casez_tmp_86 = rob_uop_3_21_dst_rtype;
      5'b10110:
        casez_tmp_86 = rob_uop_3_22_dst_rtype;
      5'b10111:
        casez_tmp_86 = rob_uop_3_23_dst_rtype;
      5'b11000:
        casez_tmp_86 = rob_uop_3_24_dst_rtype;
      5'b11001:
        casez_tmp_86 = rob_uop_3_25_dst_rtype;
      5'b11010:
        casez_tmp_86 = rob_uop_3_26_dst_rtype;
      5'b11011:
        casez_tmp_86 = rob_uop_3_27_dst_rtype;
      5'b11100:
        casez_tmp_86 = rob_uop_3_28_dst_rtype;
      5'b11101:
        casez_tmp_86 = rob_uop_3_29_dst_rtype;
      5'b11110:
        casez_tmp_86 = rob_uop_3_30_dst_rtype;
      default:
        casez_tmp_86 = rob_uop_3_31_dst_rtype;
    endcase
  end // always @(*)
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_87 = rob_uop_3_0_fp_val;
      5'b00001:
        casez_tmp_87 = rob_uop_3_1_fp_val;
      5'b00010:
        casez_tmp_87 = rob_uop_3_2_fp_val;
      5'b00011:
        casez_tmp_87 = rob_uop_3_3_fp_val;
      5'b00100:
        casez_tmp_87 = rob_uop_3_4_fp_val;
      5'b00101:
        casez_tmp_87 = rob_uop_3_5_fp_val;
      5'b00110:
        casez_tmp_87 = rob_uop_3_6_fp_val;
      5'b00111:
        casez_tmp_87 = rob_uop_3_7_fp_val;
      5'b01000:
        casez_tmp_87 = rob_uop_3_8_fp_val;
      5'b01001:
        casez_tmp_87 = rob_uop_3_9_fp_val;
      5'b01010:
        casez_tmp_87 = rob_uop_3_10_fp_val;
      5'b01011:
        casez_tmp_87 = rob_uop_3_11_fp_val;
      5'b01100:
        casez_tmp_87 = rob_uop_3_12_fp_val;
      5'b01101:
        casez_tmp_87 = rob_uop_3_13_fp_val;
      5'b01110:
        casez_tmp_87 = rob_uop_3_14_fp_val;
      5'b01111:
        casez_tmp_87 = rob_uop_3_15_fp_val;
      5'b10000:
        casez_tmp_87 = rob_uop_3_16_fp_val;
      5'b10001:
        casez_tmp_87 = rob_uop_3_17_fp_val;
      5'b10010:
        casez_tmp_87 = rob_uop_3_18_fp_val;
      5'b10011:
        casez_tmp_87 = rob_uop_3_19_fp_val;
      5'b10100:
        casez_tmp_87 = rob_uop_3_20_fp_val;
      5'b10101:
        casez_tmp_87 = rob_uop_3_21_fp_val;
      5'b10110:
        casez_tmp_87 = rob_uop_3_22_fp_val;
      5'b10111:
        casez_tmp_87 = rob_uop_3_23_fp_val;
      5'b11000:
        casez_tmp_87 = rob_uop_3_24_fp_val;
      5'b11001:
        casez_tmp_87 = rob_uop_3_25_fp_val;
      5'b11010:
        casez_tmp_87 = rob_uop_3_26_fp_val;
      5'b11011:
        casez_tmp_87 = rob_uop_3_27_fp_val;
      5'b11100:
        casez_tmp_87 = rob_uop_3_28_fp_val;
      5'b11101:
        casez_tmp_87 = rob_uop_3_29_fp_val;
      5'b11110:
        casez_tmp_87 = rob_uop_3_30_fp_val;
      default:
        casez_tmp_87 = rob_uop_3_31_fp_val;
    endcase
  end // always @(*)
  wire        rbk_row_3 = _io_commit_rollback_T_3 & ~full;
  always @(*) begin
    casez (com_idx)
      5'b00000:
        casez_tmp_88 = rob_val_3_0;
      5'b00001:
        casez_tmp_88 = rob_val_3_1;
      5'b00010:
        casez_tmp_88 = rob_val_3_2;
      5'b00011:
        casez_tmp_88 = rob_val_3_3;
      5'b00100:
        casez_tmp_88 = rob_val_3_4;
      5'b00101:
        casez_tmp_88 = rob_val_3_5;
      5'b00110:
        casez_tmp_88 = rob_val_3_6;
      5'b00111:
        casez_tmp_88 = rob_val_3_7;
      5'b01000:
        casez_tmp_88 = rob_val_3_8;
      5'b01001:
        casez_tmp_88 = rob_val_3_9;
      5'b01010:
        casez_tmp_88 = rob_val_3_10;
      5'b01011:
        casez_tmp_88 = rob_val_3_11;
      5'b01100:
        casez_tmp_88 = rob_val_3_12;
      5'b01101:
        casez_tmp_88 = rob_val_3_13;
      5'b01110:
        casez_tmp_88 = rob_val_3_14;
      5'b01111:
        casez_tmp_88 = rob_val_3_15;
      5'b10000:
        casez_tmp_88 = rob_val_3_16;
      5'b10001:
        casez_tmp_88 = rob_val_3_17;
      5'b10010:
        casez_tmp_88 = rob_val_3_18;
      5'b10011:
        casez_tmp_88 = rob_val_3_19;
      5'b10100:
        casez_tmp_88 = rob_val_3_20;
      5'b10101:
        casez_tmp_88 = rob_val_3_21;
      5'b10110:
        casez_tmp_88 = rob_val_3_22;
      5'b10111:
        casez_tmp_88 = rob_val_3_23;
      5'b11000:
        casez_tmp_88 = rob_val_3_24;
      5'b11001:
        casez_tmp_88 = rob_val_3_25;
      5'b11010:
        casez_tmp_88 = rob_val_3_26;
      5'b11011:
        casez_tmp_88 = rob_val_3_27;
      5'b11100:
        casez_tmp_88 = rob_val_3_28;
      5'b11101:
        casez_tmp_88 = rob_val_3_29;
      5'b11110:
        casez_tmp_88 = rob_val_3_30;
      default:
        casez_tmp_88 = rob_val_3_31;
    endcase
  end // always @(*)
  wire        _io_commit_rbk_valids_3_output = rbk_row_3 & casez_tmp_88;
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_89 = rob_fflags_3_0;
      5'b00001:
        casez_tmp_89 = rob_fflags_3_1;
      5'b00010:
        casez_tmp_89 = rob_fflags_3_2;
      5'b00011:
        casez_tmp_89 = rob_fflags_3_3;
      5'b00100:
        casez_tmp_89 = rob_fflags_3_4;
      5'b00101:
        casez_tmp_89 = rob_fflags_3_5;
      5'b00110:
        casez_tmp_89 = rob_fflags_3_6;
      5'b00111:
        casez_tmp_89 = rob_fflags_3_7;
      5'b01000:
        casez_tmp_89 = rob_fflags_3_8;
      5'b01001:
        casez_tmp_89 = rob_fflags_3_9;
      5'b01010:
        casez_tmp_89 = rob_fflags_3_10;
      5'b01011:
        casez_tmp_89 = rob_fflags_3_11;
      5'b01100:
        casez_tmp_89 = rob_fflags_3_12;
      5'b01101:
        casez_tmp_89 = rob_fflags_3_13;
      5'b01110:
        casez_tmp_89 = rob_fflags_3_14;
      5'b01111:
        casez_tmp_89 = rob_fflags_3_15;
      5'b10000:
        casez_tmp_89 = rob_fflags_3_16;
      5'b10001:
        casez_tmp_89 = rob_fflags_3_17;
      5'b10010:
        casez_tmp_89 = rob_fflags_3_18;
      5'b10011:
        casez_tmp_89 = rob_fflags_3_19;
      5'b10100:
        casez_tmp_89 = rob_fflags_3_20;
      5'b10101:
        casez_tmp_89 = rob_fflags_3_21;
      5'b10110:
        casez_tmp_89 = rob_fflags_3_22;
      5'b10111:
        casez_tmp_89 = rob_fflags_3_23;
      5'b11000:
        casez_tmp_89 = rob_fflags_3_24;
      5'b11001:
        casez_tmp_89 = rob_fflags_3_25;
      5'b11010:
        casez_tmp_89 = rob_fflags_3_26;
      5'b11011:
        casez_tmp_89 = rob_fflags_3_27;
      5'b11100:
        casez_tmp_89 = rob_fflags_3_28;
      5'b11101:
        casez_tmp_89 = rob_fflags_3_29;
      5'b11110:
        casez_tmp_89 = rob_fflags_3_30;
      default:
        casez_tmp_89 = rob_fflags_3_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (rob_head)
      5'b00000:
        casez_tmp_90 = rob_uop_3_0_uses_ldq;
      5'b00001:
        casez_tmp_90 = rob_uop_3_1_uses_ldq;
      5'b00010:
        casez_tmp_90 = rob_uop_3_2_uses_ldq;
      5'b00011:
        casez_tmp_90 = rob_uop_3_3_uses_ldq;
      5'b00100:
        casez_tmp_90 = rob_uop_3_4_uses_ldq;
      5'b00101:
        casez_tmp_90 = rob_uop_3_5_uses_ldq;
      5'b00110:
        casez_tmp_90 = rob_uop_3_6_uses_ldq;
      5'b00111:
        casez_tmp_90 = rob_uop_3_7_uses_ldq;
      5'b01000:
        casez_tmp_90 = rob_uop_3_8_uses_ldq;
      5'b01001:
        casez_tmp_90 = rob_uop_3_9_uses_ldq;
      5'b01010:
        casez_tmp_90 = rob_uop_3_10_uses_ldq;
      5'b01011:
        casez_tmp_90 = rob_uop_3_11_uses_ldq;
      5'b01100:
        casez_tmp_90 = rob_uop_3_12_uses_ldq;
      5'b01101:
        casez_tmp_90 = rob_uop_3_13_uses_ldq;
      5'b01110:
        casez_tmp_90 = rob_uop_3_14_uses_ldq;
      5'b01111:
        casez_tmp_90 = rob_uop_3_15_uses_ldq;
      5'b10000:
        casez_tmp_90 = rob_uop_3_16_uses_ldq;
      5'b10001:
        casez_tmp_90 = rob_uop_3_17_uses_ldq;
      5'b10010:
        casez_tmp_90 = rob_uop_3_18_uses_ldq;
      5'b10011:
        casez_tmp_90 = rob_uop_3_19_uses_ldq;
      5'b10100:
        casez_tmp_90 = rob_uop_3_20_uses_ldq;
      5'b10101:
        casez_tmp_90 = rob_uop_3_21_uses_ldq;
      5'b10110:
        casez_tmp_90 = rob_uop_3_22_uses_ldq;
      5'b10111:
        casez_tmp_90 = rob_uop_3_23_uses_ldq;
      5'b11000:
        casez_tmp_90 = rob_uop_3_24_uses_ldq;
      5'b11001:
        casez_tmp_90 = rob_uop_3_25_uses_ldq;
      5'b11010:
        casez_tmp_90 = rob_uop_3_26_uses_ldq;
      5'b11011:
        casez_tmp_90 = rob_uop_3_27_uses_ldq;
      5'b11100:
        casez_tmp_90 = rob_uop_3_28_uses_ldq;
      5'b11101:
        casez_tmp_90 = rob_uop_3_29_uses_ldq;
      5'b11110:
        casez_tmp_90 = rob_uop_3_30_uses_ldq;
      default:
        casez_tmp_90 = rob_uop_3_31_uses_ldq;
    endcase
  end // always @(*)
  reg         block_commit_REG_1;
  wire        exception_thrown = can_throw_exception_3 & ~_GEN_1 & ~_io_commit_valids_2_output | can_throw_exception_2 & ~_GEN_0 & ~_io_commit_valids_1_output | can_throw_exception_1 & ~_GEN & ~_io_commit_valids_0_output | can_throw_exception_0 & ~block_commit;
  wire        is_mini_exception = r_xcpt_uop_exc_cause == 64'h10 | r_xcpt_uop_exc_cause == 64'h11;
  wire [5:0]  com_xcpt_uop_ftq_idx = casez_tmp ? casez_tmp_14 : casez_tmp_2 ? casez_tmp_34 : casez_tmp_5 ? casez_tmp_54 : casez_tmp_74;
  wire        com_xcpt_uop_edge_inst = casez_tmp ? casez_tmp_15 : casez_tmp_2 ? casez_tmp_35 : casez_tmp_5 ? casez_tmp_55 : casez_tmp_75;
  wire [5:0]  com_xcpt_uop_pc_lob = casez_tmp ? casez_tmp_16 : casez_tmp_2 ? casez_tmp_36 : casez_tmp_5 ? casez_tmp_56 : casez_tmp_76;
  wire        flush_commit_mask_0 = _io_commit_valids_0_output & casez_tmp_23;
  wire        flush_commit_mask_1 = _io_commit_valids_1_output & casez_tmp_43;
  wire        flush_commit_mask_2 = _io_commit_valids_2_output & casez_tmp_63;
  wire        flush_commit_mask_3 = _io_commit_valids_3_output & casez_tmp_83;
  wire        flush_commit = flush_commit_mask_0 | flush_commit_mask_1 | flush_commit_mask_2 | flush_commit_mask_3;
  wire        _io_flush_valid_output = exception_thrown | flush_commit;
  wire        _fflags_val_0_T = _io_commit_valids_0_output & casez_tmp_27;
  wire        fflags_val_0 = _fflags_val_0_T & ~casez_tmp_21;
  wire        _fflags_val_1_T = _io_commit_valids_1_output & casez_tmp_47;
  wire        fflags_val_1 = _fflags_val_1_T & ~casez_tmp_41;
  wire        _fflags_val_2_T = _io_commit_valids_2_output & casez_tmp_67;
  wire        fflags_val_2 = _fflags_val_2_T & ~casez_tmp_61;
  wire        _fflags_val_3_T = _io_commit_valids_3_output & casez_tmp_87;
  wire        fflags_val_3 = _fflags_val_3_T & ~casez_tmp_81;
  wire        enq_xcpts_0 = io_enq_valids_0 & io_enq_uops_0_exception;
  wire        enq_xcpts_1 = io_enq_valids_1 & io_enq_uops_1_exception;
  wire        enq_xcpts_2 = io_enq_valids_2 & io_enq_uops_2_exception;
  wire [1:0]  idx = enq_xcpts_0 ? 2'h0 : enq_xcpts_1 ? 2'h1 : {1'h1, ~enq_xcpts_2};
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_91 = io_enq_uops_0_br_mask;
      2'b01:
        casez_tmp_91 = io_enq_uops_1_br_mask;
      2'b10:
        casez_tmp_91 = io_enq_uops_2_br_mask;
      default:
        casez_tmp_91 = io_enq_uops_3_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_92 = io_enq_uops_0_pc_lob;
      2'b01:
        casez_tmp_92 = io_enq_uops_1_pc_lob;
      2'b10:
        casez_tmp_92 = io_enq_uops_2_pc_lob;
      default:
        casez_tmp_92 = io_enq_uops_3_pc_lob;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_93 = io_enq_uops_0_rob_idx;
      2'b01:
        casez_tmp_93 = io_enq_uops_1_rob_idx;
      2'b10:
        casez_tmp_93 = io_enq_uops_2_rob_idx;
      default:
        casez_tmp_93 = io_enq_uops_3_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (idx)
      2'b00:
        casez_tmp_94 = io_enq_uops_0_exc_cause;
      2'b01:
        casez_tmp_94 = io_enq_uops_1_exc_cause;
      2'b10:
        casez_tmp_94 = io_enq_uops_2_exc_cause;
      default:
        casez_tmp_94 = io_enq_uops_3_exc_cause;
    endcase
  end // always @(*)
  wire        _finished_committing_row_T_7 = rob_head == rob_tail;
  wire        empty = _finished_committing_row_T_7 & {casez_tmp_8, casez_tmp_5, casez_tmp_2, casez_tmp} == 4'h0;
  reg         r_partial_row;
  wire        finished_committing_row = (|{_io_commit_valids_3_output, _io_commit_valids_2_output, _io_commit_valids_1_output, _io_commit_valids_0_output}) & ({_io_commit_valids_3_output, _io_commit_valids_2_output, _io_commit_valids_1_output, _io_commit_valids_0_output} ^ {casez_tmp_8, casez_tmp_5, casez_tmp_2, casez_tmp}) == 4'h0 & ~(r_partial_row & _finished_committing_row_T_7 & ~maybe_full);
  wire        _io_ready_T = rob_state == 2'h1;
  wire [3:0]  _GEN_2284 = {io_enq_valids_3, io_enq_valids_2, io_enq_valids_1, io_enq_valids_0};
  wire        _GEN_2285 = _io_commit_rollback_T_3 & (rob_tail != rob_head | maybe_full);
  wire        rob_deq = _GEN_2285 | finished_committing_row;
  reg         REG;
  reg         REG_1;
  reg         REG_2;
  wire [1:0]  _GEN_54139 = empty ? 2'h1 : rob_state;
  always @(*) begin
    casez (rob_state)
      2'b00:
        casez_tmp_95 = 2'h1;
      2'b01:
        casez_tmp_95 = REG_1 ? 2'h2 : io_enq_valids_3 & io_enq_uops_3_is_unique | io_enq_valids_2 & io_enq_uops_2_is_unique | io_enq_valids_1 & io_enq_uops_1_is_unique | io_enq_valids_0 & io_enq_uops_0_is_unique ? 2'h3 : rob_state;
      2'b10:
        casez_tmp_95 = _GEN_54139;
      default:
        casez_tmp_95 = REG_2 ? 2'h2 : _GEN_54139;
    endcase
  end // always @(*)
  always @(*) begin
    casez (casez_tmp ? 2'h0 : casez_tmp_2 ? 2'h1 : {1'h1, ~casez_tmp_5})
      2'b00:
        casez_tmp_96 = casez_tmp_30;
      2'b01:
        casez_tmp_96 = casez_tmp_50;
      2'b10:
        casez_tmp_96 = casez_tmp_70;
      default:
        casez_tmp_96 = casez_tmp_90;
    endcase
  end // always @(*)
  reg         io_com_load_is_at_rob_head_REG;
  wire [2:0]  _rob_head_lsb_T_8 = casez_tmp ? 3'h0 : casez_tmp_2 ? 3'h1 : casez_tmp_5 ? 3'h2 : {casez_tmp_8, 2'h0};
  wire [2:0]  _GEN_2286 = {io_enq_valids_2, io_enq_valids_1, io_enq_valids_0} | {io_enq_valids_3, io_enq_valids_2, io_enq_valids_1};
  wire [1:0]  _GEN_2287 = _GEN_2286[1:0] | {io_enq_valids_3, io_enq_valids_2};
  wire [2:0]  _rob_tail_lsb_T_8 = ~{_GEN_2286[2], _GEN_2287[1], _GEN_2287[0] | io_enq_valids_3};
  wire        _GEN_2288 = rob_head == 5'h1;
  wire        _GEN_2289 = rob_head == 5'h2;
  wire        _GEN_2290 = rob_head == 5'h3;
  wire        _GEN_2291 = rob_head == 5'h4;
  wire        _GEN_2292 = rob_head == 5'h5;
  wire        _GEN_2293 = rob_head == 5'h6;
  wire        _GEN_2294 = rob_head == 5'h7;
  wire        _GEN_2295 = rob_head == 5'h8;
  wire        _GEN_2296 = rob_head == 5'h9;
  wire        _GEN_2297 = rob_head == 5'hA;
  wire        _GEN_2298 = rob_head == 5'hB;
  wire        _GEN_2299 = rob_head == 5'hC;
  wire        _GEN_2300 = rob_head == 5'hD;
  wire        _GEN_2301 = rob_head == 5'hE;
  wire        _GEN_2302 = rob_head == 5'hF;
  wire        _GEN_2303 = rob_head == 5'h10;
  wire        _GEN_2304 = rob_head == 5'h11;
  wire        _GEN_2305 = rob_head == 5'h12;
  wire        _GEN_2306 = rob_head == 5'h13;
  wire        _GEN_2307 = rob_head == 5'h14;
  wire        _GEN_2308 = rob_head == 5'h15;
  wire        _GEN_2309 = rob_head == 5'h16;
  wire        _GEN_2310 = rob_head == 5'h17;
  wire        _GEN_2311 = rob_head == 5'h18;
  wire        _GEN_2312 = rob_head == 5'h19;
  wire        _GEN_2313 = rob_head == 5'h1A;
  wire        _GEN_2314 = rob_head == 5'h1B;
  wire        _GEN_2315 = rob_head == 5'h1C;
  wire        _GEN_2316 = rob_head == 5'h1D;
  wire        _GEN_2317 = rob_head == 5'h1E;
  wire        _GEN_2828 = _GEN_33 | rob_val__0;
  wire        _GEN_2829 = _GEN_34 | rob_val__1;
  wire        _GEN_2830 = _GEN_35 | rob_val__2;
  wire        _GEN_2831 = _GEN_36 | rob_val__3;
  wire        _GEN_2832 = _GEN_37 | rob_val__4;
  wire        _GEN_2833 = _GEN_38 | rob_val__5;
  wire        _GEN_2834 = _GEN_39 | rob_val__6;
  wire        _GEN_2835 = _GEN_40 | rob_val__7;
  wire        _GEN_2836 = _GEN_41 | rob_val__8;
  wire        _GEN_2837 = _GEN_42 | rob_val__9;
  wire        _GEN_2838 = _GEN_43 | rob_val__10;
  wire        _GEN_2839 = _GEN_44 | rob_val__11;
  wire        _GEN_2840 = _GEN_45 | rob_val__12;
  wire        _GEN_2841 = _GEN_46 | rob_val__13;
  wire        _GEN_2842 = _GEN_47 | rob_val__14;
  wire        _GEN_2843 = _GEN_48 | rob_val__15;
  wire        _GEN_2844 = _GEN_49 | rob_val__16;
  wire        _GEN_2845 = _GEN_50 | rob_val__17;
  wire        _GEN_2846 = _GEN_51 | rob_val__18;
  wire        _GEN_2847 = _GEN_52 | rob_val__19;
  wire        _GEN_2848 = _GEN_53 | rob_val__20;
  wire        _GEN_2849 = _GEN_54 | rob_val__21;
  wire        _GEN_2850 = _GEN_55 | rob_val__22;
  wire        _GEN_2851 = _GEN_56 | rob_val__23;
  wire        _GEN_2852 = _GEN_57 | rob_val__24;
  wire        _GEN_2853 = _GEN_58 | rob_val__25;
  wire        _GEN_2854 = _GEN_59 | rob_val__26;
  wire        _GEN_2855 = _GEN_60 | rob_val__27;
  wire        _GEN_2856 = _GEN_61 | rob_val__28;
  wire        _GEN_2857 = _GEN_62 | rob_val__29;
  wire        _GEN_2858 = _GEN_63 | rob_val__30;
  wire        _GEN_2859 = _GEN_64 | rob_val__31;
  wire        _GEN_2318 = rob_head == 5'h0;
  wire        _GEN_16192 = _GEN_898 | rob_val_1_0;
  wire        _GEN_16193 = _GEN_899 | rob_val_1_1;
  wire        _GEN_16194 = _GEN_900 | rob_val_1_2;
  wire        _GEN_16195 = _GEN_901 | rob_val_1_3;
  wire        _GEN_16196 = _GEN_902 | rob_val_1_4;
  wire        _GEN_16197 = _GEN_903 | rob_val_1_5;
  wire        _GEN_16198 = _GEN_904 | rob_val_1_6;
  wire        _GEN_16199 = _GEN_905 | rob_val_1_7;
  wire        _GEN_16200 = _GEN_906 | rob_val_1_8;
  wire        _GEN_16201 = _GEN_907 | rob_val_1_9;
  wire        _GEN_16202 = _GEN_908 | rob_val_1_10;
  wire        _GEN_16203 = _GEN_909 | rob_val_1_11;
  wire        _GEN_16204 = _GEN_910 | rob_val_1_12;
  wire        _GEN_16205 = _GEN_911 | rob_val_1_13;
  wire        _GEN_16206 = _GEN_912 | rob_val_1_14;
  wire        _GEN_16207 = _GEN_913 | rob_val_1_15;
  wire        _GEN_16208 = _GEN_914 | rob_val_1_16;
  wire        _GEN_16209 = _GEN_915 | rob_val_1_17;
  wire        _GEN_16210 = _GEN_916 | rob_val_1_18;
  wire        _GEN_16211 = _GEN_917 | rob_val_1_19;
  wire        _GEN_16212 = _GEN_918 | rob_val_1_20;
  wire        _GEN_16213 = _GEN_919 | rob_val_1_21;
  wire        _GEN_16214 = _GEN_920 | rob_val_1_22;
  wire        _GEN_16215 = _GEN_921 | rob_val_1_23;
  wire        _GEN_16216 = _GEN_922 | rob_val_1_24;
  wire        _GEN_16217 = _GEN_923 | rob_val_1_25;
  wire        _GEN_16218 = _GEN_924 | rob_val_1_26;
  wire        _GEN_16219 = _GEN_925 | rob_val_1_27;
  wire        _GEN_16220 = _GEN_926 | rob_val_1_28;
  wire        _GEN_16221 = _GEN_927 | rob_val_1_29;
  wire        _GEN_16222 = _GEN_928 | rob_val_1_30;
  wire        _GEN_16223 = _GEN_929 | rob_val_1_31;
  wire        _GEN_29556 = _GEN_1360 | rob_val_2_0;
  wire        _GEN_29557 = _GEN_1361 | rob_val_2_1;
  wire        _GEN_29558 = _GEN_1362 | rob_val_2_2;
  wire        _GEN_29559 = _GEN_1363 | rob_val_2_3;
  wire        _GEN_29560 = _GEN_1364 | rob_val_2_4;
  wire        _GEN_29561 = _GEN_1365 | rob_val_2_5;
  wire        _GEN_29562 = _GEN_1366 | rob_val_2_6;
  wire        _GEN_29563 = _GEN_1367 | rob_val_2_7;
  wire        _GEN_29564 = _GEN_1368 | rob_val_2_8;
  wire        _GEN_29565 = _GEN_1369 | rob_val_2_9;
  wire        _GEN_29566 = _GEN_1370 | rob_val_2_10;
  wire        _GEN_29567 = _GEN_1371 | rob_val_2_11;
  wire        _GEN_29568 = _GEN_1372 | rob_val_2_12;
  wire        _GEN_29569 = _GEN_1373 | rob_val_2_13;
  wire        _GEN_29570 = _GEN_1374 | rob_val_2_14;
  wire        _GEN_29571 = _GEN_1375 | rob_val_2_15;
  wire        _GEN_29572 = _GEN_1376 | rob_val_2_16;
  wire        _GEN_29573 = _GEN_1377 | rob_val_2_17;
  wire        _GEN_29574 = _GEN_1378 | rob_val_2_18;
  wire        _GEN_29575 = _GEN_1379 | rob_val_2_19;
  wire        _GEN_29576 = _GEN_1380 | rob_val_2_20;
  wire        _GEN_29577 = _GEN_1381 | rob_val_2_21;
  wire        _GEN_29578 = _GEN_1382 | rob_val_2_22;
  wire        _GEN_29579 = _GEN_1383 | rob_val_2_23;
  wire        _GEN_29580 = _GEN_1384 | rob_val_2_24;
  wire        _GEN_29581 = _GEN_1385 | rob_val_2_25;
  wire        _GEN_29582 = _GEN_1386 | rob_val_2_26;
  wire        _GEN_29583 = _GEN_1387 | rob_val_2_27;
  wire        _GEN_29584 = _GEN_1388 | rob_val_2_28;
  wire        _GEN_29585 = _GEN_1389 | rob_val_2_29;
  wire        _GEN_29586 = _GEN_1390 | rob_val_2_30;
  wire        _GEN_29587 = _GEN_1391 | rob_val_2_31;
  wire        _GEN_42920 = _GEN_1822 | rob_val_3_0;
  wire        _GEN_42921 = _GEN_1823 | rob_val_3_1;
  wire        _GEN_42922 = _GEN_1824 | rob_val_3_2;
  wire        _GEN_42923 = _GEN_1825 | rob_val_3_3;
  wire        _GEN_42924 = _GEN_1826 | rob_val_3_4;
  wire        _GEN_42925 = _GEN_1827 | rob_val_3_5;
  wire        _GEN_42926 = _GEN_1828 | rob_val_3_6;
  wire        _GEN_42927 = _GEN_1829 | rob_val_3_7;
  wire        _GEN_42928 = _GEN_1830 | rob_val_3_8;
  wire        _GEN_42929 = _GEN_1831 | rob_val_3_9;
  wire        _GEN_42930 = _GEN_1832 | rob_val_3_10;
  wire        _GEN_42931 = _GEN_1833 | rob_val_3_11;
  wire        _GEN_42932 = _GEN_1834 | rob_val_3_12;
  wire        _GEN_42933 = _GEN_1835 | rob_val_3_13;
  wire        _GEN_42934 = _GEN_1836 | rob_val_3_14;
  wire        _GEN_42935 = _GEN_1837 | rob_val_3_15;
  wire        _GEN_42936 = _GEN_1838 | rob_val_3_16;
  wire        _GEN_42937 = _GEN_1839 | rob_val_3_17;
  wire        _GEN_42938 = _GEN_1840 | rob_val_3_18;
  wire        _GEN_42939 = _GEN_1841 | rob_val_3_19;
  wire        _GEN_42940 = _GEN_1842 | rob_val_3_20;
  wire        _GEN_42941 = _GEN_1843 | rob_val_3_21;
  wire        _GEN_42942 = _GEN_1844 | rob_val_3_22;
  wire        _GEN_42943 = _GEN_1845 | rob_val_3_23;
  wire        _GEN_42944 = _GEN_1846 | rob_val_3_24;
  wire        _GEN_42945 = _GEN_1847 | rob_val_3_25;
  wire        _GEN_42946 = _GEN_1848 | rob_val_3_26;
  wire        _GEN_42947 = _GEN_1849 | rob_val_3_27;
  wire        _GEN_42948 = _GEN_1850 | rob_val_3_28;
  wire        _GEN_42949 = _GEN_1851 | rob_val_3_29;
  wire        _GEN_42950 = _GEN_1852 | rob_val_3_30;
  wire        _GEN_42951 = _GEN_1853 | rob_val_3_31;
  wire        _GEN_2319 = _io_commit_rollback_T_3 & _full_T & ~maybe_full;
  wire        _GEN_54123 = (|_GEN_2284) & ~io_enq_partial_stall;
  wire        _rob_bsy_T = io_enq_uops_0_is_fence | io_enq_uops_0_is_fencei;
  wire        _GEN_2860 = _GEN_33 ? ~_rob_bsy_T : rob_bsy__0;
  wire        _GEN_2861 = _GEN_34 ? ~_rob_bsy_T : rob_bsy__1;
  wire        _GEN_2862 = _GEN_35 ? ~_rob_bsy_T : rob_bsy__2;
  wire        _GEN_2863 = _GEN_36 ? ~_rob_bsy_T : rob_bsy__3;
  wire        _GEN_2864 = _GEN_37 ? ~_rob_bsy_T : rob_bsy__4;
  wire        _GEN_2865 = _GEN_38 ? ~_rob_bsy_T : rob_bsy__5;
  wire        _GEN_2866 = _GEN_39 ? ~_rob_bsy_T : rob_bsy__6;
  wire        _GEN_2867 = _GEN_40 ? ~_rob_bsy_T : rob_bsy__7;
  wire        _GEN_2868 = _GEN_41 ? ~_rob_bsy_T : rob_bsy__8;
  wire        _GEN_2869 = _GEN_42 ? ~_rob_bsy_T : rob_bsy__9;
  wire        _GEN_2870 = _GEN_43 ? ~_rob_bsy_T : rob_bsy__10;
  wire        _GEN_2871 = _GEN_44 ? ~_rob_bsy_T : rob_bsy__11;
  wire        _GEN_2872 = _GEN_45 ? ~_rob_bsy_T : rob_bsy__12;
  wire        _GEN_2873 = _GEN_46 ? ~_rob_bsy_T : rob_bsy__13;
  wire        _GEN_2874 = _GEN_47 ? ~_rob_bsy_T : rob_bsy__14;
  wire        _GEN_2875 = _GEN_48 ? ~_rob_bsy_T : rob_bsy__15;
  wire        _GEN_2876 = _GEN_49 ? ~_rob_bsy_T : rob_bsy__16;
  wire        _GEN_2877 = _GEN_50 ? ~_rob_bsy_T : rob_bsy__17;
  wire        _GEN_2878 = _GEN_51 ? ~_rob_bsy_T : rob_bsy__18;
  wire        _GEN_2879 = _GEN_52 ? ~_rob_bsy_T : rob_bsy__19;
  wire        _GEN_2880 = _GEN_53 ? ~_rob_bsy_T : rob_bsy__20;
  wire        _GEN_2881 = _GEN_54 ? ~_rob_bsy_T : rob_bsy__21;
  wire        _GEN_2882 = _GEN_55 ? ~_rob_bsy_T : rob_bsy__22;
  wire        _GEN_2883 = _GEN_56 ? ~_rob_bsy_T : rob_bsy__23;
  wire        _GEN_2884 = _GEN_57 ? ~_rob_bsy_T : rob_bsy__24;
  wire        _GEN_2885 = _GEN_58 ? ~_rob_bsy_T : rob_bsy__25;
  wire        _GEN_2886 = _GEN_59 ? ~_rob_bsy_T : rob_bsy__26;
  wire        _GEN_2887 = _GEN_60 ? ~_rob_bsy_T : rob_bsy__27;
  wire        _GEN_2888 = _GEN_61 ? ~_rob_bsy_T : rob_bsy__28;
  wire        _GEN_2889 = _GEN_62 ? ~_rob_bsy_T : rob_bsy__29;
  wire        _GEN_2890 = _GEN_63 ? ~_rob_bsy_T : rob_bsy__30;
  wire        _GEN_2891 = _GEN_64 ? ~_rob_bsy_T : rob_bsy__31;
  wire        _GEN_5836 = _GEN_129 ? ~_GEN_131 & _GEN_2860 : ~_GEN_97 & _GEN_2860;
  wire        _GEN_5837 = _GEN_129 ? ~_GEN_133 & _GEN_2861 : ~_GEN_98 & _GEN_2861;
  wire        _GEN_5838 = _GEN_129 ? ~_GEN_135 & _GEN_2862 : ~_GEN_99 & _GEN_2862;
  wire        _GEN_5839 = _GEN_129 ? ~_GEN_137 & _GEN_2863 : ~_GEN_100 & _GEN_2863;
  wire        _GEN_5840 = _GEN_129 ? ~_GEN_139 & _GEN_2864 : ~_GEN_101 & _GEN_2864;
  wire        _GEN_5841 = _GEN_129 ? ~_GEN_141 & _GEN_2865 : ~_GEN_102 & _GEN_2865;
  wire        _GEN_5842 = _GEN_129 ? ~_GEN_143 & _GEN_2866 : ~_GEN_103 & _GEN_2866;
  wire        _GEN_5843 = _GEN_129 ? ~_GEN_145 & _GEN_2867 : ~_GEN_104 & _GEN_2867;
  wire        _GEN_5844 = _GEN_129 ? ~_GEN_147 & _GEN_2868 : ~_GEN_105 & _GEN_2868;
  wire        _GEN_5845 = _GEN_129 ? ~_GEN_149 & _GEN_2869 : ~_GEN_106 & _GEN_2869;
  wire        _GEN_5846 = _GEN_129 ? ~_GEN_151 & _GEN_2870 : ~_GEN_107 & _GEN_2870;
  wire        _GEN_5847 = _GEN_129 ? ~_GEN_153 & _GEN_2871 : ~_GEN_108 & _GEN_2871;
  wire        _GEN_5848 = _GEN_129 ? ~_GEN_155 & _GEN_2872 : ~_GEN_109 & _GEN_2872;
  wire        _GEN_5849 = _GEN_129 ? ~_GEN_157 & _GEN_2873 : ~_GEN_110 & _GEN_2873;
  wire        _GEN_5850 = _GEN_129 ? ~_GEN_159 & _GEN_2874 : ~_GEN_111 & _GEN_2874;
  wire        _GEN_5851 = _GEN_129 ? ~_GEN_161 & _GEN_2875 : ~_GEN_112 & _GEN_2875;
  wire        _GEN_5852 = _GEN_129 ? ~_GEN_163 & _GEN_2876 : ~_GEN_113 & _GEN_2876;
  wire        _GEN_5853 = _GEN_129 ? ~_GEN_165 & _GEN_2877 : ~_GEN_114 & _GEN_2877;
  wire        _GEN_5854 = _GEN_129 ? ~_GEN_167 & _GEN_2878 : ~_GEN_115 & _GEN_2878;
  wire        _GEN_5855 = _GEN_129 ? ~_GEN_169 & _GEN_2879 : ~_GEN_116 & _GEN_2879;
  wire        _GEN_5856 = _GEN_129 ? ~_GEN_171 & _GEN_2880 : ~_GEN_117 & _GEN_2880;
  wire        _GEN_5857 = _GEN_129 ? ~_GEN_173 & _GEN_2881 : ~_GEN_118 & _GEN_2881;
  wire        _GEN_5858 = _GEN_129 ? ~_GEN_175 & _GEN_2882 : ~_GEN_119 & _GEN_2882;
  wire        _GEN_5859 = _GEN_129 ? ~_GEN_177 & _GEN_2883 : ~_GEN_120 & _GEN_2883;
  wire        _GEN_5860 = _GEN_129 ? ~_GEN_179 & _GEN_2884 : ~_GEN_121 & _GEN_2884;
  wire        _GEN_5861 = _GEN_129 ? ~_GEN_181 & _GEN_2885 : ~_GEN_122 & _GEN_2885;
  wire        _GEN_5862 = _GEN_129 ? ~_GEN_183 & _GEN_2886 : ~_GEN_123 & _GEN_2886;
  wire        _GEN_5863 = _GEN_129 ? ~_GEN_185 & _GEN_2887 : ~_GEN_124 & _GEN_2887;
  wire        _GEN_5864 = _GEN_129 ? ~_GEN_187 & _GEN_2888 : ~_GEN_125 & _GEN_2888;
  wire        _GEN_5865 = _GEN_129 ? ~_GEN_189 & _GEN_2889 : ~_GEN_126 & _GEN_2889;
  wire        _GEN_5866 = _GEN_129 ? ~_GEN_191 & _GEN_2890 : ~_GEN_127 & _GEN_2890;
  wire        _GEN_5867 = _GEN_129 ? ~_GEN_192 & _GEN_2891 : ~_GEN_128 & _GEN_2891;
  wire        _GEN_6220 = _GEN_257 ? ~_GEN_259 & _GEN_5836 : ~_GEN_225 & _GEN_5836;
  wire        _GEN_6221 = _GEN_257 ? ~_GEN_261 & _GEN_5837 : ~_GEN_226 & _GEN_5837;
  wire        _GEN_6222 = _GEN_257 ? ~_GEN_263 & _GEN_5838 : ~_GEN_227 & _GEN_5838;
  wire        _GEN_6223 = _GEN_257 ? ~_GEN_265 & _GEN_5839 : ~_GEN_228 & _GEN_5839;
  wire        _GEN_6224 = _GEN_257 ? ~_GEN_267 & _GEN_5840 : ~_GEN_229 & _GEN_5840;
  wire        _GEN_6225 = _GEN_257 ? ~_GEN_269 & _GEN_5841 : ~_GEN_230 & _GEN_5841;
  wire        _GEN_6226 = _GEN_257 ? ~_GEN_271 & _GEN_5842 : ~_GEN_231 & _GEN_5842;
  wire        _GEN_6227 = _GEN_257 ? ~_GEN_273 & _GEN_5843 : ~_GEN_232 & _GEN_5843;
  wire        _GEN_6228 = _GEN_257 ? ~_GEN_275 & _GEN_5844 : ~_GEN_233 & _GEN_5844;
  wire        _GEN_6229 = _GEN_257 ? ~_GEN_277 & _GEN_5845 : ~_GEN_234 & _GEN_5845;
  wire        _GEN_6230 = _GEN_257 ? ~_GEN_279 & _GEN_5846 : ~_GEN_235 & _GEN_5846;
  wire        _GEN_6231 = _GEN_257 ? ~_GEN_281 & _GEN_5847 : ~_GEN_236 & _GEN_5847;
  wire        _GEN_6232 = _GEN_257 ? ~_GEN_283 & _GEN_5848 : ~_GEN_237 & _GEN_5848;
  wire        _GEN_6233 = _GEN_257 ? ~_GEN_285 & _GEN_5849 : ~_GEN_238 & _GEN_5849;
  wire        _GEN_6234 = _GEN_257 ? ~_GEN_287 & _GEN_5850 : ~_GEN_239 & _GEN_5850;
  wire        _GEN_6235 = _GEN_257 ? ~_GEN_289 & _GEN_5851 : ~_GEN_240 & _GEN_5851;
  wire        _GEN_6236 = _GEN_257 ? ~_GEN_291 & _GEN_5852 : ~_GEN_241 & _GEN_5852;
  wire        _GEN_6237 = _GEN_257 ? ~_GEN_293 & _GEN_5853 : ~_GEN_242 & _GEN_5853;
  wire        _GEN_6238 = _GEN_257 ? ~_GEN_295 & _GEN_5854 : ~_GEN_243 & _GEN_5854;
  wire        _GEN_6239 = _GEN_257 ? ~_GEN_297 & _GEN_5855 : ~_GEN_244 & _GEN_5855;
  wire        _GEN_6240 = _GEN_257 ? ~_GEN_299 & _GEN_5856 : ~_GEN_245 & _GEN_5856;
  wire        _GEN_6241 = _GEN_257 ? ~_GEN_301 & _GEN_5857 : ~_GEN_246 & _GEN_5857;
  wire        _GEN_6242 = _GEN_257 ? ~_GEN_303 & _GEN_5858 : ~_GEN_247 & _GEN_5858;
  wire        _GEN_6243 = _GEN_257 ? ~_GEN_305 & _GEN_5859 : ~_GEN_248 & _GEN_5859;
  wire        _GEN_6244 = _GEN_257 ? ~_GEN_307 & _GEN_5860 : ~_GEN_249 & _GEN_5860;
  wire        _GEN_6245 = _GEN_257 ? ~_GEN_309 & _GEN_5861 : ~_GEN_250 & _GEN_5861;
  wire        _GEN_6246 = _GEN_257 ? ~_GEN_311 & _GEN_5862 : ~_GEN_251 & _GEN_5862;
  wire        _GEN_6247 = _GEN_257 ? ~_GEN_313 & _GEN_5863 : ~_GEN_252 & _GEN_5863;
  wire        _GEN_6248 = _GEN_257 ? ~_GEN_315 & _GEN_5864 : ~_GEN_253 & _GEN_5864;
  wire        _GEN_6249 = _GEN_257 ? ~_GEN_317 & _GEN_5865 : ~_GEN_254 & _GEN_5865;
  wire        _GEN_6250 = _GEN_257 ? ~_GEN_319 & _GEN_5866 : ~_GEN_255 & _GEN_5866;
  wire        _GEN_6251 = _GEN_257 ? ~_GEN_320 & _GEN_5867 : ~_GEN_256 & _GEN_5867;
  wire        _GEN_6604 = _GEN_385 ? ~_GEN_387 & _GEN_6220 : ~_GEN_353 & _GEN_6220;
  wire        _GEN_6605 = _GEN_385 ? ~_GEN_389 & _GEN_6221 : ~_GEN_354 & _GEN_6221;
  wire        _GEN_6606 = _GEN_385 ? ~_GEN_391 & _GEN_6222 : ~_GEN_355 & _GEN_6222;
  wire        _GEN_6607 = _GEN_385 ? ~_GEN_393 & _GEN_6223 : ~_GEN_356 & _GEN_6223;
  wire        _GEN_6608 = _GEN_385 ? ~_GEN_395 & _GEN_6224 : ~_GEN_357 & _GEN_6224;
  wire        _GEN_6609 = _GEN_385 ? ~_GEN_397 & _GEN_6225 : ~_GEN_358 & _GEN_6225;
  wire        _GEN_6610 = _GEN_385 ? ~_GEN_399 & _GEN_6226 : ~_GEN_359 & _GEN_6226;
  wire        _GEN_6611 = _GEN_385 ? ~_GEN_401 & _GEN_6227 : ~_GEN_360 & _GEN_6227;
  wire        _GEN_6612 = _GEN_385 ? ~_GEN_403 & _GEN_6228 : ~_GEN_361 & _GEN_6228;
  wire        _GEN_6613 = _GEN_385 ? ~_GEN_405 & _GEN_6229 : ~_GEN_362 & _GEN_6229;
  wire        _GEN_6614 = _GEN_385 ? ~_GEN_407 & _GEN_6230 : ~_GEN_363 & _GEN_6230;
  wire        _GEN_6615 = _GEN_385 ? ~_GEN_409 & _GEN_6231 : ~_GEN_364 & _GEN_6231;
  wire        _GEN_6616 = _GEN_385 ? ~_GEN_411 & _GEN_6232 : ~_GEN_365 & _GEN_6232;
  wire        _GEN_6617 = _GEN_385 ? ~_GEN_413 & _GEN_6233 : ~_GEN_366 & _GEN_6233;
  wire        _GEN_6618 = _GEN_385 ? ~_GEN_415 & _GEN_6234 : ~_GEN_367 & _GEN_6234;
  wire        _GEN_6619 = _GEN_385 ? ~_GEN_417 & _GEN_6235 : ~_GEN_368 & _GEN_6235;
  wire        _GEN_6620 = _GEN_385 ? ~_GEN_419 & _GEN_6236 : ~_GEN_369 & _GEN_6236;
  wire        _GEN_6621 = _GEN_385 ? ~_GEN_421 & _GEN_6237 : ~_GEN_370 & _GEN_6237;
  wire        _GEN_6622 = _GEN_385 ? ~_GEN_423 & _GEN_6238 : ~_GEN_371 & _GEN_6238;
  wire        _GEN_6623 = _GEN_385 ? ~_GEN_425 & _GEN_6239 : ~_GEN_372 & _GEN_6239;
  wire        _GEN_6624 = _GEN_385 ? ~_GEN_427 & _GEN_6240 : ~_GEN_373 & _GEN_6240;
  wire        _GEN_6625 = _GEN_385 ? ~_GEN_429 & _GEN_6241 : ~_GEN_374 & _GEN_6241;
  wire        _GEN_6626 = _GEN_385 ? ~_GEN_431 & _GEN_6242 : ~_GEN_375 & _GEN_6242;
  wire        _GEN_6627 = _GEN_385 ? ~_GEN_433 & _GEN_6243 : ~_GEN_376 & _GEN_6243;
  wire        _GEN_6628 = _GEN_385 ? ~_GEN_435 & _GEN_6244 : ~_GEN_377 & _GEN_6244;
  wire        _GEN_6629 = _GEN_385 ? ~_GEN_437 & _GEN_6245 : ~_GEN_378 & _GEN_6245;
  wire        _GEN_6630 = _GEN_385 ? ~_GEN_439 & _GEN_6246 : ~_GEN_379 & _GEN_6246;
  wire        _GEN_6631 = _GEN_385 ? ~_GEN_441 & _GEN_6247 : ~_GEN_380 & _GEN_6247;
  wire        _GEN_6632 = _GEN_385 ? ~_GEN_443 & _GEN_6248 : ~_GEN_381 & _GEN_6248;
  wire        _GEN_6633 = _GEN_385 ? ~_GEN_445 & _GEN_6249 : ~_GEN_382 & _GEN_6249;
  wire        _GEN_6634 = _GEN_385 ? ~_GEN_447 & _GEN_6250 : ~_GEN_383 & _GEN_6250;
  wire        _GEN_6635 = _GEN_385 ? ~_GEN_448 & _GEN_6251 : ~_GEN_384 & _GEN_6251;
  wire        _GEN_6988 = _GEN_513 ? ~_GEN_515 & _GEN_6604 : ~_GEN_481 & _GEN_6604;
  wire        _GEN_6989 = _GEN_513 ? ~_GEN_517 & _GEN_6605 : ~_GEN_482 & _GEN_6605;
  wire        _GEN_6990 = _GEN_513 ? ~_GEN_519 & _GEN_6606 : ~_GEN_483 & _GEN_6606;
  wire        _GEN_6991 = _GEN_513 ? ~_GEN_521 & _GEN_6607 : ~_GEN_484 & _GEN_6607;
  wire        _GEN_6992 = _GEN_513 ? ~_GEN_523 & _GEN_6608 : ~_GEN_485 & _GEN_6608;
  wire        _GEN_6993 = _GEN_513 ? ~_GEN_525 & _GEN_6609 : ~_GEN_486 & _GEN_6609;
  wire        _GEN_6994 = _GEN_513 ? ~_GEN_527 & _GEN_6610 : ~_GEN_487 & _GEN_6610;
  wire        _GEN_6995 = _GEN_513 ? ~_GEN_529 & _GEN_6611 : ~_GEN_488 & _GEN_6611;
  wire        _GEN_6996 = _GEN_513 ? ~_GEN_531 & _GEN_6612 : ~_GEN_489 & _GEN_6612;
  wire        _GEN_6997 = _GEN_513 ? ~_GEN_533 & _GEN_6613 : ~_GEN_490 & _GEN_6613;
  wire        _GEN_6998 = _GEN_513 ? ~_GEN_535 & _GEN_6614 : ~_GEN_491 & _GEN_6614;
  wire        _GEN_6999 = _GEN_513 ? ~_GEN_537 & _GEN_6615 : ~_GEN_492 & _GEN_6615;
  wire        _GEN_7000 = _GEN_513 ? ~_GEN_539 & _GEN_6616 : ~_GEN_493 & _GEN_6616;
  wire        _GEN_7001 = _GEN_513 ? ~_GEN_541 & _GEN_6617 : ~_GEN_494 & _GEN_6617;
  wire        _GEN_7002 = _GEN_513 ? ~_GEN_543 & _GEN_6618 : ~_GEN_495 & _GEN_6618;
  wire        _GEN_7003 = _GEN_513 ? ~_GEN_545 & _GEN_6619 : ~_GEN_496 & _GEN_6619;
  wire        _GEN_7004 = _GEN_513 ? ~_GEN_547 & _GEN_6620 : ~_GEN_497 & _GEN_6620;
  wire        _GEN_7005 = _GEN_513 ? ~_GEN_549 & _GEN_6621 : ~_GEN_498 & _GEN_6621;
  wire        _GEN_7006 = _GEN_513 ? ~_GEN_551 & _GEN_6622 : ~_GEN_499 & _GEN_6622;
  wire        _GEN_7007 = _GEN_513 ? ~_GEN_553 & _GEN_6623 : ~_GEN_500 & _GEN_6623;
  wire        _GEN_7008 = _GEN_513 ? ~_GEN_555 & _GEN_6624 : ~_GEN_501 & _GEN_6624;
  wire        _GEN_7009 = _GEN_513 ? ~_GEN_557 & _GEN_6625 : ~_GEN_502 & _GEN_6625;
  wire        _GEN_7010 = _GEN_513 ? ~_GEN_559 & _GEN_6626 : ~_GEN_503 & _GEN_6626;
  wire        _GEN_7011 = _GEN_513 ? ~_GEN_561 & _GEN_6627 : ~_GEN_504 & _GEN_6627;
  wire        _GEN_7012 = _GEN_513 ? ~_GEN_563 & _GEN_6628 : ~_GEN_505 & _GEN_6628;
  wire        _GEN_7013 = _GEN_513 ? ~_GEN_565 & _GEN_6629 : ~_GEN_506 & _GEN_6629;
  wire        _GEN_7014 = _GEN_513 ? ~_GEN_567 & _GEN_6630 : ~_GEN_507 & _GEN_6630;
  wire        _GEN_7015 = _GEN_513 ? ~_GEN_569 & _GEN_6631 : ~_GEN_508 & _GEN_6631;
  wire        _GEN_7016 = _GEN_513 ? ~_GEN_571 & _GEN_6632 : ~_GEN_509 & _GEN_6632;
  wire        _GEN_7017 = _GEN_513 ? ~_GEN_573 & _GEN_6633 : ~_GEN_510 & _GEN_6633;
  wire        _GEN_7018 = _GEN_513 ? ~_GEN_575 & _GEN_6634 : ~_GEN_511 & _GEN_6634;
  wire        _GEN_7019 = _GEN_513 ? ~_GEN_576 & _GEN_6635 : ~_GEN_512 & _GEN_6635;
  wire        _GEN_7372 = _GEN_641 ? ~_GEN_643 & _GEN_6988 : ~_GEN_609 & _GEN_6988;
  wire        _GEN_7373 = _GEN_641 ? ~_GEN_645 & _GEN_6989 : ~_GEN_610 & _GEN_6989;
  wire        _GEN_7374 = _GEN_641 ? ~_GEN_647 & _GEN_6990 : ~_GEN_611 & _GEN_6990;
  wire        _GEN_7375 = _GEN_641 ? ~_GEN_649 & _GEN_6991 : ~_GEN_612 & _GEN_6991;
  wire        _GEN_7376 = _GEN_641 ? ~_GEN_651 & _GEN_6992 : ~_GEN_613 & _GEN_6992;
  wire        _GEN_7377 = _GEN_641 ? ~_GEN_653 & _GEN_6993 : ~_GEN_614 & _GEN_6993;
  wire        _GEN_7378 = _GEN_641 ? ~_GEN_655 & _GEN_6994 : ~_GEN_615 & _GEN_6994;
  wire        _GEN_7379 = _GEN_641 ? ~_GEN_657 & _GEN_6995 : ~_GEN_616 & _GEN_6995;
  wire        _GEN_7380 = _GEN_641 ? ~_GEN_659 & _GEN_6996 : ~_GEN_617 & _GEN_6996;
  wire        _GEN_7381 = _GEN_641 ? ~_GEN_661 & _GEN_6997 : ~_GEN_618 & _GEN_6997;
  wire        _GEN_7382 = _GEN_641 ? ~_GEN_663 & _GEN_6998 : ~_GEN_619 & _GEN_6998;
  wire        _GEN_7383 = _GEN_641 ? ~_GEN_665 & _GEN_6999 : ~_GEN_620 & _GEN_6999;
  wire        _GEN_7384 = _GEN_641 ? ~_GEN_667 & _GEN_7000 : ~_GEN_621 & _GEN_7000;
  wire        _GEN_7385 = _GEN_641 ? ~_GEN_669 & _GEN_7001 : ~_GEN_622 & _GEN_7001;
  wire        _GEN_7386 = _GEN_641 ? ~_GEN_671 & _GEN_7002 : ~_GEN_623 & _GEN_7002;
  wire        _GEN_7387 = _GEN_641 ? ~_GEN_673 & _GEN_7003 : ~_GEN_624 & _GEN_7003;
  wire        _GEN_7388 = _GEN_641 ? ~_GEN_675 & _GEN_7004 : ~_GEN_625 & _GEN_7004;
  wire        _GEN_7389 = _GEN_641 ? ~_GEN_677 & _GEN_7005 : ~_GEN_626 & _GEN_7005;
  wire        _GEN_7390 = _GEN_641 ? ~_GEN_679 & _GEN_7006 : ~_GEN_627 & _GEN_7006;
  wire        _GEN_7391 = _GEN_641 ? ~_GEN_681 & _GEN_7007 : ~_GEN_628 & _GEN_7007;
  wire        _GEN_7392 = _GEN_641 ? ~_GEN_683 & _GEN_7008 : ~_GEN_629 & _GEN_7008;
  wire        _GEN_7393 = _GEN_641 ? ~_GEN_685 & _GEN_7009 : ~_GEN_630 & _GEN_7009;
  wire        _GEN_7394 = _GEN_641 ? ~_GEN_687 & _GEN_7010 : ~_GEN_631 & _GEN_7010;
  wire        _GEN_7395 = _GEN_641 ? ~_GEN_689 & _GEN_7011 : ~_GEN_632 & _GEN_7011;
  wire        _GEN_7396 = _GEN_641 ? ~_GEN_691 & _GEN_7012 : ~_GEN_633 & _GEN_7012;
  wire        _GEN_7397 = _GEN_641 ? ~_GEN_693 & _GEN_7013 : ~_GEN_634 & _GEN_7013;
  wire        _GEN_7398 = _GEN_641 ? ~_GEN_695 & _GEN_7014 : ~_GEN_635 & _GEN_7014;
  wire        _GEN_7399 = _GEN_641 ? ~_GEN_697 & _GEN_7015 : ~_GEN_636 & _GEN_7015;
  wire        _GEN_7400 = _GEN_641 ? ~_GEN_699 & _GEN_7016 : ~_GEN_637 & _GEN_7016;
  wire        _GEN_7401 = _GEN_641 ? ~_GEN_701 & _GEN_7017 : ~_GEN_638 & _GEN_7017;
  wire        _GEN_7402 = _GEN_641 ? ~_GEN_703 & _GEN_7018 : ~_GEN_639 & _GEN_7018;
  wire        _GEN_7403 = _GEN_641 ? ~_GEN_704 & _GEN_7019 : ~_GEN_640 & _GEN_7019;
  wire        _GEN_2320 = io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_2321 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_2322 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_2323 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_2324 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_2325 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_2326 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_2327 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_2328 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_2329 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_2330 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_2331 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_2332 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_2333 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_2334 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_2335 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_2336 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_2337 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_2338 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_2339 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_2340 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_2341 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_2342 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_2343 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_2344 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_2345 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_2346 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_2347 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_2348 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_2349 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_2350 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_2351 = io_fflags_0_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_2352 = io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_2353 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_2354 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_2355 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_2356 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_2357 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_2358 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_2359 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_2360 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_2361 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_2362 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_2363 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_2364 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_2365 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_2366 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_2367 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_2368 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_2369 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_2370 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_2371 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_2372 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_2373 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_2374 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_2375 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_2376 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_2377 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_2378 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_2379 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_2380 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_2381 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_2382 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_2383 = io_fflags_2_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_2384 = io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h0;
  wire        _GEN_2385 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_2386 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_2387 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_2388 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_2389 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_2390 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_2391 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_2392 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_2393 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_2394 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_2395 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_2396 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_2397 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_2398 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_2399 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_2400 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_2401 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_2402 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_2403 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_2404 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_2405 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_2406 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_2407 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_2408 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_2409 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_2410 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_2411 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_2412 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_2413 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_2414 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_2415 = io_fflags_3_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_2416 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h0;
  wire        _GEN_2417 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1;
  wire        _GEN_2418 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h2;
  wire        _GEN_2419 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h3;
  wire        _GEN_2420 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h4;
  wire        _GEN_2421 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h5;
  wire        _GEN_2422 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h6;
  wire        _GEN_2423 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h7;
  wire        _GEN_2424 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h8;
  wire        _GEN_2425 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h9;
  wire        _GEN_2426 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hA;
  wire        _GEN_2427 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hB;
  wire        _GEN_2428 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hC;
  wire        _GEN_2429 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hD;
  wire        _GEN_2430 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hE;
  wire        _GEN_2431 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'hF;
  wire        _GEN_2432 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h10;
  wire        _GEN_2433 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h11;
  wire        _GEN_2434 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h12;
  wire        _GEN_2435 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h13;
  wire        _GEN_2436 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h14;
  wire        _GEN_2437 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h15;
  wire        _GEN_2438 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h16;
  wire        _GEN_2439 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h17;
  wire        _GEN_2440 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h18;
  wire        _GEN_2441 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h19;
  wire        _GEN_2442 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1A;
  wire        _GEN_2443 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1B;
  wire        _GEN_2444 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1C;
  wire        _GEN_2445 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1D;
  wire        _GEN_2446 = io_lxcpt_bits_uop_rob_idx[6:2] == 5'h1E;
  wire        _GEN_2447 = com_idx == 5'h1;
  wire        _GEN_2448 = com_idx == 5'h2;
  wire        _GEN_2449 = com_idx == 5'h3;
  wire        _GEN_2450 = com_idx == 5'h4;
  wire        _GEN_2451 = com_idx == 5'h5;
  wire        _GEN_2452 = com_idx == 5'h6;
  wire        _GEN_2453 = com_idx == 5'h7;
  wire        _GEN_2454 = com_idx == 5'h8;
  wire        _GEN_2455 = com_idx == 5'h9;
  wire        _GEN_2456 = com_idx == 5'hA;
  wire        _GEN_2457 = com_idx == 5'hB;
  wire        _GEN_2458 = com_idx == 5'hC;
  wire        _GEN_2459 = com_idx == 5'hD;
  wire        _GEN_2460 = com_idx == 5'hE;
  wire        _GEN_2461 = com_idx == 5'hF;
  wire        _GEN_2462 = com_idx == 5'h10;
  wire        _GEN_2463 = com_idx == 5'h11;
  wire        _GEN_2464 = com_idx == 5'h12;
  wire        _GEN_2465 = com_idx == 5'h13;
  wire        _GEN_2466 = com_idx == 5'h14;
  wire        _GEN_2467 = com_idx == 5'h15;
  wire        _GEN_2468 = com_idx == 5'h16;
  wire        _GEN_2469 = com_idx == 5'h17;
  wire        _GEN_2470 = com_idx == 5'h18;
  wire        _GEN_2471 = com_idx == 5'h19;
  wire        _GEN_2472 = com_idx == 5'h1A;
  wire        _GEN_2473 = com_idx == 5'h1B;
  wire        _GEN_2474 = com_idx == 5'h1C;
  wire        _GEN_2475 = com_idx == 5'h1D;
  wire        _GEN_2476 = com_idx == 5'h1E;
  wire        _GEN_2477 = com_idx == 5'h0;
  wire        _GEN_2478 = rbk_row & _GEN_2477;
  wire        _GEN_2479 = rbk_row & _GEN_2447;
  wire        _GEN_2480 = rbk_row & _GEN_2448;
  wire        _GEN_2481 = rbk_row & _GEN_2449;
  wire        _GEN_2482 = rbk_row & _GEN_2450;
  wire        _GEN_2483 = rbk_row & _GEN_2451;
  wire        _GEN_2484 = rbk_row & _GEN_2452;
  wire        _GEN_2485 = rbk_row & _GEN_2453;
  wire        _GEN_2486 = rbk_row & _GEN_2454;
  wire        _GEN_2487 = rbk_row & _GEN_2455;
  wire        _GEN_2488 = rbk_row & _GEN_2456;
  wire        _GEN_2489 = rbk_row & _GEN_2457;
  wire        _GEN_2490 = rbk_row & _GEN_2458;
  wire        _GEN_2491 = rbk_row & _GEN_2459;
  wire        _GEN_2492 = rbk_row & _GEN_2460;
  wire        _GEN_2493 = rbk_row & _GEN_2461;
  wire        _GEN_2494 = rbk_row & _GEN_2462;
  wire        _GEN_2495 = rbk_row & _GEN_2463;
  wire        _GEN_2496 = rbk_row & _GEN_2464;
  wire        _GEN_2497 = rbk_row & _GEN_2465;
  wire        _GEN_2498 = rbk_row & _GEN_2466;
  wire        _GEN_2499 = rbk_row & _GEN_2467;
  wire        _GEN_2500 = rbk_row & _GEN_2468;
  wire        _GEN_2501 = rbk_row & _GEN_2469;
  wire        _GEN_2502 = rbk_row & _GEN_2470;
  wire        _GEN_2503 = rbk_row & _GEN_2471;
  wire        _GEN_2504 = rbk_row & _GEN_2472;
  wire        _GEN_2505 = rbk_row & _GEN_2473;
  wire        _GEN_2506 = rbk_row & _GEN_2474;
  wire        _GEN_2507 = rbk_row & _GEN_2475;
  wire        _GEN_2508 = rbk_row & _GEN_2476;
  wire        _GEN_2509 = rbk_row & (&com_idx);
  wire [19:0] _GEN_2510 = io_brupdate_b1_mispredict_mask & rob_uop__0_br_mask;
  wire [19:0] _GEN_2511 = io_brupdate_b1_mispredict_mask & rob_uop__1_br_mask;
  wire [19:0] _GEN_2512 = io_brupdate_b1_mispredict_mask & rob_uop__2_br_mask;
  wire [19:0] _GEN_2513 = io_brupdate_b1_mispredict_mask & rob_uop__3_br_mask;
  wire [19:0] _GEN_2514 = io_brupdate_b1_mispredict_mask & rob_uop__4_br_mask;
  wire [19:0] _GEN_2515 = io_brupdate_b1_mispredict_mask & rob_uop__5_br_mask;
  wire [19:0] _GEN_2516 = io_brupdate_b1_mispredict_mask & rob_uop__6_br_mask;
  wire [19:0] _GEN_2517 = io_brupdate_b1_mispredict_mask & rob_uop__7_br_mask;
  wire [19:0] _GEN_2518 = io_brupdate_b1_mispredict_mask & rob_uop__8_br_mask;
  wire [19:0] _GEN_2519 = io_brupdate_b1_mispredict_mask & rob_uop__9_br_mask;
  wire [19:0] _GEN_2520 = io_brupdate_b1_mispredict_mask & rob_uop__10_br_mask;
  wire [19:0] _GEN_2521 = io_brupdate_b1_mispredict_mask & rob_uop__11_br_mask;
  wire [19:0] _GEN_2522 = io_brupdate_b1_mispredict_mask & rob_uop__12_br_mask;
  wire [19:0] _GEN_2523 = io_brupdate_b1_mispredict_mask & rob_uop__13_br_mask;
  wire [19:0] _GEN_2524 = io_brupdate_b1_mispredict_mask & rob_uop__14_br_mask;
  wire [19:0] _GEN_2525 = io_brupdate_b1_mispredict_mask & rob_uop__15_br_mask;
  wire [19:0] _GEN_2526 = io_brupdate_b1_mispredict_mask & rob_uop__16_br_mask;
  wire [19:0] _GEN_2527 = io_brupdate_b1_mispredict_mask & rob_uop__17_br_mask;
  wire [19:0] _GEN_2528 = io_brupdate_b1_mispredict_mask & rob_uop__18_br_mask;
  wire [19:0] _GEN_2529 = io_brupdate_b1_mispredict_mask & rob_uop__19_br_mask;
  wire [19:0] _GEN_2530 = io_brupdate_b1_mispredict_mask & rob_uop__20_br_mask;
  wire [19:0] _GEN_2531 = io_brupdate_b1_mispredict_mask & rob_uop__21_br_mask;
  wire [19:0] _GEN_2532 = io_brupdate_b1_mispredict_mask & rob_uop__22_br_mask;
  wire [19:0] _GEN_2533 = io_brupdate_b1_mispredict_mask & rob_uop__23_br_mask;
  wire [19:0] _GEN_2534 = io_brupdate_b1_mispredict_mask & rob_uop__24_br_mask;
  wire [19:0] _GEN_2535 = io_brupdate_b1_mispredict_mask & rob_uop__25_br_mask;
  wire [19:0] _GEN_2536 = io_brupdate_b1_mispredict_mask & rob_uop__26_br_mask;
  wire [19:0] _GEN_2537 = io_brupdate_b1_mispredict_mask & rob_uop__27_br_mask;
  wire [19:0] _GEN_2538 = io_brupdate_b1_mispredict_mask & rob_uop__28_br_mask;
  wire [19:0] _GEN_2539 = io_brupdate_b1_mispredict_mask & rob_uop__29_br_mask;
  wire [19:0] _GEN_2540 = io_brupdate_b1_mispredict_mask & rob_uop__30_br_mask;
  wire [19:0] _GEN_2541 = io_brupdate_b1_mispredict_mask & rob_uop__31_br_mask;
  wire        _rob_bsy_T_2 = io_enq_uops_1_is_fence | io_enq_uops_1_is_fencei;
  wire        _GEN_16224 = _GEN_898 ? ~_rob_bsy_T_2 : rob_bsy_1_0;
  wire        _GEN_16225 = _GEN_899 ? ~_rob_bsy_T_2 : rob_bsy_1_1;
  wire        _GEN_16226 = _GEN_900 ? ~_rob_bsy_T_2 : rob_bsy_1_2;
  wire        _GEN_16227 = _GEN_901 ? ~_rob_bsy_T_2 : rob_bsy_1_3;
  wire        _GEN_16228 = _GEN_902 ? ~_rob_bsy_T_2 : rob_bsy_1_4;
  wire        _GEN_16229 = _GEN_903 ? ~_rob_bsy_T_2 : rob_bsy_1_5;
  wire        _GEN_16230 = _GEN_904 ? ~_rob_bsy_T_2 : rob_bsy_1_6;
  wire        _GEN_16231 = _GEN_905 ? ~_rob_bsy_T_2 : rob_bsy_1_7;
  wire        _GEN_16232 = _GEN_906 ? ~_rob_bsy_T_2 : rob_bsy_1_8;
  wire        _GEN_16233 = _GEN_907 ? ~_rob_bsy_T_2 : rob_bsy_1_9;
  wire        _GEN_16234 = _GEN_908 ? ~_rob_bsy_T_2 : rob_bsy_1_10;
  wire        _GEN_16235 = _GEN_909 ? ~_rob_bsy_T_2 : rob_bsy_1_11;
  wire        _GEN_16236 = _GEN_910 ? ~_rob_bsy_T_2 : rob_bsy_1_12;
  wire        _GEN_16237 = _GEN_911 ? ~_rob_bsy_T_2 : rob_bsy_1_13;
  wire        _GEN_16238 = _GEN_912 ? ~_rob_bsy_T_2 : rob_bsy_1_14;
  wire        _GEN_16239 = _GEN_913 ? ~_rob_bsy_T_2 : rob_bsy_1_15;
  wire        _GEN_16240 = _GEN_914 ? ~_rob_bsy_T_2 : rob_bsy_1_16;
  wire        _GEN_16241 = _GEN_915 ? ~_rob_bsy_T_2 : rob_bsy_1_17;
  wire        _GEN_16242 = _GEN_916 ? ~_rob_bsy_T_2 : rob_bsy_1_18;
  wire        _GEN_16243 = _GEN_917 ? ~_rob_bsy_T_2 : rob_bsy_1_19;
  wire        _GEN_16244 = _GEN_918 ? ~_rob_bsy_T_2 : rob_bsy_1_20;
  wire        _GEN_16245 = _GEN_919 ? ~_rob_bsy_T_2 : rob_bsy_1_21;
  wire        _GEN_16246 = _GEN_920 ? ~_rob_bsy_T_2 : rob_bsy_1_22;
  wire        _GEN_16247 = _GEN_921 ? ~_rob_bsy_T_2 : rob_bsy_1_23;
  wire        _GEN_16248 = _GEN_922 ? ~_rob_bsy_T_2 : rob_bsy_1_24;
  wire        _GEN_16249 = _GEN_923 ? ~_rob_bsy_T_2 : rob_bsy_1_25;
  wire        _GEN_16250 = _GEN_924 ? ~_rob_bsy_T_2 : rob_bsy_1_26;
  wire        _GEN_16251 = _GEN_925 ? ~_rob_bsy_T_2 : rob_bsy_1_27;
  wire        _GEN_16252 = _GEN_926 ? ~_rob_bsy_T_2 : rob_bsy_1_28;
  wire        _GEN_16253 = _GEN_927 ? ~_rob_bsy_T_2 : rob_bsy_1_29;
  wire        _GEN_16254 = _GEN_928 ? ~_rob_bsy_T_2 : rob_bsy_1_30;
  wire        _GEN_16255 = _GEN_929 ? ~_rob_bsy_T_2 : rob_bsy_1_31;
  wire        _GEN_19200 = _GEN_963 ? ~_GEN_964 & _GEN_16224 : ~_GEN_931 & _GEN_16224;
  wire        _GEN_19201 = _GEN_963 ? ~_GEN_965 & _GEN_16225 : ~_GEN_932 & _GEN_16225;
  wire        _GEN_19202 = _GEN_963 ? ~_GEN_966 & _GEN_16226 : ~_GEN_933 & _GEN_16226;
  wire        _GEN_19203 = _GEN_963 ? ~_GEN_967 & _GEN_16227 : ~_GEN_934 & _GEN_16227;
  wire        _GEN_19204 = _GEN_963 ? ~_GEN_968 & _GEN_16228 : ~_GEN_935 & _GEN_16228;
  wire        _GEN_19205 = _GEN_963 ? ~_GEN_969 & _GEN_16229 : ~_GEN_936 & _GEN_16229;
  wire        _GEN_19206 = _GEN_963 ? ~_GEN_970 & _GEN_16230 : ~_GEN_937 & _GEN_16230;
  wire        _GEN_19207 = _GEN_963 ? ~_GEN_971 & _GEN_16231 : ~_GEN_938 & _GEN_16231;
  wire        _GEN_19208 = _GEN_963 ? ~_GEN_972 & _GEN_16232 : ~_GEN_939 & _GEN_16232;
  wire        _GEN_19209 = _GEN_963 ? ~_GEN_973 & _GEN_16233 : ~_GEN_940 & _GEN_16233;
  wire        _GEN_19210 = _GEN_963 ? ~_GEN_974 & _GEN_16234 : ~_GEN_941 & _GEN_16234;
  wire        _GEN_19211 = _GEN_963 ? ~_GEN_975 & _GEN_16235 : ~_GEN_942 & _GEN_16235;
  wire        _GEN_19212 = _GEN_963 ? ~_GEN_976 & _GEN_16236 : ~_GEN_943 & _GEN_16236;
  wire        _GEN_19213 = _GEN_963 ? ~_GEN_977 & _GEN_16237 : ~_GEN_944 & _GEN_16237;
  wire        _GEN_19214 = _GEN_963 ? ~_GEN_978 & _GEN_16238 : ~_GEN_945 & _GEN_16238;
  wire        _GEN_19215 = _GEN_963 ? ~_GEN_979 & _GEN_16239 : ~_GEN_946 & _GEN_16239;
  wire        _GEN_19216 = _GEN_963 ? ~_GEN_980 & _GEN_16240 : ~_GEN_947 & _GEN_16240;
  wire        _GEN_19217 = _GEN_963 ? ~_GEN_981 & _GEN_16241 : ~_GEN_948 & _GEN_16241;
  wire        _GEN_19218 = _GEN_963 ? ~_GEN_982 & _GEN_16242 : ~_GEN_949 & _GEN_16242;
  wire        _GEN_19219 = _GEN_963 ? ~_GEN_983 & _GEN_16243 : ~_GEN_950 & _GEN_16243;
  wire        _GEN_19220 = _GEN_963 ? ~_GEN_984 & _GEN_16244 : ~_GEN_951 & _GEN_16244;
  wire        _GEN_19221 = _GEN_963 ? ~_GEN_985 & _GEN_16245 : ~_GEN_952 & _GEN_16245;
  wire        _GEN_19222 = _GEN_963 ? ~_GEN_986 & _GEN_16246 : ~_GEN_953 & _GEN_16246;
  wire        _GEN_19223 = _GEN_963 ? ~_GEN_987 & _GEN_16247 : ~_GEN_954 & _GEN_16247;
  wire        _GEN_19224 = _GEN_963 ? ~_GEN_988 & _GEN_16248 : ~_GEN_955 & _GEN_16248;
  wire        _GEN_19225 = _GEN_963 ? ~_GEN_989 & _GEN_16249 : ~_GEN_956 & _GEN_16249;
  wire        _GEN_19226 = _GEN_963 ? ~_GEN_990 & _GEN_16250 : ~_GEN_957 & _GEN_16250;
  wire        _GEN_19227 = _GEN_963 ? ~_GEN_991 & _GEN_16251 : ~_GEN_958 & _GEN_16251;
  wire        _GEN_19228 = _GEN_963 ? ~_GEN_992 & _GEN_16252 : ~_GEN_959 & _GEN_16252;
  wire        _GEN_19229 = _GEN_963 ? ~_GEN_993 & _GEN_16253 : ~_GEN_960 & _GEN_16253;
  wire        _GEN_19230 = _GEN_963 ? ~_GEN_994 & _GEN_16254 : ~_GEN_961 & _GEN_16254;
  wire        _GEN_19231 = _GEN_963 ? ~_GEN_995 & _GEN_16255 : ~_GEN_962 & _GEN_16255;
  wire        _GEN_19584 = _GEN_1029 ? ~_GEN_1030 & _GEN_19200 : ~_GEN_997 & _GEN_19200;
  wire        _GEN_19585 = _GEN_1029 ? ~_GEN_1031 & _GEN_19201 : ~_GEN_998 & _GEN_19201;
  wire        _GEN_19586 = _GEN_1029 ? ~_GEN_1032 & _GEN_19202 : ~_GEN_999 & _GEN_19202;
  wire        _GEN_19587 = _GEN_1029 ? ~_GEN_1033 & _GEN_19203 : ~_GEN_1000 & _GEN_19203;
  wire        _GEN_19588 = _GEN_1029 ? ~_GEN_1034 & _GEN_19204 : ~_GEN_1001 & _GEN_19204;
  wire        _GEN_19589 = _GEN_1029 ? ~_GEN_1035 & _GEN_19205 : ~_GEN_1002 & _GEN_19205;
  wire        _GEN_19590 = _GEN_1029 ? ~_GEN_1036 & _GEN_19206 : ~_GEN_1003 & _GEN_19206;
  wire        _GEN_19591 = _GEN_1029 ? ~_GEN_1037 & _GEN_19207 : ~_GEN_1004 & _GEN_19207;
  wire        _GEN_19592 = _GEN_1029 ? ~_GEN_1038 & _GEN_19208 : ~_GEN_1005 & _GEN_19208;
  wire        _GEN_19593 = _GEN_1029 ? ~_GEN_1039 & _GEN_19209 : ~_GEN_1006 & _GEN_19209;
  wire        _GEN_19594 = _GEN_1029 ? ~_GEN_1040 & _GEN_19210 : ~_GEN_1007 & _GEN_19210;
  wire        _GEN_19595 = _GEN_1029 ? ~_GEN_1041 & _GEN_19211 : ~_GEN_1008 & _GEN_19211;
  wire        _GEN_19596 = _GEN_1029 ? ~_GEN_1042 & _GEN_19212 : ~_GEN_1009 & _GEN_19212;
  wire        _GEN_19597 = _GEN_1029 ? ~_GEN_1043 & _GEN_19213 : ~_GEN_1010 & _GEN_19213;
  wire        _GEN_19598 = _GEN_1029 ? ~_GEN_1044 & _GEN_19214 : ~_GEN_1011 & _GEN_19214;
  wire        _GEN_19599 = _GEN_1029 ? ~_GEN_1045 & _GEN_19215 : ~_GEN_1012 & _GEN_19215;
  wire        _GEN_19600 = _GEN_1029 ? ~_GEN_1046 & _GEN_19216 : ~_GEN_1013 & _GEN_19216;
  wire        _GEN_19601 = _GEN_1029 ? ~_GEN_1047 & _GEN_19217 : ~_GEN_1014 & _GEN_19217;
  wire        _GEN_19602 = _GEN_1029 ? ~_GEN_1048 & _GEN_19218 : ~_GEN_1015 & _GEN_19218;
  wire        _GEN_19603 = _GEN_1029 ? ~_GEN_1049 & _GEN_19219 : ~_GEN_1016 & _GEN_19219;
  wire        _GEN_19604 = _GEN_1029 ? ~_GEN_1050 & _GEN_19220 : ~_GEN_1017 & _GEN_19220;
  wire        _GEN_19605 = _GEN_1029 ? ~_GEN_1051 & _GEN_19221 : ~_GEN_1018 & _GEN_19221;
  wire        _GEN_19606 = _GEN_1029 ? ~_GEN_1052 & _GEN_19222 : ~_GEN_1019 & _GEN_19222;
  wire        _GEN_19607 = _GEN_1029 ? ~_GEN_1053 & _GEN_19223 : ~_GEN_1020 & _GEN_19223;
  wire        _GEN_19608 = _GEN_1029 ? ~_GEN_1054 & _GEN_19224 : ~_GEN_1021 & _GEN_19224;
  wire        _GEN_19609 = _GEN_1029 ? ~_GEN_1055 & _GEN_19225 : ~_GEN_1022 & _GEN_19225;
  wire        _GEN_19610 = _GEN_1029 ? ~_GEN_1056 & _GEN_19226 : ~_GEN_1023 & _GEN_19226;
  wire        _GEN_19611 = _GEN_1029 ? ~_GEN_1057 & _GEN_19227 : ~_GEN_1024 & _GEN_19227;
  wire        _GEN_19612 = _GEN_1029 ? ~_GEN_1058 & _GEN_19228 : ~_GEN_1025 & _GEN_19228;
  wire        _GEN_19613 = _GEN_1029 ? ~_GEN_1059 & _GEN_19229 : ~_GEN_1026 & _GEN_19229;
  wire        _GEN_19614 = _GEN_1029 ? ~_GEN_1060 & _GEN_19230 : ~_GEN_1027 & _GEN_19230;
  wire        _GEN_19615 = _GEN_1029 ? ~_GEN_1061 & _GEN_19231 : ~_GEN_1028 & _GEN_19231;
  wire        _GEN_19968 = _GEN_1095 ? ~_GEN_1096 & _GEN_19584 : ~_GEN_1063 & _GEN_19584;
  wire        _GEN_19969 = _GEN_1095 ? ~_GEN_1097 & _GEN_19585 : ~_GEN_1064 & _GEN_19585;
  wire        _GEN_19970 = _GEN_1095 ? ~_GEN_1098 & _GEN_19586 : ~_GEN_1065 & _GEN_19586;
  wire        _GEN_19971 = _GEN_1095 ? ~_GEN_1099 & _GEN_19587 : ~_GEN_1066 & _GEN_19587;
  wire        _GEN_19972 = _GEN_1095 ? ~_GEN_1100 & _GEN_19588 : ~_GEN_1067 & _GEN_19588;
  wire        _GEN_19973 = _GEN_1095 ? ~_GEN_1101 & _GEN_19589 : ~_GEN_1068 & _GEN_19589;
  wire        _GEN_19974 = _GEN_1095 ? ~_GEN_1102 & _GEN_19590 : ~_GEN_1069 & _GEN_19590;
  wire        _GEN_19975 = _GEN_1095 ? ~_GEN_1103 & _GEN_19591 : ~_GEN_1070 & _GEN_19591;
  wire        _GEN_19976 = _GEN_1095 ? ~_GEN_1104 & _GEN_19592 : ~_GEN_1071 & _GEN_19592;
  wire        _GEN_19977 = _GEN_1095 ? ~_GEN_1105 & _GEN_19593 : ~_GEN_1072 & _GEN_19593;
  wire        _GEN_19978 = _GEN_1095 ? ~_GEN_1106 & _GEN_19594 : ~_GEN_1073 & _GEN_19594;
  wire        _GEN_19979 = _GEN_1095 ? ~_GEN_1107 & _GEN_19595 : ~_GEN_1074 & _GEN_19595;
  wire        _GEN_19980 = _GEN_1095 ? ~_GEN_1108 & _GEN_19596 : ~_GEN_1075 & _GEN_19596;
  wire        _GEN_19981 = _GEN_1095 ? ~_GEN_1109 & _GEN_19597 : ~_GEN_1076 & _GEN_19597;
  wire        _GEN_19982 = _GEN_1095 ? ~_GEN_1110 & _GEN_19598 : ~_GEN_1077 & _GEN_19598;
  wire        _GEN_19983 = _GEN_1095 ? ~_GEN_1111 & _GEN_19599 : ~_GEN_1078 & _GEN_19599;
  wire        _GEN_19984 = _GEN_1095 ? ~_GEN_1112 & _GEN_19600 : ~_GEN_1079 & _GEN_19600;
  wire        _GEN_19985 = _GEN_1095 ? ~_GEN_1113 & _GEN_19601 : ~_GEN_1080 & _GEN_19601;
  wire        _GEN_19986 = _GEN_1095 ? ~_GEN_1114 & _GEN_19602 : ~_GEN_1081 & _GEN_19602;
  wire        _GEN_19987 = _GEN_1095 ? ~_GEN_1115 & _GEN_19603 : ~_GEN_1082 & _GEN_19603;
  wire        _GEN_19988 = _GEN_1095 ? ~_GEN_1116 & _GEN_19604 : ~_GEN_1083 & _GEN_19604;
  wire        _GEN_19989 = _GEN_1095 ? ~_GEN_1117 & _GEN_19605 : ~_GEN_1084 & _GEN_19605;
  wire        _GEN_19990 = _GEN_1095 ? ~_GEN_1118 & _GEN_19606 : ~_GEN_1085 & _GEN_19606;
  wire        _GEN_19991 = _GEN_1095 ? ~_GEN_1119 & _GEN_19607 : ~_GEN_1086 & _GEN_19607;
  wire        _GEN_19992 = _GEN_1095 ? ~_GEN_1120 & _GEN_19608 : ~_GEN_1087 & _GEN_19608;
  wire        _GEN_19993 = _GEN_1095 ? ~_GEN_1121 & _GEN_19609 : ~_GEN_1088 & _GEN_19609;
  wire        _GEN_19994 = _GEN_1095 ? ~_GEN_1122 & _GEN_19610 : ~_GEN_1089 & _GEN_19610;
  wire        _GEN_19995 = _GEN_1095 ? ~_GEN_1123 & _GEN_19611 : ~_GEN_1090 & _GEN_19611;
  wire        _GEN_19996 = _GEN_1095 ? ~_GEN_1124 & _GEN_19612 : ~_GEN_1091 & _GEN_19612;
  wire        _GEN_19997 = _GEN_1095 ? ~_GEN_1125 & _GEN_19613 : ~_GEN_1092 & _GEN_19613;
  wire        _GEN_19998 = _GEN_1095 ? ~_GEN_1126 & _GEN_19614 : ~_GEN_1093 & _GEN_19614;
  wire        _GEN_19999 = _GEN_1095 ? ~_GEN_1127 & _GEN_19615 : ~_GEN_1094 & _GEN_19615;
  wire        _GEN_20352 = _GEN_1161 ? ~_GEN_1162 & _GEN_19968 : ~_GEN_1129 & _GEN_19968;
  wire        _GEN_20353 = _GEN_1161 ? ~_GEN_1163 & _GEN_19969 : ~_GEN_1130 & _GEN_19969;
  wire        _GEN_20354 = _GEN_1161 ? ~_GEN_1164 & _GEN_19970 : ~_GEN_1131 & _GEN_19970;
  wire        _GEN_20355 = _GEN_1161 ? ~_GEN_1165 & _GEN_19971 : ~_GEN_1132 & _GEN_19971;
  wire        _GEN_20356 = _GEN_1161 ? ~_GEN_1166 & _GEN_19972 : ~_GEN_1133 & _GEN_19972;
  wire        _GEN_20357 = _GEN_1161 ? ~_GEN_1167 & _GEN_19973 : ~_GEN_1134 & _GEN_19973;
  wire        _GEN_20358 = _GEN_1161 ? ~_GEN_1168 & _GEN_19974 : ~_GEN_1135 & _GEN_19974;
  wire        _GEN_20359 = _GEN_1161 ? ~_GEN_1169 & _GEN_19975 : ~_GEN_1136 & _GEN_19975;
  wire        _GEN_20360 = _GEN_1161 ? ~_GEN_1170 & _GEN_19976 : ~_GEN_1137 & _GEN_19976;
  wire        _GEN_20361 = _GEN_1161 ? ~_GEN_1171 & _GEN_19977 : ~_GEN_1138 & _GEN_19977;
  wire        _GEN_20362 = _GEN_1161 ? ~_GEN_1172 & _GEN_19978 : ~_GEN_1139 & _GEN_19978;
  wire        _GEN_20363 = _GEN_1161 ? ~_GEN_1173 & _GEN_19979 : ~_GEN_1140 & _GEN_19979;
  wire        _GEN_20364 = _GEN_1161 ? ~_GEN_1174 & _GEN_19980 : ~_GEN_1141 & _GEN_19980;
  wire        _GEN_20365 = _GEN_1161 ? ~_GEN_1175 & _GEN_19981 : ~_GEN_1142 & _GEN_19981;
  wire        _GEN_20366 = _GEN_1161 ? ~_GEN_1176 & _GEN_19982 : ~_GEN_1143 & _GEN_19982;
  wire        _GEN_20367 = _GEN_1161 ? ~_GEN_1177 & _GEN_19983 : ~_GEN_1144 & _GEN_19983;
  wire        _GEN_20368 = _GEN_1161 ? ~_GEN_1178 & _GEN_19984 : ~_GEN_1145 & _GEN_19984;
  wire        _GEN_20369 = _GEN_1161 ? ~_GEN_1179 & _GEN_19985 : ~_GEN_1146 & _GEN_19985;
  wire        _GEN_20370 = _GEN_1161 ? ~_GEN_1180 & _GEN_19986 : ~_GEN_1147 & _GEN_19986;
  wire        _GEN_20371 = _GEN_1161 ? ~_GEN_1181 & _GEN_19987 : ~_GEN_1148 & _GEN_19987;
  wire        _GEN_20372 = _GEN_1161 ? ~_GEN_1182 & _GEN_19988 : ~_GEN_1149 & _GEN_19988;
  wire        _GEN_20373 = _GEN_1161 ? ~_GEN_1183 & _GEN_19989 : ~_GEN_1150 & _GEN_19989;
  wire        _GEN_20374 = _GEN_1161 ? ~_GEN_1184 & _GEN_19990 : ~_GEN_1151 & _GEN_19990;
  wire        _GEN_20375 = _GEN_1161 ? ~_GEN_1185 & _GEN_19991 : ~_GEN_1152 & _GEN_19991;
  wire        _GEN_20376 = _GEN_1161 ? ~_GEN_1186 & _GEN_19992 : ~_GEN_1153 & _GEN_19992;
  wire        _GEN_20377 = _GEN_1161 ? ~_GEN_1187 & _GEN_19993 : ~_GEN_1154 & _GEN_19993;
  wire        _GEN_20378 = _GEN_1161 ? ~_GEN_1188 & _GEN_19994 : ~_GEN_1155 & _GEN_19994;
  wire        _GEN_20379 = _GEN_1161 ? ~_GEN_1189 & _GEN_19995 : ~_GEN_1156 & _GEN_19995;
  wire        _GEN_20380 = _GEN_1161 ? ~_GEN_1190 & _GEN_19996 : ~_GEN_1157 & _GEN_19996;
  wire        _GEN_20381 = _GEN_1161 ? ~_GEN_1191 & _GEN_19997 : ~_GEN_1158 & _GEN_19997;
  wire        _GEN_20382 = _GEN_1161 ? ~_GEN_1192 & _GEN_19998 : ~_GEN_1159 & _GEN_19998;
  wire        _GEN_20383 = _GEN_1161 ? ~_GEN_1193 & _GEN_19999 : ~_GEN_1160 & _GEN_19999;
  wire        _GEN_20736 = _GEN_1227 ? ~_GEN_1228 & _GEN_20352 : ~_GEN_1195 & _GEN_20352;
  wire        _GEN_20737 = _GEN_1227 ? ~_GEN_1229 & _GEN_20353 : ~_GEN_1196 & _GEN_20353;
  wire        _GEN_20738 = _GEN_1227 ? ~_GEN_1230 & _GEN_20354 : ~_GEN_1197 & _GEN_20354;
  wire        _GEN_20739 = _GEN_1227 ? ~_GEN_1231 & _GEN_20355 : ~_GEN_1198 & _GEN_20355;
  wire        _GEN_20740 = _GEN_1227 ? ~_GEN_1232 & _GEN_20356 : ~_GEN_1199 & _GEN_20356;
  wire        _GEN_20741 = _GEN_1227 ? ~_GEN_1233 & _GEN_20357 : ~_GEN_1200 & _GEN_20357;
  wire        _GEN_20742 = _GEN_1227 ? ~_GEN_1234 & _GEN_20358 : ~_GEN_1201 & _GEN_20358;
  wire        _GEN_20743 = _GEN_1227 ? ~_GEN_1235 & _GEN_20359 : ~_GEN_1202 & _GEN_20359;
  wire        _GEN_20744 = _GEN_1227 ? ~_GEN_1236 & _GEN_20360 : ~_GEN_1203 & _GEN_20360;
  wire        _GEN_20745 = _GEN_1227 ? ~_GEN_1237 & _GEN_20361 : ~_GEN_1204 & _GEN_20361;
  wire        _GEN_20746 = _GEN_1227 ? ~_GEN_1238 & _GEN_20362 : ~_GEN_1205 & _GEN_20362;
  wire        _GEN_20747 = _GEN_1227 ? ~_GEN_1239 & _GEN_20363 : ~_GEN_1206 & _GEN_20363;
  wire        _GEN_20748 = _GEN_1227 ? ~_GEN_1240 & _GEN_20364 : ~_GEN_1207 & _GEN_20364;
  wire        _GEN_20749 = _GEN_1227 ? ~_GEN_1241 & _GEN_20365 : ~_GEN_1208 & _GEN_20365;
  wire        _GEN_20750 = _GEN_1227 ? ~_GEN_1242 & _GEN_20366 : ~_GEN_1209 & _GEN_20366;
  wire        _GEN_20751 = _GEN_1227 ? ~_GEN_1243 & _GEN_20367 : ~_GEN_1210 & _GEN_20367;
  wire        _GEN_20752 = _GEN_1227 ? ~_GEN_1244 & _GEN_20368 : ~_GEN_1211 & _GEN_20368;
  wire        _GEN_20753 = _GEN_1227 ? ~_GEN_1245 & _GEN_20369 : ~_GEN_1212 & _GEN_20369;
  wire        _GEN_20754 = _GEN_1227 ? ~_GEN_1246 & _GEN_20370 : ~_GEN_1213 & _GEN_20370;
  wire        _GEN_20755 = _GEN_1227 ? ~_GEN_1247 & _GEN_20371 : ~_GEN_1214 & _GEN_20371;
  wire        _GEN_20756 = _GEN_1227 ? ~_GEN_1248 & _GEN_20372 : ~_GEN_1215 & _GEN_20372;
  wire        _GEN_20757 = _GEN_1227 ? ~_GEN_1249 & _GEN_20373 : ~_GEN_1216 & _GEN_20373;
  wire        _GEN_20758 = _GEN_1227 ? ~_GEN_1250 & _GEN_20374 : ~_GEN_1217 & _GEN_20374;
  wire        _GEN_20759 = _GEN_1227 ? ~_GEN_1251 & _GEN_20375 : ~_GEN_1218 & _GEN_20375;
  wire        _GEN_20760 = _GEN_1227 ? ~_GEN_1252 & _GEN_20376 : ~_GEN_1219 & _GEN_20376;
  wire        _GEN_20761 = _GEN_1227 ? ~_GEN_1253 & _GEN_20377 : ~_GEN_1220 & _GEN_20377;
  wire        _GEN_20762 = _GEN_1227 ? ~_GEN_1254 & _GEN_20378 : ~_GEN_1221 & _GEN_20378;
  wire        _GEN_20763 = _GEN_1227 ? ~_GEN_1255 & _GEN_20379 : ~_GEN_1222 & _GEN_20379;
  wire        _GEN_20764 = _GEN_1227 ? ~_GEN_1256 & _GEN_20380 : ~_GEN_1223 & _GEN_20380;
  wire        _GEN_20765 = _GEN_1227 ? ~_GEN_1257 & _GEN_20381 : ~_GEN_1224 & _GEN_20381;
  wire        _GEN_20766 = _GEN_1227 ? ~_GEN_1258 & _GEN_20382 : ~_GEN_1225 & _GEN_20382;
  wire        _GEN_20767 = _GEN_1227 ? ~_GEN_1259 & _GEN_20383 : ~_GEN_1226 & _GEN_20383;
  wire        _GEN_2542 = io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_2543 = io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_2544 = io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h1;
  wire        _GEN_2545 = rbk_row_1 & _GEN_2477;
  wire        _GEN_2546 = rbk_row_1 & _GEN_2447;
  wire        _GEN_2547 = rbk_row_1 & _GEN_2448;
  wire        _GEN_2548 = rbk_row_1 & _GEN_2449;
  wire        _GEN_2549 = rbk_row_1 & _GEN_2450;
  wire        _GEN_2550 = rbk_row_1 & _GEN_2451;
  wire        _GEN_2551 = rbk_row_1 & _GEN_2452;
  wire        _GEN_2552 = rbk_row_1 & _GEN_2453;
  wire        _GEN_2553 = rbk_row_1 & _GEN_2454;
  wire        _GEN_2554 = rbk_row_1 & _GEN_2455;
  wire        _GEN_2555 = rbk_row_1 & _GEN_2456;
  wire        _GEN_2556 = rbk_row_1 & _GEN_2457;
  wire        _GEN_2557 = rbk_row_1 & _GEN_2458;
  wire        _GEN_2558 = rbk_row_1 & _GEN_2459;
  wire        _GEN_2559 = rbk_row_1 & _GEN_2460;
  wire        _GEN_2560 = rbk_row_1 & _GEN_2461;
  wire        _GEN_2561 = rbk_row_1 & _GEN_2462;
  wire        _GEN_2562 = rbk_row_1 & _GEN_2463;
  wire        _GEN_2563 = rbk_row_1 & _GEN_2464;
  wire        _GEN_2564 = rbk_row_1 & _GEN_2465;
  wire        _GEN_2565 = rbk_row_1 & _GEN_2466;
  wire        _GEN_2566 = rbk_row_1 & _GEN_2467;
  wire        _GEN_2567 = rbk_row_1 & _GEN_2468;
  wire        _GEN_2568 = rbk_row_1 & _GEN_2469;
  wire        _GEN_2569 = rbk_row_1 & _GEN_2470;
  wire        _GEN_2570 = rbk_row_1 & _GEN_2471;
  wire        _GEN_2571 = rbk_row_1 & _GEN_2472;
  wire        _GEN_2572 = rbk_row_1 & _GEN_2473;
  wire        _GEN_2573 = rbk_row_1 & _GEN_2474;
  wire        _GEN_2574 = rbk_row_1 & _GEN_2475;
  wire        _GEN_2575 = rbk_row_1 & _GEN_2476;
  wire        _GEN_2576 = rbk_row_1 & (&com_idx);
  wire [19:0] _GEN_2577 = io_brupdate_b1_mispredict_mask & rob_uop_1_0_br_mask;
  wire [19:0] _GEN_2578 = io_brupdate_b1_mispredict_mask & rob_uop_1_1_br_mask;
  wire [19:0] _GEN_2579 = io_brupdate_b1_mispredict_mask & rob_uop_1_2_br_mask;
  wire [19:0] _GEN_2580 = io_brupdate_b1_mispredict_mask & rob_uop_1_3_br_mask;
  wire [19:0] _GEN_2581 = io_brupdate_b1_mispredict_mask & rob_uop_1_4_br_mask;
  wire [19:0] _GEN_2582 = io_brupdate_b1_mispredict_mask & rob_uop_1_5_br_mask;
  wire [19:0] _GEN_2583 = io_brupdate_b1_mispredict_mask & rob_uop_1_6_br_mask;
  wire [19:0] _GEN_2584 = io_brupdate_b1_mispredict_mask & rob_uop_1_7_br_mask;
  wire [19:0] _GEN_2585 = io_brupdate_b1_mispredict_mask & rob_uop_1_8_br_mask;
  wire [19:0] _GEN_2586 = io_brupdate_b1_mispredict_mask & rob_uop_1_9_br_mask;
  wire [19:0] _GEN_2587 = io_brupdate_b1_mispredict_mask & rob_uop_1_10_br_mask;
  wire [19:0] _GEN_2588 = io_brupdate_b1_mispredict_mask & rob_uop_1_11_br_mask;
  wire [19:0] _GEN_2589 = io_brupdate_b1_mispredict_mask & rob_uop_1_12_br_mask;
  wire [19:0] _GEN_2590 = io_brupdate_b1_mispredict_mask & rob_uop_1_13_br_mask;
  wire [19:0] _GEN_2591 = io_brupdate_b1_mispredict_mask & rob_uop_1_14_br_mask;
  wire [19:0] _GEN_2592 = io_brupdate_b1_mispredict_mask & rob_uop_1_15_br_mask;
  wire [19:0] _GEN_2593 = io_brupdate_b1_mispredict_mask & rob_uop_1_16_br_mask;
  wire [19:0] _GEN_2594 = io_brupdate_b1_mispredict_mask & rob_uop_1_17_br_mask;
  wire [19:0] _GEN_2595 = io_brupdate_b1_mispredict_mask & rob_uop_1_18_br_mask;
  wire [19:0] _GEN_2596 = io_brupdate_b1_mispredict_mask & rob_uop_1_19_br_mask;
  wire [19:0] _GEN_2597 = io_brupdate_b1_mispredict_mask & rob_uop_1_20_br_mask;
  wire [19:0] _GEN_2598 = io_brupdate_b1_mispredict_mask & rob_uop_1_21_br_mask;
  wire [19:0] _GEN_2599 = io_brupdate_b1_mispredict_mask & rob_uop_1_22_br_mask;
  wire [19:0] _GEN_2600 = io_brupdate_b1_mispredict_mask & rob_uop_1_23_br_mask;
  wire [19:0] _GEN_2601 = io_brupdate_b1_mispredict_mask & rob_uop_1_24_br_mask;
  wire [19:0] _GEN_2602 = io_brupdate_b1_mispredict_mask & rob_uop_1_25_br_mask;
  wire [19:0] _GEN_2603 = io_brupdate_b1_mispredict_mask & rob_uop_1_26_br_mask;
  wire [19:0] _GEN_2604 = io_brupdate_b1_mispredict_mask & rob_uop_1_27_br_mask;
  wire [19:0] _GEN_2605 = io_brupdate_b1_mispredict_mask & rob_uop_1_28_br_mask;
  wire [19:0] _GEN_2606 = io_brupdate_b1_mispredict_mask & rob_uop_1_29_br_mask;
  wire [19:0] _GEN_2607 = io_brupdate_b1_mispredict_mask & rob_uop_1_30_br_mask;
  wire [19:0] _GEN_2608 = io_brupdate_b1_mispredict_mask & rob_uop_1_31_br_mask;
  wire        _rob_bsy_T_4 = io_enq_uops_2_is_fence | io_enq_uops_2_is_fencei;
  wire        _GEN_29588 = _GEN_1360 ? ~_rob_bsy_T_4 : rob_bsy_2_0;
  wire        _GEN_29589 = _GEN_1361 ? ~_rob_bsy_T_4 : rob_bsy_2_1;
  wire        _GEN_29590 = _GEN_1362 ? ~_rob_bsy_T_4 : rob_bsy_2_2;
  wire        _GEN_29591 = _GEN_1363 ? ~_rob_bsy_T_4 : rob_bsy_2_3;
  wire        _GEN_29592 = _GEN_1364 ? ~_rob_bsy_T_4 : rob_bsy_2_4;
  wire        _GEN_29593 = _GEN_1365 ? ~_rob_bsy_T_4 : rob_bsy_2_5;
  wire        _GEN_29594 = _GEN_1366 ? ~_rob_bsy_T_4 : rob_bsy_2_6;
  wire        _GEN_29595 = _GEN_1367 ? ~_rob_bsy_T_4 : rob_bsy_2_7;
  wire        _GEN_29596 = _GEN_1368 ? ~_rob_bsy_T_4 : rob_bsy_2_8;
  wire        _GEN_29597 = _GEN_1369 ? ~_rob_bsy_T_4 : rob_bsy_2_9;
  wire        _GEN_29598 = _GEN_1370 ? ~_rob_bsy_T_4 : rob_bsy_2_10;
  wire        _GEN_29599 = _GEN_1371 ? ~_rob_bsy_T_4 : rob_bsy_2_11;
  wire        _GEN_29600 = _GEN_1372 ? ~_rob_bsy_T_4 : rob_bsy_2_12;
  wire        _GEN_29601 = _GEN_1373 ? ~_rob_bsy_T_4 : rob_bsy_2_13;
  wire        _GEN_29602 = _GEN_1374 ? ~_rob_bsy_T_4 : rob_bsy_2_14;
  wire        _GEN_29603 = _GEN_1375 ? ~_rob_bsy_T_4 : rob_bsy_2_15;
  wire        _GEN_29604 = _GEN_1376 ? ~_rob_bsy_T_4 : rob_bsy_2_16;
  wire        _GEN_29605 = _GEN_1377 ? ~_rob_bsy_T_4 : rob_bsy_2_17;
  wire        _GEN_29606 = _GEN_1378 ? ~_rob_bsy_T_4 : rob_bsy_2_18;
  wire        _GEN_29607 = _GEN_1379 ? ~_rob_bsy_T_4 : rob_bsy_2_19;
  wire        _GEN_29608 = _GEN_1380 ? ~_rob_bsy_T_4 : rob_bsy_2_20;
  wire        _GEN_29609 = _GEN_1381 ? ~_rob_bsy_T_4 : rob_bsy_2_21;
  wire        _GEN_29610 = _GEN_1382 ? ~_rob_bsy_T_4 : rob_bsy_2_22;
  wire        _GEN_29611 = _GEN_1383 ? ~_rob_bsy_T_4 : rob_bsy_2_23;
  wire        _GEN_29612 = _GEN_1384 ? ~_rob_bsy_T_4 : rob_bsy_2_24;
  wire        _GEN_29613 = _GEN_1385 ? ~_rob_bsy_T_4 : rob_bsy_2_25;
  wire        _GEN_29614 = _GEN_1386 ? ~_rob_bsy_T_4 : rob_bsy_2_26;
  wire        _GEN_29615 = _GEN_1387 ? ~_rob_bsy_T_4 : rob_bsy_2_27;
  wire        _GEN_29616 = _GEN_1388 ? ~_rob_bsy_T_4 : rob_bsy_2_28;
  wire        _GEN_29617 = _GEN_1389 ? ~_rob_bsy_T_4 : rob_bsy_2_29;
  wire        _GEN_29618 = _GEN_1390 ? ~_rob_bsy_T_4 : rob_bsy_2_30;
  wire        _GEN_29619 = _GEN_1391 ? ~_rob_bsy_T_4 : rob_bsy_2_31;
  wire        _GEN_32564 = _GEN_1425 ? ~_GEN_1426 & _GEN_29588 : ~_GEN_1393 & _GEN_29588;
  wire        _GEN_32565 = _GEN_1425 ? ~_GEN_1427 & _GEN_29589 : ~_GEN_1394 & _GEN_29589;
  wire        _GEN_32566 = _GEN_1425 ? ~_GEN_1428 & _GEN_29590 : ~_GEN_1395 & _GEN_29590;
  wire        _GEN_32567 = _GEN_1425 ? ~_GEN_1429 & _GEN_29591 : ~_GEN_1396 & _GEN_29591;
  wire        _GEN_32568 = _GEN_1425 ? ~_GEN_1430 & _GEN_29592 : ~_GEN_1397 & _GEN_29592;
  wire        _GEN_32569 = _GEN_1425 ? ~_GEN_1431 & _GEN_29593 : ~_GEN_1398 & _GEN_29593;
  wire        _GEN_32570 = _GEN_1425 ? ~_GEN_1432 & _GEN_29594 : ~_GEN_1399 & _GEN_29594;
  wire        _GEN_32571 = _GEN_1425 ? ~_GEN_1433 & _GEN_29595 : ~_GEN_1400 & _GEN_29595;
  wire        _GEN_32572 = _GEN_1425 ? ~_GEN_1434 & _GEN_29596 : ~_GEN_1401 & _GEN_29596;
  wire        _GEN_32573 = _GEN_1425 ? ~_GEN_1435 & _GEN_29597 : ~_GEN_1402 & _GEN_29597;
  wire        _GEN_32574 = _GEN_1425 ? ~_GEN_1436 & _GEN_29598 : ~_GEN_1403 & _GEN_29598;
  wire        _GEN_32575 = _GEN_1425 ? ~_GEN_1437 & _GEN_29599 : ~_GEN_1404 & _GEN_29599;
  wire        _GEN_32576 = _GEN_1425 ? ~_GEN_1438 & _GEN_29600 : ~_GEN_1405 & _GEN_29600;
  wire        _GEN_32577 = _GEN_1425 ? ~_GEN_1439 & _GEN_29601 : ~_GEN_1406 & _GEN_29601;
  wire        _GEN_32578 = _GEN_1425 ? ~_GEN_1440 & _GEN_29602 : ~_GEN_1407 & _GEN_29602;
  wire        _GEN_32579 = _GEN_1425 ? ~_GEN_1441 & _GEN_29603 : ~_GEN_1408 & _GEN_29603;
  wire        _GEN_32580 = _GEN_1425 ? ~_GEN_1442 & _GEN_29604 : ~_GEN_1409 & _GEN_29604;
  wire        _GEN_32581 = _GEN_1425 ? ~_GEN_1443 & _GEN_29605 : ~_GEN_1410 & _GEN_29605;
  wire        _GEN_32582 = _GEN_1425 ? ~_GEN_1444 & _GEN_29606 : ~_GEN_1411 & _GEN_29606;
  wire        _GEN_32583 = _GEN_1425 ? ~_GEN_1445 & _GEN_29607 : ~_GEN_1412 & _GEN_29607;
  wire        _GEN_32584 = _GEN_1425 ? ~_GEN_1446 & _GEN_29608 : ~_GEN_1413 & _GEN_29608;
  wire        _GEN_32585 = _GEN_1425 ? ~_GEN_1447 & _GEN_29609 : ~_GEN_1414 & _GEN_29609;
  wire        _GEN_32586 = _GEN_1425 ? ~_GEN_1448 & _GEN_29610 : ~_GEN_1415 & _GEN_29610;
  wire        _GEN_32587 = _GEN_1425 ? ~_GEN_1449 & _GEN_29611 : ~_GEN_1416 & _GEN_29611;
  wire        _GEN_32588 = _GEN_1425 ? ~_GEN_1450 & _GEN_29612 : ~_GEN_1417 & _GEN_29612;
  wire        _GEN_32589 = _GEN_1425 ? ~_GEN_1451 & _GEN_29613 : ~_GEN_1418 & _GEN_29613;
  wire        _GEN_32590 = _GEN_1425 ? ~_GEN_1452 & _GEN_29614 : ~_GEN_1419 & _GEN_29614;
  wire        _GEN_32591 = _GEN_1425 ? ~_GEN_1453 & _GEN_29615 : ~_GEN_1420 & _GEN_29615;
  wire        _GEN_32592 = _GEN_1425 ? ~_GEN_1454 & _GEN_29616 : ~_GEN_1421 & _GEN_29616;
  wire        _GEN_32593 = _GEN_1425 ? ~_GEN_1455 & _GEN_29617 : ~_GEN_1422 & _GEN_29617;
  wire        _GEN_32594 = _GEN_1425 ? ~_GEN_1456 & _GEN_29618 : ~_GEN_1423 & _GEN_29618;
  wire        _GEN_32595 = _GEN_1425 ? ~_GEN_1457 & _GEN_29619 : ~_GEN_1424 & _GEN_29619;
  wire        _GEN_32948 = _GEN_1491 ? ~_GEN_1492 & _GEN_32564 : ~_GEN_1459 & _GEN_32564;
  wire        _GEN_32949 = _GEN_1491 ? ~_GEN_1493 & _GEN_32565 : ~_GEN_1460 & _GEN_32565;
  wire        _GEN_32950 = _GEN_1491 ? ~_GEN_1494 & _GEN_32566 : ~_GEN_1461 & _GEN_32566;
  wire        _GEN_32951 = _GEN_1491 ? ~_GEN_1495 & _GEN_32567 : ~_GEN_1462 & _GEN_32567;
  wire        _GEN_32952 = _GEN_1491 ? ~_GEN_1496 & _GEN_32568 : ~_GEN_1463 & _GEN_32568;
  wire        _GEN_32953 = _GEN_1491 ? ~_GEN_1497 & _GEN_32569 : ~_GEN_1464 & _GEN_32569;
  wire        _GEN_32954 = _GEN_1491 ? ~_GEN_1498 & _GEN_32570 : ~_GEN_1465 & _GEN_32570;
  wire        _GEN_32955 = _GEN_1491 ? ~_GEN_1499 & _GEN_32571 : ~_GEN_1466 & _GEN_32571;
  wire        _GEN_32956 = _GEN_1491 ? ~_GEN_1500 & _GEN_32572 : ~_GEN_1467 & _GEN_32572;
  wire        _GEN_32957 = _GEN_1491 ? ~_GEN_1501 & _GEN_32573 : ~_GEN_1468 & _GEN_32573;
  wire        _GEN_32958 = _GEN_1491 ? ~_GEN_1502 & _GEN_32574 : ~_GEN_1469 & _GEN_32574;
  wire        _GEN_32959 = _GEN_1491 ? ~_GEN_1503 & _GEN_32575 : ~_GEN_1470 & _GEN_32575;
  wire        _GEN_32960 = _GEN_1491 ? ~_GEN_1504 & _GEN_32576 : ~_GEN_1471 & _GEN_32576;
  wire        _GEN_32961 = _GEN_1491 ? ~_GEN_1505 & _GEN_32577 : ~_GEN_1472 & _GEN_32577;
  wire        _GEN_32962 = _GEN_1491 ? ~_GEN_1506 & _GEN_32578 : ~_GEN_1473 & _GEN_32578;
  wire        _GEN_32963 = _GEN_1491 ? ~_GEN_1507 & _GEN_32579 : ~_GEN_1474 & _GEN_32579;
  wire        _GEN_32964 = _GEN_1491 ? ~_GEN_1508 & _GEN_32580 : ~_GEN_1475 & _GEN_32580;
  wire        _GEN_32965 = _GEN_1491 ? ~_GEN_1509 & _GEN_32581 : ~_GEN_1476 & _GEN_32581;
  wire        _GEN_32966 = _GEN_1491 ? ~_GEN_1510 & _GEN_32582 : ~_GEN_1477 & _GEN_32582;
  wire        _GEN_32967 = _GEN_1491 ? ~_GEN_1511 & _GEN_32583 : ~_GEN_1478 & _GEN_32583;
  wire        _GEN_32968 = _GEN_1491 ? ~_GEN_1512 & _GEN_32584 : ~_GEN_1479 & _GEN_32584;
  wire        _GEN_32969 = _GEN_1491 ? ~_GEN_1513 & _GEN_32585 : ~_GEN_1480 & _GEN_32585;
  wire        _GEN_32970 = _GEN_1491 ? ~_GEN_1514 & _GEN_32586 : ~_GEN_1481 & _GEN_32586;
  wire        _GEN_32971 = _GEN_1491 ? ~_GEN_1515 & _GEN_32587 : ~_GEN_1482 & _GEN_32587;
  wire        _GEN_32972 = _GEN_1491 ? ~_GEN_1516 & _GEN_32588 : ~_GEN_1483 & _GEN_32588;
  wire        _GEN_32973 = _GEN_1491 ? ~_GEN_1517 & _GEN_32589 : ~_GEN_1484 & _GEN_32589;
  wire        _GEN_32974 = _GEN_1491 ? ~_GEN_1518 & _GEN_32590 : ~_GEN_1485 & _GEN_32590;
  wire        _GEN_32975 = _GEN_1491 ? ~_GEN_1519 & _GEN_32591 : ~_GEN_1486 & _GEN_32591;
  wire        _GEN_32976 = _GEN_1491 ? ~_GEN_1520 & _GEN_32592 : ~_GEN_1487 & _GEN_32592;
  wire        _GEN_32977 = _GEN_1491 ? ~_GEN_1521 & _GEN_32593 : ~_GEN_1488 & _GEN_32593;
  wire        _GEN_32978 = _GEN_1491 ? ~_GEN_1522 & _GEN_32594 : ~_GEN_1489 & _GEN_32594;
  wire        _GEN_32979 = _GEN_1491 ? ~_GEN_1523 & _GEN_32595 : ~_GEN_1490 & _GEN_32595;
  wire        _GEN_33332 = _GEN_1557 ? ~_GEN_1558 & _GEN_32948 : ~_GEN_1525 & _GEN_32948;
  wire        _GEN_33333 = _GEN_1557 ? ~_GEN_1559 & _GEN_32949 : ~_GEN_1526 & _GEN_32949;
  wire        _GEN_33334 = _GEN_1557 ? ~_GEN_1560 & _GEN_32950 : ~_GEN_1527 & _GEN_32950;
  wire        _GEN_33335 = _GEN_1557 ? ~_GEN_1561 & _GEN_32951 : ~_GEN_1528 & _GEN_32951;
  wire        _GEN_33336 = _GEN_1557 ? ~_GEN_1562 & _GEN_32952 : ~_GEN_1529 & _GEN_32952;
  wire        _GEN_33337 = _GEN_1557 ? ~_GEN_1563 & _GEN_32953 : ~_GEN_1530 & _GEN_32953;
  wire        _GEN_33338 = _GEN_1557 ? ~_GEN_1564 & _GEN_32954 : ~_GEN_1531 & _GEN_32954;
  wire        _GEN_33339 = _GEN_1557 ? ~_GEN_1565 & _GEN_32955 : ~_GEN_1532 & _GEN_32955;
  wire        _GEN_33340 = _GEN_1557 ? ~_GEN_1566 & _GEN_32956 : ~_GEN_1533 & _GEN_32956;
  wire        _GEN_33341 = _GEN_1557 ? ~_GEN_1567 & _GEN_32957 : ~_GEN_1534 & _GEN_32957;
  wire        _GEN_33342 = _GEN_1557 ? ~_GEN_1568 & _GEN_32958 : ~_GEN_1535 & _GEN_32958;
  wire        _GEN_33343 = _GEN_1557 ? ~_GEN_1569 & _GEN_32959 : ~_GEN_1536 & _GEN_32959;
  wire        _GEN_33344 = _GEN_1557 ? ~_GEN_1570 & _GEN_32960 : ~_GEN_1537 & _GEN_32960;
  wire        _GEN_33345 = _GEN_1557 ? ~_GEN_1571 & _GEN_32961 : ~_GEN_1538 & _GEN_32961;
  wire        _GEN_33346 = _GEN_1557 ? ~_GEN_1572 & _GEN_32962 : ~_GEN_1539 & _GEN_32962;
  wire        _GEN_33347 = _GEN_1557 ? ~_GEN_1573 & _GEN_32963 : ~_GEN_1540 & _GEN_32963;
  wire        _GEN_33348 = _GEN_1557 ? ~_GEN_1574 & _GEN_32964 : ~_GEN_1541 & _GEN_32964;
  wire        _GEN_33349 = _GEN_1557 ? ~_GEN_1575 & _GEN_32965 : ~_GEN_1542 & _GEN_32965;
  wire        _GEN_33350 = _GEN_1557 ? ~_GEN_1576 & _GEN_32966 : ~_GEN_1543 & _GEN_32966;
  wire        _GEN_33351 = _GEN_1557 ? ~_GEN_1577 & _GEN_32967 : ~_GEN_1544 & _GEN_32967;
  wire        _GEN_33352 = _GEN_1557 ? ~_GEN_1578 & _GEN_32968 : ~_GEN_1545 & _GEN_32968;
  wire        _GEN_33353 = _GEN_1557 ? ~_GEN_1579 & _GEN_32969 : ~_GEN_1546 & _GEN_32969;
  wire        _GEN_33354 = _GEN_1557 ? ~_GEN_1580 & _GEN_32970 : ~_GEN_1547 & _GEN_32970;
  wire        _GEN_33355 = _GEN_1557 ? ~_GEN_1581 & _GEN_32971 : ~_GEN_1548 & _GEN_32971;
  wire        _GEN_33356 = _GEN_1557 ? ~_GEN_1582 & _GEN_32972 : ~_GEN_1549 & _GEN_32972;
  wire        _GEN_33357 = _GEN_1557 ? ~_GEN_1583 & _GEN_32973 : ~_GEN_1550 & _GEN_32973;
  wire        _GEN_33358 = _GEN_1557 ? ~_GEN_1584 & _GEN_32974 : ~_GEN_1551 & _GEN_32974;
  wire        _GEN_33359 = _GEN_1557 ? ~_GEN_1585 & _GEN_32975 : ~_GEN_1552 & _GEN_32975;
  wire        _GEN_33360 = _GEN_1557 ? ~_GEN_1586 & _GEN_32976 : ~_GEN_1553 & _GEN_32976;
  wire        _GEN_33361 = _GEN_1557 ? ~_GEN_1587 & _GEN_32977 : ~_GEN_1554 & _GEN_32977;
  wire        _GEN_33362 = _GEN_1557 ? ~_GEN_1588 & _GEN_32978 : ~_GEN_1555 & _GEN_32978;
  wire        _GEN_33363 = _GEN_1557 ? ~_GEN_1589 & _GEN_32979 : ~_GEN_1556 & _GEN_32979;
  wire        _GEN_33716 = _GEN_1623 ? ~_GEN_1624 & _GEN_33332 : ~_GEN_1591 & _GEN_33332;
  wire        _GEN_33717 = _GEN_1623 ? ~_GEN_1625 & _GEN_33333 : ~_GEN_1592 & _GEN_33333;
  wire        _GEN_33718 = _GEN_1623 ? ~_GEN_1626 & _GEN_33334 : ~_GEN_1593 & _GEN_33334;
  wire        _GEN_33719 = _GEN_1623 ? ~_GEN_1627 & _GEN_33335 : ~_GEN_1594 & _GEN_33335;
  wire        _GEN_33720 = _GEN_1623 ? ~_GEN_1628 & _GEN_33336 : ~_GEN_1595 & _GEN_33336;
  wire        _GEN_33721 = _GEN_1623 ? ~_GEN_1629 & _GEN_33337 : ~_GEN_1596 & _GEN_33337;
  wire        _GEN_33722 = _GEN_1623 ? ~_GEN_1630 & _GEN_33338 : ~_GEN_1597 & _GEN_33338;
  wire        _GEN_33723 = _GEN_1623 ? ~_GEN_1631 & _GEN_33339 : ~_GEN_1598 & _GEN_33339;
  wire        _GEN_33724 = _GEN_1623 ? ~_GEN_1632 & _GEN_33340 : ~_GEN_1599 & _GEN_33340;
  wire        _GEN_33725 = _GEN_1623 ? ~_GEN_1633 & _GEN_33341 : ~_GEN_1600 & _GEN_33341;
  wire        _GEN_33726 = _GEN_1623 ? ~_GEN_1634 & _GEN_33342 : ~_GEN_1601 & _GEN_33342;
  wire        _GEN_33727 = _GEN_1623 ? ~_GEN_1635 & _GEN_33343 : ~_GEN_1602 & _GEN_33343;
  wire        _GEN_33728 = _GEN_1623 ? ~_GEN_1636 & _GEN_33344 : ~_GEN_1603 & _GEN_33344;
  wire        _GEN_33729 = _GEN_1623 ? ~_GEN_1637 & _GEN_33345 : ~_GEN_1604 & _GEN_33345;
  wire        _GEN_33730 = _GEN_1623 ? ~_GEN_1638 & _GEN_33346 : ~_GEN_1605 & _GEN_33346;
  wire        _GEN_33731 = _GEN_1623 ? ~_GEN_1639 & _GEN_33347 : ~_GEN_1606 & _GEN_33347;
  wire        _GEN_33732 = _GEN_1623 ? ~_GEN_1640 & _GEN_33348 : ~_GEN_1607 & _GEN_33348;
  wire        _GEN_33733 = _GEN_1623 ? ~_GEN_1641 & _GEN_33349 : ~_GEN_1608 & _GEN_33349;
  wire        _GEN_33734 = _GEN_1623 ? ~_GEN_1642 & _GEN_33350 : ~_GEN_1609 & _GEN_33350;
  wire        _GEN_33735 = _GEN_1623 ? ~_GEN_1643 & _GEN_33351 : ~_GEN_1610 & _GEN_33351;
  wire        _GEN_33736 = _GEN_1623 ? ~_GEN_1644 & _GEN_33352 : ~_GEN_1611 & _GEN_33352;
  wire        _GEN_33737 = _GEN_1623 ? ~_GEN_1645 & _GEN_33353 : ~_GEN_1612 & _GEN_33353;
  wire        _GEN_33738 = _GEN_1623 ? ~_GEN_1646 & _GEN_33354 : ~_GEN_1613 & _GEN_33354;
  wire        _GEN_33739 = _GEN_1623 ? ~_GEN_1647 & _GEN_33355 : ~_GEN_1614 & _GEN_33355;
  wire        _GEN_33740 = _GEN_1623 ? ~_GEN_1648 & _GEN_33356 : ~_GEN_1615 & _GEN_33356;
  wire        _GEN_33741 = _GEN_1623 ? ~_GEN_1649 & _GEN_33357 : ~_GEN_1616 & _GEN_33357;
  wire        _GEN_33742 = _GEN_1623 ? ~_GEN_1650 & _GEN_33358 : ~_GEN_1617 & _GEN_33358;
  wire        _GEN_33743 = _GEN_1623 ? ~_GEN_1651 & _GEN_33359 : ~_GEN_1618 & _GEN_33359;
  wire        _GEN_33744 = _GEN_1623 ? ~_GEN_1652 & _GEN_33360 : ~_GEN_1619 & _GEN_33360;
  wire        _GEN_33745 = _GEN_1623 ? ~_GEN_1653 & _GEN_33361 : ~_GEN_1620 & _GEN_33361;
  wire        _GEN_33746 = _GEN_1623 ? ~_GEN_1654 & _GEN_33362 : ~_GEN_1621 & _GEN_33362;
  wire        _GEN_33747 = _GEN_1623 ? ~_GEN_1655 & _GEN_33363 : ~_GEN_1622 & _GEN_33363;
  wire        _GEN_34100 = _GEN_1689 ? ~_GEN_1690 & _GEN_33716 : ~_GEN_1657 & _GEN_33716;
  wire        _GEN_34101 = _GEN_1689 ? ~_GEN_1691 & _GEN_33717 : ~_GEN_1658 & _GEN_33717;
  wire        _GEN_34102 = _GEN_1689 ? ~_GEN_1692 & _GEN_33718 : ~_GEN_1659 & _GEN_33718;
  wire        _GEN_34103 = _GEN_1689 ? ~_GEN_1693 & _GEN_33719 : ~_GEN_1660 & _GEN_33719;
  wire        _GEN_34104 = _GEN_1689 ? ~_GEN_1694 & _GEN_33720 : ~_GEN_1661 & _GEN_33720;
  wire        _GEN_34105 = _GEN_1689 ? ~_GEN_1695 & _GEN_33721 : ~_GEN_1662 & _GEN_33721;
  wire        _GEN_34106 = _GEN_1689 ? ~_GEN_1696 & _GEN_33722 : ~_GEN_1663 & _GEN_33722;
  wire        _GEN_34107 = _GEN_1689 ? ~_GEN_1697 & _GEN_33723 : ~_GEN_1664 & _GEN_33723;
  wire        _GEN_34108 = _GEN_1689 ? ~_GEN_1698 & _GEN_33724 : ~_GEN_1665 & _GEN_33724;
  wire        _GEN_34109 = _GEN_1689 ? ~_GEN_1699 & _GEN_33725 : ~_GEN_1666 & _GEN_33725;
  wire        _GEN_34110 = _GEN_1689 ? ~_GEN_1700 & _GEN_33726 : ~_GEN_1667 & _GEN_33726;
  wire        _GEN_34111 = _GEN_1689 ? ~_GEN_1701 & _GEN_33727 : ~_GEN_1668 & _GEN_33727;
  wire        _GEN_34112 = _GEN_1689 ? ~_GEN_1702 & _GEN_33728 : ~_GEN_1669 & _GEN_33728;
  wire        _GEN_34113 = _GEN_1689 ? ~_GEN_1703 & _GEN_33729 : ~_GEN_1670 & _GEN_33729;
  wire        _GEN_34114 = _GEN_1689 ? ~_GEN_1704 & _GEN_33730 : ~_GEN_1671 & _GEN_33730;
  wire        _GEN_34115 = _GEN_1689 ? ~_GEN_1705 & _GEN_33731 : ~_GEN_1672 & _GEN_33731;
  wire        _GEN_34116 = _GEN_1689 ? ~_GEN_1706 & _GEN_33732 : ~_GEN_1673 & _GEN_33732;
  wire        _GEN_34117 = _GEN_1689 ? ~_GEN_1707 & _GEN_33733 : ~_GEN_1674 & _GEN_33733;
  wire        _GEN_34118 = _GEN_1689 ? ~_GEN_1708 & _GEN_33734 : ~_GEN_1675 & _GEN_33734;
  wire        _GEN_34119 = _GEN_1689 ? ~_GEN_1709 & _GEN_33735 : ~_GEN_1676 & _GEN_33735;
  wire        _GEN_34120 = _GEN_1689 ? ~_GEN_1710 & _GEN_33736 : ~_GEN_1677 & _GEN_33736;
  wire        _GEN_34121 = _GEN_1689 ? ~_GEN_1711 & _GEN_33737 : ~_GEN_1678 & _GEN_33737;
  wire        _GEN_34122 = _GEN_1689 ? ~_GEN_1712 & _GEN_33738 : ~_GEN_1679 & _GEN_33738;
  wire        _GEN_34123 = _GEN_1689 ? ~_GEN_1713 & _GEN_33739 : ~_GEN_1680 & _GEN_33739;
  wire        _GEN_34124 = _GEN_1689 ? ~_GEN_1714 & _GEN_33740 : ~_GEN_1681 & _GEN_33740;
  wire        _GEN_34125 = _GEN_1689 ? ~_GEN_1715 & _GEN_33741 : ~_GEN_1682 & _GEN_33741;
  wire        _GEN_34126 = _GEN_1689 ? ~_GEN_1716 & _GEN_33742 : ~_GEN_1683 & _GEN_33742;
  wire        _GEN_34127 = _GEN_1689 ? ~_GEN_1717 & _GEN_33743 : ~_GEN_1684 & _GEN_33743;
  wire        _GEN_34128 = _GEN_1689 ? ~_GEN_1718 & _GEN_33744 : ~_GEN_1685 & _GEN_33744;
  wire        _GEN_34129 = _GEN_1689 ? ~_GEN_1719 & _GEN_33745 : ~_GEN_1686 & _GEN_33745;
  wire        _GEN_34130 = _GEN_1689 ? ~_GEN_1720 & _GEN_33746 : ~_GEN_1687 & _GEN_33746;
  wire        _GEN_34131 = _GEN_1689 ? ~_GEN_1721 & _GEN_33747 : ~_GEN_1688 & _GEN_33747;
  wire        _GEN_2609 = io_fflags_0_valid & io_fflags_0_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_2610 = io_fflags_2_valid & io_fflags_2_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_2611 = io_fflags_3_valid & io_fflags_3_bits_uop_rob_idx[1:0] == 2'h2;
  wire        _GEN_2612 = rbk_row_2 & _GEN_2477;
  wire        _GEN_2613 = rbk_row_2 & _GEN_2447;
  wire        _GEN_2614 = rbk_row_2 & _GEN_2448;
  wire        _GEN_2615 = rbk_row_2 & _GEN_2449;
  wire        _GEN_2616 = rbk_row_2 & _GEN_2450;
  wire        _GEN_2617 = rbk_row_2 & _GEN_2451;
  wire        _GEN_2618 = rbk_row_2 & _GEN_2452;
  wire        _GEN_2619 = rbk_row_2 & _GEN_2453;
  wire        _GEN_2620 = rbk_row_2 & _GEN_2454;
  wire        _GEN_2621 = rbk_row_2 & _GEN_2455;
  wire        _GEN_2622 = rbk_row_2 & _GEN_2456;
  wire        _GEN_2623 = rbk_row_2 & _GEN_2457;
  wire        _GEN_2624 = rbk_row_2 & _GEN_2458;
  wire        _GEN_2625 = rbk_row_2 & _GEN_2459;
  wire        _GEN_2626 = rbk_row_2 & _GEN_2460;
  wire        _GEN_2627 = rbk_row_2 & _GEN_2461;
  wire        _GEN_2628 = rbk_row_2 & _GEN_2462;
  wire        _GEN_2629 = rbk_row_2 & _GEN_2463;
  wire        _GEN_2630 = rbk_row_2 & _GEN_2464;
  wire        _GEN_2631 = rbk_row_2 & _GEN_2465;
  wire        _GEN_2632 = rbk_row_2 & _GEN_2466;
  wire        _GEN_2633 = rbk_row_2 & _GEN_2467;
  wire        _GEN_2634 = rbk_row_2 & _GEN_2468;
  wire        _GEN_2635 = rbk_row_2 & _GEN_2469;
  wire        _GEN_2636 = rbk_row_2 & _GEN_2470;
  wire        _GEN_2637 = rbk_row_2 & _GEN_2471;
  wire        _GEN_2638 = rbk_row_2 & _GEN_2472;
  wire        _GEN_2639 = rbk_row_2 & _GEN_2473;
  wire        _GEN_2640 = rbk_row_2 & _GEN_2474;
  wire        _GEN_2641 = rbk_row_2 & _GEN_2475;
  wire        _GEN_2642 = rbk_row_2 & _GEN_2476;
  wire        _GEN_2643 = rbk_row_2 & (&com_idx);
  wire [19:0] _GEN_2644 = io_brupdate_b1_mispredict_mask & rob_uop_2_0_br_mask;
  wire [19:0] _GEN_2645 = io_brupdate_b1_mispredict_mask & rob_uop_2_1_br_mask;
  wire [19:0] _GEN_2646 = io_brupdate_b1_mispredict_mask & rob_uop_2_2_br_mask;
  wire [19:0] _GEN_2647 = io_brupdate_b1_mispredict_mask & rob_uop_2_3_br_mask;
  wire [19:0] _GEN_2648 = io_brupdate_b1_mispredict_mask & rob_uop_2_4_br_mask;
  wire [19:0] _GEN_2649 = io_brupdate_b1_mispredict_mask & rob_uop_2_5_br_mask;
  wire [19:0] _GEN_2650 = io_brupdate_b1_mispredict_mask & rob_uop_2_6_br_mask;
  wire [19:0] _GEN_2651 = io_brupdate_b1_mispredict_mask & rob_uop_2_7_br_mask;
  wire [19:0] _GEN_2652 = io_brupdate_b1_mispredict_mask & rob_uop_2_8_br_mask;
  wire [19:0] _GEN_2653 = io_brupdate_b1_mispredict_mask & rob_uop_2_9_br_mask;
  wire [19:0] _GEN_2654 = io_brupdate_b1_mispredict_mask & rob_uop_2_10_br_mask;
  wire [19:0] _GEN_2655 = io_brupdate_b1_mispredict_mask & rob_uop_2_11_br_mask;
  wire [19:0] _GEN_2656 = io_brupdate_b1_mispredict_mask & rob_uop_2_12_br_mask;
  wire [19:0] _GEN_2657 = io_brupdate_b1_mispredict_mask & rob_uop_2_13_br_mask;
  wire [19:0] _GEN_2658 = io_brupdate_b1_mispredict_mask & rob_uop_2_14_br_mask;
  wire [19:0] _GEN_2659 = io_brupdate_b1_mispredict_mask & rob_uop_2_15_br_mask;
  wire [19:0] _GEN_2660 = io_brupdate_b1_mispredict_mask & rob_uop_2_16_br_mask;
  wire [19:0] _GEN_2661 = io_brupdate_b1_mispredict_mask & rob_uop_2_17_br_mask;
  wire [19:0] _GEN_2662 = io_brupdate_b1_mispredict_mask & rob_uop_2_18_br_mask;
  wire [19:0] _GEN_2663 = io_brupdate_b1_mispredict_mask & rob_uop_2_19_br_mask;
  wire [19:0] _GEN_2664 = io_brupdate_b1_mispredict_mask & rob_uop_2_20_br_mask;
  wire [19:0] _GEN_2665 = io_brupdate_b1_mispredict_mask & rob_uop_2_21_br_mask;
  wire [19:0] _GEN_2666 = io_brupdate_b1_mispredict_mask & rob_uop_2_22_br_mask;
  wire [19:0] _GEN_2667 = io_brupdate_b1_mispredict_mask & rob_uop_2_23_br_mask;
  wire [19:0] _GEN_2668 = io_brupdate_b1_mispredict_mask & rob_uop_2_24_br_mask;
  wire [19:0] _GEN_2669 = io_brupdate_b1_mispredict_mask & rob_uop_2_25_br_mask;
  wire [19:0] _GEN_2670 = io_brupdate_b1_mispredict_mask & rob_uop_2_26_br_mask;
  wire [19:0] _GEN_2671 = io_brupdate_b1_mispredict_mask & rob_uop_2_27_br_mask;
  wire [19:0] _GEN_2672 = io_brupdate_b1_mispredict_mask & rob_uop_2_28_br_mask;
  wire [19:0] _GEN_2673 = io_brupdate_b1_mispredict_mask & rob_uop_2_29_br_mask;
  wire [19:0] _GEN_2674 = io_brupdate_b1_mispredict_mask & rob_uop_2_30_br_mask;
  wire [19:0] _GEN_2675 = io_brupdate_b1_mispredict_mask & rob_uop_2_31_br_mask;
  wire        _rob_bsy_T_6 = io_enq_uops_3_is_fence | io_enq_uops_3_is_fencei;
  wire        _GEN_42952 = _GEN_1822 ? ~_rob_bsy_T_6 : rob_bsy_3_0;
  wire        _GEN_42953 = _GEN_1823 ? ~_rob_bsy_T_6 : rob_bsy_3_1;
  wire        _GEN_42954 = _GEN_1824 ? ~_rob_bsy_T_6 : rob_bsy_3_2;
  wire        _GEN_42955 = _GEN_1825 ? ~_rob_bsy_T_6 : rob_bsy_3_3;
  wire        _GEN_42956 = _GEN_1826 ? ~_rob_bsy_T_6 : rob_bsy_3_4;
  wire        _GEN_42957 = _GEN_1827 ? ~_rob_bsy_T_6 : rob_bsy_3_5;
  wire        _GEN_42958 = _GEN_1828 ? ~_rob_bsy_T_6 : rob_bsy_3_6;
  wire        _GEN_42959 = _GEN_1829 ? ~_rob_bsy_T_6 : rob_bsy_3_7;
  wire        _GEN_42960 = _GEN_1830 ? ~_rob_bsy_T_6 : rob_bsy_3_8;
  wire        _GEN_42961 = _GEN_1831 ? ~_rob_bsy_T_6 : rob_bsy_3_9;
  wire        _GEN_42962 = _GEN_1832 ? ~_rob_bsy_T_6 : rob_bsy_3_10;
  wire        _GEN_42963 = _GEN_1833 ? ~_rob_bsy_T_6 : rob_bsy_3_11;
  wire        _GEN_42964 = _GEN_1834 ? ~_rob_bsy_T_6 : rob_bsy_3_12;
  wire        _GEN_42965 = _GEN_1835 ? ~_rob_bsy_T_6 : rob_bsy_3_13;
  wire        _GEN_42966 = _GEN_1836 ? ~_rob_bsy_T_6 : rob_bsy_3_14;
  wire        _GEN_42967 = _GEN_1837 ? ~_rob_bsy_T_6 : rob_bsy_3_15;
  wire        _GEN_42968 = _GEN_1838 ? ~_rob_bsy_T_6 : rob_bsy_3_16;
  wire        _GEN_42969 = _GEN_1839 ? ~_rob_bsy_T_6 : rob_bsy_3_17;
  wire        _GEN_42970 = _GEN_1840 ? ~_rob_bsy_T_6 : rob_bsy_3_18;
  wire        _GEN_42971 = _GEN_1841 ? ~_rob_bsy_T_6 : rob_bsy_3_19;
  wire        _GEN_42972 = _GEN_1842 ? ~_rob_bsy_T_6 : rob_bsy_3_20;
  wire        _GEN_42973 = _GEN_1843 ? ~_rob_bsy_T_6 : rob_bsy_3_21;
  wire        _GEN_42974 = _GEN_1844 ? ~_rob_bsy_T_6 : rob_bsy_3_22;
  wire        _GEN_42975 = _GEN_1845 ? ~_rob_bsy_T_6 : rob_bsy_3_23;
  wire        _GEN_42976 = _GEN_1846 ? ~_rob_bsy_T_6 : rob_bsy_3_24;
  wire        _GEN_42977 = _GEN_1847 ? ~_rob_bsy_T_6 : rob_bsy_3_25;
  wire        _GEN_42978 = _GEN_1848 ? ~_rob_bsy_T_6 : rob_bsy_3_26;
  wire        _GEN_42979 = _GEN_1849 ? ~_rob_bsy_T_6 : rob_bsy_3_27;
  wire        _GEN_42980 = _GEN_1850 ? ~_rob_bsy_T_6 : rob_bsy_3_28;
  wire        _GEN_42981 = _GEN_1851 ? ~_rob_bsy_T_6 : rob_bsy_3_29;
  wire        _GEN_42982 = _GEN_1852 ? ~_rob_bsy_T_6 : rob_bsy_3_30;
  wire        _GEN_42983 = _GEN_1853 ? ~_rob_bsy_T_6 : rob_bsy_3_31;
  wire        _GEN_45928 = _GEN_1887 ? ~_GEN_1888 & _GEN_42952 : ~_GEN_1855 & _GEN_42952;
  wire        _GEN_45929 = _GEN_1887 ? ~_GEN_1889 & _GEN_42953 : ~_GEN_1856 & _GEN_42953;
  wire        _GEN_45930 = _GEN_1887 ? ~_GEN_1890 & _GEN_42954 : ~_GEN_1857 & _GEN_42954;
  wire        _GEN_45931 = _GEN_1887 ? ~_GEN_1891 & _GEN_42955 : ~_GEN_1858 & _GEN_42955;
  wire        _GEN_45932 = _GEN_1887 ? ~_GEN_1892 & _GEN_42956 : ~_GEN_1859 & _GEN_42956;
  wire        _GEN_45933 = _GEN_1887 ? ~_GEN_1893 & _GEN_42957 : ~_GEN_1860 & _GEN_42957;
  wire        _GEN_45934 = _GEN_1887 ? ~_GEN_1894 & _GEN_42958 : ~_GEN_1861 & _GEN_42958;
  wire        _GEN_45935 = _GEN_1887 ? ~_GEN_1895 & _GEN_42959 : ~_GEN_1862 & _GEN_42959;
  wire        _GEN_45936 = _GEN_1887 ? ~_GEN_1896 & _GEN_42960 : ~_GEN_1863 & _GEN_42960;
  wire        _GEN_45937 = _GEN_1887 ? ~_GEN_1897 & _GEN_42961 : ~_GEN_1864 & _GEN_42961;
  wire        _GEN_45938 = _GEN_1887 ? ~_GEN_1898 & _GEN_42962 : ~_GEN_1865 & _GEN_42962;
  wire        _GEN_45939 = _GEN_1887 ? ~_GEN_1899 & _GEN_42963 : ~_GEN_1866 & _GEN_42963;
  wire        _GEN_45940 = _GEN_1887 ? ~_GEN_1900 & _GEN_42964 : ~_GEN_1867 & _GEN_42964;
  wire        _GEN_45941 = _GEN_1887 ? ~_GEN_1901 & _GEN_42965 : ~_GEN_1868 & _GEN_42965;
  wire        _GEN_45942 = _GEN_1887 ? ~_GEN_1902 & _GEN_42966 : ~_GEN_1869 & _GEN_42966;
  wire        _GEN_45943 = _GEN_1887 ? ~_GEN_1903 & _GEN_42967 : ~_GEN_1870 & _GEN_42967;
  wire        _GEN_45944 = _GEN_1887 ? ~_GEN_1904 & _GEN_42968 : ~_GEN_1871 & _GEN_42968;
  wire        _GEN_45945 = _GEN_1887 ? ~_GEN_1905 & _GEN_42969 : ~_GEN_1872 & _GEN_42969;
  wire        _GEN_45946 = _GEN_1887 ? ~_GEN_1906 & _GEN_42970 : ~_GEN_1873 & _GEN_42970;
  wire        _GEN_45947 = _GEN_1887 ? ~_GEN_1907 & _GEN_42971 : ~_GEN_1874 & _GEN_42971;
  wire        _GEN_45948 = _GEN_1887 ? ~_GEN_1908 & _GEN_42972 : ~_GEN_1875 & _GEN_42972;
  wire        _GEN_45949 = _GEN_1887 ? ~_GEN_1909 & _GEN_42973 : ~_GEN_1876 & _GEN_42973;
  wire        _GEN_45950 = _GEN_1887 ? ~_GEN_1910 & _GEN_42974 : ~_GEN_1877 & _GEN_42974;
  wire        _GEN_45951 = _GEN_1887 ? ~_GEN_1911 & _GEN_42975 : ~_GEN_1878 & _GEN_42975;
  wire        _GEN_45952 = _GEN_1887 ? ~_GEN_1912 & _GEN_42976 : ~_GEN_1879 & _GEN_42976;
  wire        _GEN_45953 = _GEN_1887 ? ~_GEN_1913 & _GEN_42977 : ~_GEN_1880 & _GEN_42977;
  wire        _GEN_45954 = _GEN_1887 ? ~_GEN_1914 & _GEN_42978 : ~_GEN_1881 & _GEN_42978;
  wire        _GEN_45955 = _GEN_1887 ? ~_GEN_1915 & _GEN_42979 : ~_GEN_1882 & _GEN_42979;
  wire        _GEN_45956 = _GEN_1887 ? ~_GEN_1916 & _GEN_42980 : ~_GEN_1883 & _GEN_42980;
  wire        _GEN_45957 = _GEN_1887 ? ~_GEN_1917 & _GEN_42981 : ~_GEN_1884 & _GEN_42981;
  wire        _GEN_45958 = _GEN_1887 ? ~_GEN_1918 & _GEN_42982 : ~_GEN_1885 & _GEN_42982;
  wire        _GEN_45959 = _GEN_1887 ? ~_GEN_1919 & _GEN_42983 : ~_GEN_1886 & _GEN_42983;
  wire        _GEN_46312 = _GEN_1953 ? ~_GEN_1954 & _GEN_45928 : ~_GEN_1921 & _GEN_45928;
  wire        _GEN_46313 = _GEN_1953 ? ~_GEN_1955 & _GEN_45929 : ~_GEN_1922 & _GEN_45929;
  wire        _GEN_46314 = _GEN_1953 ? ~_GEN_1956 & _GEN_45930 : ~_GEN_1923 & _GEN_45930;
  wire        _GEN_46315 = _GEN_1953 ? ~_GEN_1957 & _GEN_45931 : ~_GEN_1924 & _GEN_45931;
  wire        _GEN_46316 = _GEN_1953 ? ~_GEN_1958 & _GEN_45932 : ~_GEN_1925 & _GEN_45932;
  wire        _GEN_46317 = _GEN_1953 ? ~_GEN_1959 & _GEN_45933 : ~_GEN_1926 & _GEN_45933;
  wire        _GEN_46318 = _GEN_1953 ? ~_GEN_1960 & _GEN_45934 : ~_GEN_1927 & _GEN_45934;
  wire        _GEN_46319 = _GEN_1953 ? ~_GEN_1961 & _GEN_45935 : ~_GEN_1928 & _GEN_45935;
  wire        _GEN_46320 = _GEN_1953 ? ~_GEN_1962 & _GEN_45936 : ~_GEN_1929 & _GEN_45936;
  wire        _GEN_46321 = _GEN_1953 ? ~_GEN_1963 & _GEN_45937 : ~_GEN_1930 & _GEN_45937;
  wire        _GEN_46322 = _GEN_1953 ? ~_GEN_1964 & _GEN_45938 : ~_GEN_1931 & _GEN_45938;
  wire        _GEN_46323 = _GEN_1953 ? ~_GEN_1965 & _GEN_45939 : ~_GEN_1932 & _GEN_45939;
  wire        _GEN_46324 = _GEN_1953 ? ~_GEN_1966 & _GEN_45940 : ~_GEN_1933 & _GEN_45940;
  wire        _GEN_46325 = _GEN_1953 ? ~_GEN_1967 & _GEN_45941 : ~_GEN_1934 & _GEN_45941;
  wire        _GEN_46326 = _GEN_1953 ? ~_GEN_1968 & _GEN_45942 : ~_GEN_1935 & _GEN_45942;
  wire        _GEN_46327 = _GEN_1953 ? ~_GEN_1969 & _GEN_45943 : ~_GEN_1936 & _GEN_45943;
  wire        _GEN_46328 = _GEN_1953 ? ~_GEN_1970 & _GEN_45944 : ~_GEN_1937 & _GEN_45944;
  wire        _GEN_46329 = _GEN_1953 ? ~_GEN_1971 & _GEN_45945 : ~_GEN_1938 & _GEN_45945;
  wire        _GEN_46330 = _GEN_1953 ? ~_GEN_1972 & _GEN_45946 : ~_GEN_1939 & _GEN_45946;
  wire        _GEN_46331 = _GEN_1953 ? ~_GEN_1973 & _GEN_45947 : ~_GEN_1940 & _GEN_45947;
  wire        _GEN_46332 = _GEN_1953 ? ~_GEN_1974 & _GEN_45948 : ~_GEN_1941 & _GEN_45948;
  wire        _GEN_46333 = _GEN_1953 ? ~_GEN_1975 & _GEN_45949 : ~_GEN_1942 & _GEN_45949;
  wire        _GEN_46334 = _GEN_1953 ? ~_GEN_1976 & _GEN_45950 : ~_GEN_1943 & _GEN_45950;
  wire        _GEN_46335 = _GEN_1953 ? ~_GEN_1977 & _GEN_45951 : ~_GEN_1944 & _GEN_45951;
  wire        _GEN_46336 = _GEN_1953 ? ~_GEN_1978 & _GEN_45952 : ~_GEN_1945 & _GEN_45952;
  wire        _GEN_46337 = _GEN_1953 ? ~_GEN_1979 & _GEN_45953 : ~_GEN_1946 & _GEN_45953;
  wire        _GEN_46338 = _GEN_1953 ? ~_GEN_1980 & _GEN_45954 : ~_GEN_1947 & _GEN_45954;
  wire        _GEN_46339 = _GEN_1953 ? ~_GEN_1981 & _GEN_45955 : ~_GEN_1948 & _GEN_45955;
  wire        _GEN_46340 = _GEN_1953 ? ~_GEN_1982 & _GEN_45956 : ~_GEN_1949 & _GEN_45956;
  wire        _GEN_46341 = _GEN_1953 ? ~_GEN_1983 & _GEN_45957 : ~_GEN_1950 & _GEN_45957;
  wire        _GEN_46342 = _GEN_1953 ? ~_GEN_1984 & _GEN_45958 : ~_GEN_1951 & _GEN_45958;
  wire        _GEN_46343 = _GEN_1953 ? ~_GEN_1985 & _GEN_45959 : ~_GEN_1952 & _GEN_45959;
  wire        _GEN_46696 = _GEN_2019 ? ~_GEN_2020 & _GEN_46312 : ~_GEN_1987 & _GEN_46312;
  wire        _GEN_46697 = _GEN_2019 ? ~_GEN_2021 & _GEN_46313 : ~_GEN_1988 & _GEN_46313;
  wire        _GEN_46698 = _GEN_2019 ? ~_GEN_2022 & _GEN_46314 : ~_GEN_1989 & _GEN_46314;
  wire        _GEN_46699 = _GEN_2019 ? ~_GEN_2023 & _GEN_46315 : ~_GEN_1990 & _GEN_46315;
  wire        _GEN_46700 = _GEN_2019 ? ~_GEN_2024 & _GEN_46316 : ~_GEN_1991 & _GEN_46316;
  wire        _GEN_46701 = _GEN_2019 ? ~_GEN_2025 & _GEN_46317 : ~_GEN_1992 & _GEN_46317;
  wire        _GEN_46702 = _GEN_2019 ? ~_GEN_2026 & _GEN_46318 : ~_GEN_1993 & _GEN_46318;
  wire        _GEN_46703 = _GEN_2019 ? ~_GEN_2027 & _GEN_46319 : ~_GEN_1994 & _GEN_46319;
  wire        _GEN_46704 = _GEN_2019 ? ~_GEN_2028 & _GEN_46320 : ~_GEN_1995 & _GEN_46320;
  wire        _GEN_46705 = _GEN_2019 ? ~_GEN_2029 & _GEN_46321 : ~_GEN_1996 & _GEN_46321;
  wire        _GEN_46706 = _GEN_2019 ? ~_GEN_2030 & _GEN_46322 : ~_GEN_1997 & _GEN_46322;
  wire        _GEN_46707 = _GEN_2019 ? ~_GEN_2031 & _GEN_46323 : ~_GEN_1998 & _GEN_46323;
  wire        _GEN_46708 = _GEN_2019 ? ~_GEN_2032 & _GEN_46324 : ~_GEN_1999 & _GEN_46324;
  wire        _GEN_46709 = _GEN_2019 ? ~_GEN_2033 & _GEN_46325 : ~_GEN_2000 & _GEN_46325;
  wire        _GEN_46710 = _GEN_2019 ? ~_GEN_2034 & _GEN_46326 : ~_GEN_2001 & _GEN_46326;
  wire        _GEN_46711 = _GEN_2019 ? ~_GEN_2035 & _GEN_46327 : ~_GEN_2002 & _GEN_46327;
  wire        _GEN_46712 = _GEN_2019 ? ~_GEN_2036 & _GEN_46328 : ~_GEN_2003 & _GEN_46328;
  wire        _GEN_46713 = _GEN_2019 ? ~_GEN_2037 & _GEN_46329 : ~_GEN_2004 & _GEN_46329;
  wire        _GEN_46714 = _GEN_2019 ? ~_GEN_2038 & _GEN_46330 : ~_GEN_2005 & _GEN_46330;
  wire        _GEN_46715 = _GEN_2019 ? ~_GEN_2039 & _GEN_46331 : ~_GEN_2006 & _GEN_46331;
  wire        _GEN_46716 = _GEN_2019 ? ~_GEN_2040 & _GEN_46332 : ~_GEN_2007 & _GEN_46332;
  wire        _GEN_46717 = _GEN_2019 ? ~_GEN_2041 & _GEN_46333 : ~_GEN_2008 & _GEN_46333;
  wire        _GEN_46718 = _GEN_2019 ? ~_GEN_2042 & _GEN_46334 : ~_GEN_2009 & _GEN_46334;
  wire        _GEN_46719 = _GEN_2019 ? ~_GEN_2043 & _GEN_46335 : ~_GEN_2010 & _GEN_46335;
  wire        _GEN_46720 = _GEN_2019 ? ~_GEN_2044 & _GEN_46336 : ~_GEN_2011 & _GEN_46336;
  wire        _GEN_46721 = _GEN_2019 ? ~_GEN_2045 & _GEN_46337 : ~_GEN_2012 & _GEN_46337;
  wire        _GEN_46722 = _GEN_2019 ? ~_GEN_2046 & _GEN_46338 : ~_GEN_2013 & _GEN_46338;
  wire        _GEN_46723 = _GEN_2019 ? ~_GEN_2047 & _GEN_46339 : ~_GEN_2014 & _GEN_46339;
  wire        _GEN_46724 = _GEN_2019 ? ~_GEN_2048 & _GEN_46340 : ~_GEN_2015 & _GEN_46340;
  wire        _GEN_46725 = _GEN_2019 ? ~_GEN_2049 & _GEN_46341 : ~_GEN_2016 & _GEN_46341;
  wire        _GEN_46726 = _GEN_2019 ? ~_GEN_2050 & _GEN_46342 : ~_GEN_2017 & _GEN_46342;
  wire        _GEN_46727 = _GEN_2019 ? ~_GEN_2051 & _GEN_46343 : ~_GEN_2018 & _GEN_46343;
  wire        _GEN_47080 = _GEN_2085 ? ~_GEN_2086 & _GEN_46696 : ~_GEN_2053 & _GEN_46696;
  wire        _GEN_47081 = _GEN_2085 ? ~_GEN_2087 & _GEN_46697 : ~_GEN_2054 & _GEN_46697;
  wire        _GEN_47082 = _GEN_2085 ? ~_GEN_2088 & _GEN_46698 : ~_GEN_2055 & _GEN_46698;
  wire        _GEN_47083 = _GEN_2085 ? ~_GEN_2089 & _GEN_46699 : ~_GEN_2056 & _GEN_46699;
  wire        _GEN_47084 = _GEN_2085 ? ~_GEN_2090 & _GEN_46700 : ~_GEN_2057 & _GEN_46700;
  wire        _GEN_47085 = _GEN_2085 ? ~_GEN_2091 & _GEN_46701 : ~_GEN_2058 & _GEN_46701;
  wire        _GEN_47086 = _GEN_2085 ? ~_GEN_2092 & _GEN_46702 : ~_GEN_2059 & _GEN_46702;
  wire        _GEN_47087 = _GEN_2085 ? ~_GEN_2093 & _GEN_46703 : ~_GEN_2060 & _GEN_46703;
  wire        _GEN_47088 = _GEN_2085 ? ~_GEN_2094 & _GEN_46704 : ~_GEN_2061 & _GEN_46704;
  wire        _GEN_47089 = _GEN_2085 ? ~_GEN_2095 & _GEN_46705 : ~_GEN_2062 & _GEN_46705;
  wire        _GEN_47090 = _GEN_2085 ? ~_GEN_2096 & _GEN_46706 : ~_GEN_2063 & _GEN_46706;
  wire        _GEN_47091 = _GEN_2085 ? ~_GEN_2097 & _GEN_46707 : ~_GEN_2064 & _GEN_46707;
  wire        _GEN_47092 = _GEN_2085 ? ~_GEN_2098 & _GEN_46708 : ~_GEN_2065 & _GEN_46708;
  wire        _GEN_47093 = _GEN_2085 ? ~_GEN_2099 & _GEN_46709 : ~_GEN_2066 & _GEN_46709;
  wire        _GEN_47094 = _GEN_2085 ? ~_GEN_2100 & _GEN_46710 : ~_GEN_2067 & _GEN_46710;
  wire        _GEN_47095 = _GEN_2085 ? ~_GEN_2101 & _GEN_46711 : ~_GEN_2068 & _GEN_46711;
  wire        _GEN_47096 = _GEN_2085 ? ~_GEN_2102 & _GEN_46712 : ~_GEN_2069 & _GEN_46712;
  wire        _GEN_47097 = _GEN_2085 ? ~_GEN_2103 & _GEN_46713 : ~_GEN_2070 & _GEN_46713;
  wire        _GEN_47098 = _GEN_2085 ? ~_GEN_2104 & _GEN_46714 : ~_GEN_2071 & _GEN_46714;
  wire        _GEN_47099 = _GEN_2085 ? ~_GEN_2105 & _GEN_46715 : ~_GEN_2072 & _GEN_46715;
  wire        _GEN_47100 = _GEN_2085 ? ~_GEN_2106 & _GEN_46716 : ~_GEN_2073 & _GEN_46716;
  wire        _GEN_47101 = _GEN_2085 ? ~_GEN_2107 & _GEN_46717 : ~_GEN_2074 & _GEN_46717;
  wire        _GEN_47102 = _GEN_2085 ? ~_GEN_2108 & _GEN_46718 : ~_GEN_2075 & _GEN_46718;
  wire        _GEN_47103 = _GEN_2085 ? ~_GEN_2109 & _GEN_46719 : ~_GEN_2076 & _GEN_46719;
  wire        _GEN_47104 = _GEN_2085 ? ~_GEN_2110 & _GEN_46720 : ~_GEN_2077 & _GEN_46720;
  wire        _GEN_47105 = _GEN_2085 ? ~_GEN_2111 & _GEN_46721 : ~_GEN_2078 & _GEN_46721;
  wire        _GEN_47106 = _GEN_2085 ? ~_GEN_2112 & _GEN_46722 : ~_GEN_2079 & _GEN_46722;
  wire        _GEN_47107 = _GEN_2085 ? ~_GEN_2113 & _GEN_46723 : ~_GEN_2080 & _GEN_46723;
  wire        _GEN_47108 = _GEN_2085 ? ~_GEN_2114 & _GEN_46724 : ~_GEN_2081 & _GEN_46724;
  wire        _GEN_47109 = _GEN_2085 ? ~_GEN_2115 & _GEN_46725 : ~_GEN_2082 & _GEN_46725;
  wire        _GEN_47110 = _GEN_2085 ? ~_GEN_2116 & _GEN_46726 : ~_GEN_2083 & _GEN_46726;
  wire        _GEN_47111 = _GEN_2085 ? ~_GEN_2117 & _GEN_46727 : ~_GEN_2084 & _GEN_46727;
  wire        _GEN_47464 = _GEN_2151 ? ~_GEN_2152 & _GEN_47080 : ~_GEN_2119 & _GEN_47080;
  wire        _GEN_47465 = _GEN_2151 ? ~_GEN_2153 & _GEN_47081 : ~_GEN_2120 & _GEN_47081;
  wire        _GEN_47466 = _GEN_2151 ? ~_GEN_2154 & _GEN_47082 : ~_GEN_2121 & _GEN_47082;
  wire        _GEN_47467 = _GEN_2151 ? ~_GEN_2155 & _GEN_47083 : ~_GEN_2122 & _GEN_47083;
  wire        _GEN_47468 = _GEN_2151 ? ~_GEN_2156 & _GEN_47084 : ~_GEN_2123 & _GEN_47084;
  wire        _GEN_47469 = _GEN_2151 ? ~_GEN_2157 & _GEN_47085 : ~_GEN_2124 & _GEN_47085;
  wire        _GEN_47470 = _GEN_2151 ? ~_GEN_2158 & _GEN_47086 : ~_GEN_2125 & _GEN_47086;
  wire        _GEN_47471 = _GEN_2151 ? ~_GEN_2159 & _GEN_47087 : ~_GEN_2126 & _GEN_47087;
  wire        _GEN_47472 = _GEN_2151 ? ~_GEN_2160 & _GEN_47088 : ~_GEN_2127 & _GEN_47088;
  wire        _GEN_47473 = _GEN_2151 ? ~_GEN_2161 & _GEN_47089 : ~_GEN_2128 & _GEN_47089;
  wire        _GEN_47474 = _GEN_2151 ? ~_GEN_2162 & _GEN_47090 : ~_GEN_2129 & _GEN_47090;
  wire        _GEN_47475 = _GEN_2151 ? ~_GEN_2163 & _GEN_47091 : ~_GEN_2130 & _GEN_47091;
  wire        _GEN_47476 = _GEN_2151 ? ~_GEN_2164 & _GEN_47092 : ~_GEN_2131 & _GEN_47092;
  wire        _GEN_47477 = _GEN_2151 ? ~_GEN_2165 & _GEN_47093 : ~_GEN_2132 & _GEN_47093;
  wire        _GEN_47478 = _GEN_2151 ? ~_GEN_2166 & _GEN_47094 : ~_GEN_2133 & _GEN_47094;
  wire        _GEN_47479 = _GEN_2151 ? ~_GEN_2167 & _GEN_47095 : ~_GEN_2134 & _GEN_47095;
  wire        _GEN_47480 = _GEN_2151 ? ~_GEN_2168 & _GEN_47096 : ~_GEN_2135 & _GEN_47096;
  wire        _GEN_47481 = _GEN_2151 ? ~_GEN_2169 & _GEN_47097 : ~_GEN_2136 & _GEN_47097;
  wire        _GEN_47482 = _GEN_2151 ? ~_GEN_2170 & _GEN_47098 : ~_GEN_2137 & _GEN_47098;
  wire        _GEN_47483 = _GEN_2151 ? ~_GEN_2171 & _GEN_47099 : ~_GEN_2138 & _GEN_47099;
  wire        _GEN_47484 = _GEN_2151 ? ~_GEN_2172 & _GEN_47100 : ~_GEN_2139 & _GEN_47100;
  wire        _GEN_47485 = _GEN_2151 ? ~_GEN_2173 & _GEN_47101 : ~_GEN_2140 & _GEN_47101;
  wire        _GEN_47486 = _GEN_2151 ? ~_GEN_2174 & _GEN_47102 : ~_GEN_2141 & _GEN_47102;
  wire        _GEN_47487 = _GEN_2151 ? ~_GEN_2175 & _GEN_47103 : ~_GEN_2142 & _GEN_47103;
  wire        _GEN_47488 = _GEN_2151 ? ~_GEN_2176 & _GEN_47104 : ~_GEN_2143 & _GEN_47104;
  wire        _GEN_47489 = _GEN_2151 ? ~_GEN_2177 & _GEN_47105 : ~_GEN_2144 & _GEN_47105;
  wire        _GEN_47490 = _GEN_2151 ? ~_GEN_2178 & _GEN_47106 : ~_GEN_2145 & _GEN_47106;
  wire        _GEN_47491 = _GEN_2151 ? ~_GEN_2179 & _GEN_47107 : ~_GEN_2146 & _GEN_47107;
  wire        _GEN_47492 = _GEN_2151 ? ~_GEN_2180 & _GEN_47108 : ~_GEN_2147 & _GEN_47108;
  wire        _GEN_47493 = _GEN_2151 ? ~_GEN_2181 & _GEN_47109 : ~_GEN_2148 & _GEN_47109;
  wire        _GEN_47494 = _GEN_2151 ? ~_GEN_2182 & _GEN_47110 : ~_GEN_2149 & _GEN_47110;
  wire        _GEN_47495 = _GEN_2151 ? ~_GEN_2183 & _GEN_47111 : ~_GEN_2150 & _GEN_47111;
  wire        _GEN_2676 = io_fflags_0_valid & (&(io_fflags_0_bits_uop_rob_idx[1:0]));
  wire        _GEN_2677 = io_fflags_2_valid & (&(io_fflags_2_bits_uop_rob_idx[1:0]));
  wire        _GEN_2678 = io_fflags_3_valid & (&(io_fflags_3_bits_uop_rob_idx[1:0]));
  wire        _GEN_2679 = rbk_row_3 & _GEN_2477;
  wire        _GEN_2680 = rbk_row_3 & _GEN_2447;
  wire        _GEN_2681 = rbk_row_3 & _GEN_2448;
  wire        _GEN_2682 = rbk_row_3 & _GEN_2449;
  wire        _GEN_2683 = rbk_row_3 & _GEN_2450;
  wire        _GEN_2684 = rbk_row_3 & _GEN_2451;
  wire        _GEN_2685 = rbk_row_3 & _GEN_2452;
  wire        _GEN_2686 = rbk_row_3 & _GEN_2453;
  wire        _GEN_2687 = rbk_row_3 & _GEN_2454;
  wire        _GEN_2688 = rbk_row_3 & _GEN_2455;
  wire        _GEN_2689 = rbk_row_3 & _GEN_2456;
  wire        _GEN_2690 = rbk_row_3 & _GEN_2457;
  wire        _GEN_2691 = rbk_row_3 & _GEN_2458;
  wire        _GEN_2692 = rbk_row_3 & _GEN_2459;
  wire        _GEN_2693 = rbk_row_3 & _GEN_2460;
  wire        _GEN_2694 = rbk_row_3 & _GEN_2461;
  wire        _GEN_2695 = rbk_row_3 & _GEN_2462;
  wire        _GEN_2696 = rbk_row_3 & _GEN_2463;
  wire        _GEN_2697 = rbk_row_3 & _GEN_2464;
  wire        _GEN_2698 = rbk_row_3 & _GEN_2465;
  wire        _GEN_2699 = rbk_row_3 & _GEN_2466;
  wire        _GEN_2700 = rbk_row_3 & _GEN_2467;
  wire        _GEN_2701 = rbk_row_3 & _GEN_2468;
  wire        _GEN_2702 = rbk_row_3 & _GEN_2469;
  wire        _GEN_2703 = rbk_row_3 & _GEN_2470;
  wire        _GEN_2704 = rbk_row_3 & _GEN_2471;
  wire        _GEN_2705 = rbk_row_3 & _GEN_2472;
  wire        _GEN_2706 = rbk_row_3 & _GEN_2473;
  wire        _GEN_2707 = rbk_row_3 & _GEN_2474;
  wire        _GEN_2708 = rbk_row_3 & _GEN_2475;
  wire        _GEN_2709 = rbk_row_3 & _GEN_2476;
  wire        _GEN_2710 = rbk_row_3 & (&com_idx);
  wire [19:0] _GEN_2711 = io_brupdate_b1_mispredict_mask & rob_uop_3_0_br_mask;
  wire [19:0] _GEN_2712 = io_brupdate_b1_mispredict_mask & rob_uop_3_1_br_mask;
  wire [19:0] _GEN_2713 = io_brupdate_b1_mispredict_mask & rob_uop_3_2_br_mask;
  wire [19:0] _GEN_2714 = io_brupdate_b1_mispredict_mask & rob_uop_3_3_br_mask;
  wire [19:0] _GEN_2715 = io_brupdate_b1_mispredict_mask & rob_uop_3_4_br_mask;
  wire [19:0] _GEN_2716 = io_brupdate_b1_mispredict_mask & rob_uop_3_5_br_mask;
  wire [19:0] _GEN_2717 = io_brupdate_b1_mispredict_mask & rob_uop_3_6_br_mask;
  wire [19:0] _GEN_2718 = io_brupdate_b1_mispredict_mask & rob_uop_3_7_br_mask;
  wire [19:0] _GEN_2719 = io_brupdate_b1_mispredict_mask & rob_uop_3_8_br_mask;
  wire [19:0] _GEN_2720 = io_brupdate_b1_mispredict_mask & rob_uop_3_9_br_mask;
  wire [19:0] _GEN_2721 = io_brupdate_b1_mispredict_mask & rob_uop_3_10_br_mask;
  wire [19:0] _GEN_2722 = io_brupdate_b1_mispredict_mask & rob_uop_3_11_br_mask;
  wire [19:0] _GEN_2723 = io_brupdate_b1_mispredict_mask & rob_uop_3_12_br_mask;
  wire [19:0] _GEN_2724 = io_brupdate_b1_mispredict_mask & rob_uop_3_13_br_mask;
  wire [19:0] _GEN_2725 = io_brupdate_b1_mispredict_mask & rob_uop_3_14_br_mask;
  wire [19:0] _GEN_2726 = io_brupdate_b1_mispredict_mask & rob_uop_3_15_br_mask;
  wire [19:0] _GEN_2727 = io_brupdate_b1_mispredict_mask & rob_uop_3_16_br_mask;
  wire [19:0] _GEN_2728 = io_brupdate_b1_mispredict_mask & rob_uop_3_17_br_mask;
  wire [19:0] _GEN_2729 = io_brupdate_b1_mispredict_mask & rob_uop_3_18_br_mask;
  wire [19:0] _GEN_2730 = io_brupdate_b1_mispredict_mask & rob_uop_3_19_br_mask;
  wire [19:0] _GEN_2731 = io_brupdate_b1_mispredict_mask & rob_uop_3_20_br_mask;
  wire [19:0] _GEN_2732 = io_brupdate_b1_mispredict_mask & rob_uop_3_21_br_mask;
  wire [19:0] _GEN_2733 = io_brupdate_b1_mispredict_mask & rob_uop_3_22_br_mask;
  wire [19:0] _GEN_2734 = io_brupdate_b1_mispredict_mask & rob_uop_3_23_br_mask;
  wire [19:0] _GEN_2735 = io_brupdate_b1_mispredict_mask & rob_uop_3_24_br_mask;
  wire [19:0] _GEN_2736 = io_brupdate_b1_mispredict_mask & rob_uop_3_25_br_mask;
  wire [19:0] _GEN_2737 = io_brupdate_b1_mispredict_mask & rob_uop_3_26_br_mask;
  wire [19:0] _GEN_2738 = io_brupdate_b1_mispredict_mask & rob_uop_3_27_br_mask;
  wire [19:0] _GEN_2739 = io_brupdate_b1_mispredict_mask & rob_uop_3_28_br_mask;
  wire [19:0] _GEN_2740 = io_brupdate_b1_mispredict_mask & rob_uop_3_29_br_mask;
  wire [19:0] _GEN_2741 = io_brupdate_b1_mispredict_mask & rob_uop_3_30_br_mask;
  wire [19:0] _GEN_2742 = io_brupdate_b1_mispredict_mask & rob_uop_3_31_br_mask;
  wire        _GEN_2743 = ~(_io_flush_valid_output | exception_thrown) & rob_state != 2'h2;
  wire        _GEN_2744 = ~r_xcpt_val | io_lxcpt_bits_uop_rob_idx < r_xcpt_uop_rob_idx ^ io_lxcpt_bits_uop_rob_idx < rob_head_idx ^ r_xcpt_uop_rob_idx < rob_head_idx;
  wire        _GEN_2745 = ~r_xcpt_val & (enq_xcpts_0 | enq_xcpts_1 | enq_xcpts_2 | io_enq_valids_3 & io_enq_uops_3_exception);
  wire [19:0] next_xcpt_uop_br_mask = _GEN_2743 ? (io_lxcpt_valid ? (_GEN_2744 ? io_lxcpt_bits_uop_br_mask : r_xcpt_uop_br_mask) : _GEN_2745 ? casez_tmp_91 : r_xcpt_uop_br_mask) : r_xcpt_uop_br_mask;
  wire        _GEN_2746 = (|_GEN_2510) | _GEN_2478;
  wire        _GEN_2747 = (|_GEN_2511) | _GEN_2479;
  wire        _GEN_2748 = (|_GEN_2512) | _GEN_2480;
  wire        _GEN_2749 = (|_GEN_2513) | _GEN_2481;
  wire        _GEN_2750 = (|_GEN_2514) | _GEN_2482;
  wire        _GEN_2751 = (|_GEN_2515) | _GEN_2483;
  wire        _GEN_2752 = (|_GEN_2516) | _GEN_2484;
  wire        _GEN_2753 = (|_GEN_2517) | _GEN_2485;
  wire        _GEN_2754 = (|_GEN_2518) | _GEN_2486;
  wire        _GEN_2755 = (|_GEN_2519) | _GEN_2487;
  wire        _GEN_2756 = (|_GEN_2520) | _GEN_2488;
  wire        _GEN_2757 = (|_GEN_2521) | _GEN_2489;
  wire        _GEN_2758 = (|_GEN_2522) | _GEN_2490;
  wire        _GEN_2759 = (|_GEN_2523) | _GEN_2491;
  wire        _GEN_2760 = (|_GEN_2524) | _GEN_2492;
  wire        _GEN_2761 = (|_GEN_2525) | _GEN_2493;
  wire        _GEN_2762 = (|_GEN_2526) | _GEN_2494;
  wire        _GEN_2763 = (|_GEN_2527) | _GEN_2495;
  wire        _GEN_2764 = (|_GEN_2528) | _GEN_2496;
  wire        _GEN_2765 = (|_GEN_2529) | _GEN_2497;
  wire        _GEN_2766 = (|_GEN_2530) | _GEN_2498;
  wire        _GEN_2767 = (|_GEN_2531) | _GEN_2499;
  wire        _GEN_2768 = (|_GEN_2532) | _GEN_2500;
  wire        _GEN_2769 = (|_GEN_2533) | _GEN_2501;
  wire        _GEN_2770 = (|_GEN_2534) | _GEN_2502;
  wire        _GEN_2771 = (|_GEN_2535) | _GEN_2503;
  wire        _GEN_2772 = (|_GEN_2536) | _GEN_2504;
  wire        _GEN_2773 = (|_GEN_2537) | _GEN_2505;
  wire        _GEN_2774 = (|_GEN_2538) | _GEN_2506;
  wire        _GEN_2775 = (|_GEN_2539) | _GEN_2507;
  wire        _GEN_2776 = (|_GEN_2540) | _GEN_2508;
  wire        _GEN_2777 = (|_GEN_2541) | _GEN_2509;
  wire        _GEN_2778 = (|_GEN_2577) | _GEN_2545;
  wire        _GEN_2779 = (|_GEN_2578) | _GEN_2546;
  wire        _GEN_2780 = (|_GEN_2579) | _GEN_2547;
  wire        _GEN_2781 = (|_GEN_2580) | _GEN_2548;
  wire        _GEN_2782 = (|_GEN_2581) | _GEN_2549;
  wire        _GEN_2783 = (|_GEN_2582) | _GEN_2550;
  wire        _GEN_2784 = (|_GEN_2583) | _GEN_2551;
  wire        _GEN_2785 = (|_GEN_2584) | _GEN_2552;
  wire        _GEN_2786 = (|_GEN_2585) | _GEN_2553;
  wire        _GEN_2787 = (|_GEN_2586) | _GEN_2554;
  wire        _GEN_2788 = (|_GEN_2587) | _GEN_2555;
  wire        _GEN_2789 = (|_GEN_2588) | _GEN_2556;
  wire        _GEN_2790 = (|_GEN_2589) | _GEN_2557;
  wire        _GEN_2791 = (|_GEN_2590) | _GEN_2558;
  wire        _GEN_2792 = (|_GEN_2591) | _GEN_2559;
  wire        _GEN_2793 = (|_GEN_2592) | _GEN_2560;
  wire        _GEN_2794 = (|_GEN_2593) | _GEN_2561;
  wire        _GEN_2795 = (|_GEN_2594) | _GEN_2562;
  wire        _GEN_2796 = (|_GEN_2595) | _GEN_2563;
  wire        _GEN_2797 = (|_GEN_2596) | _GEN_2564;
  wire        _GEN_2798 = (|_GEN_2597) | _GEN_2565;
  wire        _GEN_2799 = (|_GEN_2598) | _GEN_2566;
  wire        _GEN_2800 = (|_GEN_2599) | _GEN_2567;
  wire        _GEN_2801 = (|_GEN_2600) | _GEN_2568;
  wire        _GEN_2802 = (|_GEN_2601) | _GEN_2569;
  wire        _GEN_2803 = (|_GEN_2602) | _GEN_2570;
  wire        _GEN_2804 = (|_GEN_2603) | _GEN_2571;
  wire        _GEN_2805 = (|_GEN_2604) | _GEN_2572;
  wire        _GEN_2806 = (|_GEN_2605) | _GEN_2573;
  wire        _GEN_2807 = (|_GEN_2606) | _GEN_2574;
  wire        _GEN_2808 = (|_GEN_2607) | _GEN_2575;
  wire        _GEN_2809 = (|_GEN_2608) | _GEN_2576;
  wire        _GEN_2810 = (|_GEN_2644) | _GEN_2612;
  wire        _GEN_2811 = (|_GEN_2645) | _GEN_2613;
  wire        _GEN_2812 = (|_GEN_2646) | _GEN_2614;
  wire        _GEN_2813 = (|_GEN_2647) | _GEN_2615;
  wire        _GEN_2814 = (|_GEN_2648) | _GEN_2616;
  wire        _GEN_2815 = (|_GEN_2649) | _GEN_2617;
  wire        _GEN_2816 = (|_GEN_2650) | _GEN_2618;
  wire        _GEN_2817 = (|_GEN_2651) | _GEN_2619;
  wire        _GEN_2818 = (|_GEN_2652) | _GEN_2620;
  wire        _GEN_2819 = (|_GEN_2653) | _GEN_2621;
  wire        _GEN_2820 = (|_GEN_2654) | _GEN_2622;
  wire        _GEN_2821 = (|_GEN_2655) | _GEN_2623;
  wire        _GEN_2822 = (|_GEN_2656) | _GEN_2624;
  wire        _GEN_2823 = (|_GEN_2657) | _GEN_2625;
  wire        _GEN_2824 = (|_GEN_2658) | _GEN_2626;
  wire        _GEN_2825 = (|_GEN_2659) | _GEN_2627;
  wire        _GEN_2826 = (|_GEN_2660) | _GEN_2628;
  wire        _GEN_2827 = (|_GEN_2661) | _GEN_2629;
  wire        _GEN_2892 = (|_GEN_2662) | _GEN_2630;
  wire        _GEN_2893 = (|_GEN_2663) | _GEN_2631;
  wire        _GEN_2894 = (|_GEN_2664) | _GEN_2632;
  wire        _GEN_2895 = (|_GEN_2665) | _GEN_2633;
  wire        _GEN_2896 = (|_GEN_2666) | _GEN_2634;
  wire        _GEN_2897 = (|_GEN_2667) | _GEN_2635;
  wire        _GEN_2898 = (|_GEN_2668) | _GEN_2636;
  wire        _GEN_2899 = (|_GEN_2669) | _GEN_2637;
  wire        _GEN_2900 = (|_GEN_2670) | _GEN_2638;
  wire        _GEN_2901 = (|_GEN_2671) | _GEN_2639;
  wire        _GEN_2902 = (|_GEN_2672) | _GEN_2640;
  wire        _GEN_2903 = (|_GEN_2673) | _GEN_2641;
  wire        _GEN_2904 = (|_GEN_2674) | _GEN_2642;
  wire        _GEN_2905 = (|_GEN_2675) | _GEN_2643;
  wire        _GEN_2906 = (|_GEN_2711) | _GEN_2679;
  wire        _GEN_2907 = (|_GEN_2712) | _GEN_2680;
  wire        _GEN_2908 = (|_GEN_2713) | _GEN_2681;
  wire        _GEN_2909 = (|_GEN_2714) | _GEN_2682;
  wire        _GEN_2910 = (|_GEN_2715) | _GEN_2683;
  wire        _GEN_2911 = (|_GEN_2716) | _GEN_2684;
  wire        _GEN_2912 = (|_GEN_2717) | _GEN_2685;
  wire        _GEN_2913 = (|_GEN_2718) | _GEN_2686;
  wire        _GEN_2914 = (|_GEN_2719) | _GEN_2687;
  wire        _GEN_2915 = (|_GEN_2720) | _GEN_2688;
  wire        _GEN_2916 = (|_GEN_2721) | _GEN_2689;
  wire        _GEN_2917 = (|_GEN_2722) | _GEN_2690;
  wire        _GEN_2918 = (|_GEN_2723) | _GEN_2691;
  wire        _GEN_2919 = (|_GEN_2724) | _GEN_2692;
  wire        _GEN_2920 = (|_GEN_2725) | _GEN_2693;
  wire        _GEN_2921 = (|_GEN_2726) | _GEN_2694;
  wire        _GEN_2922 = (|_GEN_2727) | _GEN_2695;
  wire        _GEN_2923 = (|_GEN_2728) | _GEN_2696;
  wire        _GEN_2924 = (|_GEN_2729) | _GEN_2697;
  wire        _GEN_2925 = (|_GEN_2730) | _GEN_2698;
  wire        _GEN_2926 = (|_GEN_2731) | _GEN_2699;
  wire        _GEN_2927 = (|_GEN_2732) | _GEN_2700;
  wire        _GEN_2928 = (|_GEN_2733) | _GEN_2701;
  wire        _GEN_2929 = (|_GEN_2734) | _GEN_2702;
  wire        _GEN_2930 = (|_GEN_2735) | _GEN_2703;
  wire        _GEN_2931 = (|_GEN_2736) | _GEN_2704;
  wire        _GEN_2932 = (|_GEN_2737) | _GEN_2705;
  wire        _GEN_2933 = (|_GEN_2738) | _GEN_2706;
  wire        _GEN_2934 = (|_GEN_2739) | _GEN_2707;
  wire        _GEN_2935 = (|_GEN_2740) | _GEN_2708;
  wire        _GEN_2936 = (|_GEN_2741) | _GEN_2709;
  wire        _GEN_2937 = (|_GEN_2742) | _GEN_2710;
  always @(posedge clock) begin
    if (reset) begin
      rob_state <= 2'h0;
      rob_head <= 5'h0;
      rob_head_lsb <= 2'h0;
      rob_tail <= 5'h0;
      rob_tail_lsb <= 2'h0;
      maybe_full <= 1'h0;
      r_xcpt_val <= 1'h0;
      rob_val__31 <= 1'h0;
      rob_val__30 <= 1'h0;
      rob_val__29 <= 1'h0;
      rob_val__28 <= 1'h0;
      rob_val__27 <= 1'h0;
      rob_val__26 <= 1'h0;
      rob_val__25 <= 1'h0;
      rob_val__24 <= 1'h0;
      rob_val__23 <= 1'h0;
      rob_val__22 <= 1'h0;
      rob_val__21 <= 1'h0;
      rob_val__20 <= 1'h0;
      rob_val__19 <= 1'h0;
      rob_val__18 <= 1'h0;
      rob_val__17 <= 1'h0;
      rob_val__16 <= 1'h0;
      rob_val__15 <= 1'h0;
      rob_val__14 <= 1'h0;
      rob_val__13 <= 1'h0;
      rob_val__12 <= 1'h0;
      rob_val__11 <= 1'h0;
      rob_val__10 <= 1'h0;
      rob_val__9 <= 1'h0;
      rob_val__8 <= 1'h0;
      rob_val__7 <= 1'h0;
      rob_val__6 <= 1'h0;
      rob_val__5 <= 1'h0;
      rob_val__4 <= 1'h0;
      rob_val__3 <= 1'h0;
      rob_val__2 <= 1'h0;
      rob_val__1 <= 1'h0;
      rob_val__0 <= 1'h0;
      rob_val_1_31 <= 1'h0;
      rob_val_1_30 <= 1'h0;
      rob_val_1_29 <= 1'h0;
      rob_val_1_28 <= 1'h0;
      rob_val_1_27 <= 1'h0;
      rob_val_1_26 <= 1'h0;
      rob_val_1_25 <= 1'h0;
      rob_val_1_24 <= 1'h0;
      rob_val_1_23 <= 1'h0;
      rob_val_1_22 <= 1'h0;
      rob_val_1_21 <= 1'h0;
      rob_val_1_20 <= 1'h0;
      rob_val_1_19 <= 1'h0;
      rob_val_1_18 <= 1'h0;
      rob_val_1_17 <= 1'h0;
      rob_val_1_16 <= 1'h0;
      rob_val_1_15 <= 1'h0;
      rob_val_1_14 <= 1'h0;
      rob_val_1_13 <= 1'h0;
      rob_val_1_12 <= 1'h0;
      rob_val_1_11 <= 1'h0;
      rob_val_1_10 <= 1'h0;
      rob_val_1_9 <= 1'h0;
      rob_val_1_8 <= 1'h0;
      rob_val_1_7 <= 1'h0;
      rob_val_1_6 <= 1'h0;
      rob_val_1_5 <= 1'h0;
      rob_val_1_4 <= 1'h0;
      rob_val_1_3 <= 1'h0;
      rob_val_1_2 <= 1'h0;
      rob_val_1_1 <= 1'h0;
      rob_val_1_0 <= 1'h0;
      rob_val_2_31 <= 1'h0;
      rob_val_2_30 <= 1'h0;
      rob_val_2_29 <= 1'h0;
      rob_val_2_28 <= 1'h0;
      rob_val_2_27 <= 1'h0;
      rob_val_2_26 <= 1'h0;
      rob_val_2_25 <= 1'h0;
      rob_val_2_24 <= 1'h0;
      rob_val_2_23 <= 1'h0;
      rob_val_2_22 <= 1'h0;
      rob_val_2_21 <= 1'h0;
      rob_val_2_20 <= 1'h0;
      rob_val_2_19 <= 1'h0;
      rob_val_2_18 <= 1'h0;
      rob_val_2_17 <= 1'h0;
      rob_val_2_16 <= 1'h0;
      rob_val_2_15 <= 1'h0;
      rob_val_2_14 <= 1'h0;
      rob_val_2_13 <= 1'h0;
      rob_val_2_12 <= 1'h0;
      rob_val_2_11 <= 1'h0;
      rob_val_2_10 <= 1'h0;
      rob_val_2_9 <= 1'h0;
      rob_val_2_8 <= 1'h0;
      rob_val_2_7 <= 1'h0;
      rob_val_2_6 <= 1'h0;
      rob_val_2_5 <= 1'h0;
      rob_val_2_4 <= 1'h0;
      rob_val_2_3 <= 1'h0;
      rob_val_2_2 <= 1'h0;
      rob_val_2_1 <= 1'h0;
      rob_val_2_0 <= 1'h0;
      rob_val_3_31 <= 1'h0;
      rob_val_3_30 <= 1'h0;
      rob_val_3_29 <= 1'h0;
      rob_val_3_28 <= 1'h0;
      rob_val_3_27 <= 1'h0;
      rob_val_3_26 <= 1'h0;
      rob_val_3_25 <= 1'h0;
      rob_val_3_24 <= 1'h0;
      rob_val_3_23 <= 1'h0;
      rob_val_3_22 <= 1'h0;
      rob_val_3_21 <= 1'h0;
      rob_val_3_20 <= 1'h0;
      rob_val_3_19 <= 1'h0;
      rob_val_3_18 <= 1'h0;
      rob_val_3_17 <= 1'h0;
      rob_val_3_16 <= 1'h0;
      rob_val_3_15 <= 1'h0;
      rob_val_3_14 <= 1'h0;
      rob_val_3_13 <= 1'h0;
      rob_val_3_12 <= 1'h0;
      rob_val_3_11 <= 1'h0;
      rob_val_3_10 <= 1'h0;
      rob_val_3_9 <= 1'h0;
      rob_val_3_8 <= 1'h0;
      rob_val_3_7 <= 1'h0;
      rob_val_3_6 <= 1'h0;
      rob_val_3_5 <= 1'h0;
      rob_val_3_4 <= 1'h0;
      rob_val_3_3 <= 1'h0;
      rob_val_3_2 <= 1'h0;
      rob_val_3_1 <= 1'h0;
      rob_val_3_0 <= 1'h0;
      r_partial_row <= 1'h0;
    end
    else begin
      rob_state <= casez_tmp_95;
      if (finished_committing_row) begin
        rob_head <= rob_head + 5'h1;
        rob_head_lsb <= 2'h0;
      end
      else
        rob_head_lsb <= {|(_rob_head_lsb_T_8[2:1]), _rob_head_lsb_T_8[2] | _rob_head_lsb_T_8[0]};
      if (_GEN_2285) begin
        rob_tail <= rob_tail - 5'h1;
        rob_tail_lsb <= 2'h3;
      end
      else if (_GEN_2319)
        rob_tail_lsb <= rob_head_lsb;
      else begin
        if (io_brupdate_b2_mispredict)
          rob_tail <= io_brupdate_b2_uop_rob_idx[6:2] + 5'h1;
        else if (_GEN_54123)
          rob_tail <= rob_tail + 5'h1;
        if (io_brupdate_b2_mispredict | _GEN_54123)
          rob_tail_lsb <= 2'h0;
        else if ((|_GEN_2284) & io_enq_partial_stall) begin
          if (_rob_tail_lsb_T_8[0])
            rob_tail_lsb <= 2'h0;
          else if (_rob_tail_lsb_T_8[1])
            rob_tail_lsb <= 2'h1;
          else
            rob_tail_lsb <= {1'h1, ~(_rob_tail_lsb_T_8[2])};
        end
      end
      maybe_full <= ~rob_deq & (~(_GEN_2285 | _GEN_2319 | io_brupdate_b2_mispredict) & _GEN_54123 | maybe_full) | (|io_brupdate_b1_mispredict_mask);
      r_xcpt_val <= ~(_io_flush_valid_output | (|(io_brupdate_b1_mispredict_mask & next_xcpt_uop_br_mask))) & (_GEN_2743 ? (io_lxcpt_valid ? _GEN_2744 | r_xcpt_val : _GEN_2745 | r_xcpt_val) : r_xcpt_val);
      if (_io_commit_valids_0_output) begin
        rob_val__31 <= ~((&rob_head) | _GEN_2777) & _GEN_2859;
        rob_val__30 <= ~(_GEN_2317 | _GEN_2776) & _GEN_2858;
        rob_val__29 <= ~(_GEN_2316 | _GEN_2775) & _GEN_2857;
        rob_val__28 <= ~(_GEN_2315 | _GEN_2774) & _GEN_2856;
        rob_val__27 <= ~(_GEN_2314 | _GEN_2773) & _GEN_2855;
        rob_val__26 <= ~(_GEN_2313 | _GEN_2772) & _GEN_2854;
        rob_val__25 <= ~(_GEN_2312 | _GEN_2771) & _GEN_2853;
        rob_val__24 <= ~(_GEN_2311 | _GEN_2770) & _GEN_2852;
        rob_val__23 <= ~(_GEN_2310 | _GEN_2769) & _GEN_2851;
        rob_val__22 <= ~(_GEN_2309 | _GEN_2768) & _GEN_2850;
        rob_val__21 <= ~(_GEN_2308 | _GEN_2767) & _GEN_2849;
        rob_val__20 <= ~(_GEN_2307 | _GEN_2766) & _GEN_2848;
        rob_val__19 <= ~(_GEN_2306 | _GEN_2765) & _GEN_2847;
        rob_val__18 <= ~(_GEN_2305 | _GEN_2764) & _GEN_2846;
        rob_val__17 <= ~(_GEN_2304 | _GEN_2763) & _GEN_2845;
        rob_val__16 <= ~(_GEN_2303 | _GEN_2762) & _GEN_2844;
        rob_val__15 <= ~(_GEN_2302 | _GEN_2761) & _GEN_2843;
        rob_val__14 <= ~(_GEN_2301 | _GEN_2760) & _GEN_2842;
        rob_val__13 <= ~(_GEN_2300 | _GEN_2759) & _GEN_2841;
        rob_val__12 <= ~(_GEN_2299 | _GEN_2758) & _GEN_2840;
        rob_val__11 <= ~(_GEN_2298 | _GEN_2757) & _GEN_2839;
        rob_val__10 <= ~(_GEN_2297 | _GEN_2756) & _GEN_2838;
        rob_val__9 <= ~(_GEN_2296 | _GEN_2755) & _GEN_2837;
        rob_val__8 <= ~(_GEN_2295 | _GEN_2754) & _GEN_2836;
        rob_val__7 <= ~(_GEN_2294 | _GEN_2753) & _GEN_2835;
        rob_val__6 <= ~(_GEN_2293 | _GEN_2752) & _GEN_2834;
        rob_val__5 <= ~(_GEN_2292 | _GEN_2751) & _GEN_2833;
        rob_val__4 <= ~(_GEN_2291 | _GEN_2750) & _GEN_2832;
        rob_val__3 <= ~(_GEN_2290 | _GEN_2749) & _GEN_2831;
        rob_val__2 <= ~(_GEN_2289 | _GEN_2748) & _GEN_2830;
        rob_val__1 <= ~(_GEN_2288 | _GEN_2747) & _GEN_2829;
        rob_val__0 <= ~(_GEN_2318 | _GEN_2746) & _GEN_2828;
      end
      else begin
        rob_val__31 <= ~_GEN_2777 & _GEN_2859;
        rob_val__30 <= ~_GEN_2776 & _GEN_2858;
        rob_val__29 <= ~_GEN_2775 & _GEN_2857;
        rob_val__28 <= ~_GEN_2774 & _GEN_2856;
        rob_val__27 <= ~_GEN_2773 & _GEN_2855;
        rob_val__26 <= ~_GEN_2772 & _GEN_2854;
        rob_val__25 <= ~_GEN_2771 & _GEN_2853;
        rob_val__24 <= ~_GEN_2770 & _GEN_2852;
        rob_val__23 <= ~_GEN_2769 & _GEN_2851;
        rob_val__22 <= ~_GEN_2768 & _GEN_2850;
        rob_val__21 <= ~_GEN_2767 & _GEN_2849;
        rob_val__20 <= ~_GEN_2766 & _GEN_2848;
        rob_val__19 <= ~_GEN_2765 & _GEN_2847;
        rob_val__18 <= ~_GEN_2764 & _GEN_2846;
        rob_val__17 <= ~_GEN_2763 & _GEN_2845;
        rob_val__16 <= ~_GEN_2762 & _GEN_2844;
        rob_val__15 <= ~_GEN_2761 & _GEN_2843;
        rob_val__14 <= ~_GEN_2760 & _GEN_2842;
        rob_val__13 <= ~_GEN_2759 & _GEN_2841;
        rob_val__12 <= ~_GEN_2758 & _GEN_2840;
        rob_val__11 <= ~_GEN_2757 & _GEN_2839;
        rob_val__10 <= ~_GEN_2756 & _GEN_2838;
        rob_val__9 <= ~_GEN_2755 & _GEN_2837;
        rob_val__8 <= ~_GEN_2754 & _GEN_2836;
        rob_val__7 <= ~_GEN_2753 & _GEN_2835;
        rob_val__6 <= ~_GEN_2752 & _GEN_2834;
        rob_val__5 <= ~_GEN_2751 & _GEN_2833;
        rob_val__4 <= ~_GEN_2750 & _GEN_2832;
        rob_val__3 <= ~_GEN_2749 & _GEN_2831;
        rob_val__2 <= ~_GEN_2748 & _GEN_2830;
        rob_val__1 <= ~_GEN_2747 & _GEN_2829;
        rob_val__0 <= ~_GEN_2746 & _GEN_2828;
      end
      if (_io_commit_valids_1_output) begin
        rob_val_1_31 <= ~((&rob_head) | _GEN_2809) & _GEN_16223;
        rob_val_1_30 <= ~(_GEN_2317 | _GEN_2808) & _GEN_16222;
        rob_val_1_29 <= ~(_GEN_2316 | _GEN_2807) & _GEN_16221;
        rob_val_1_28 <= ~(_GEN_2315 | _GEN_2806) & _GEN_16220;
        rob_val_1_27 <= ~(_GEN_2314 | _GEN_2805) & _GEN_16219;
        rob_val_1_26 <= ~(_GEN_2313 | _GEN_2804) & _GEN_16218;
        rob_val_1_25 <= ~(_GEN_2312 | _GEN_2803) & _GEN_16217;
        rob_val_1_24 <= ~(_GEN_2311 | _GEN_2802) & _GEN_16216;
        rob_val_1_23 <= ~(_GEN_2310 | _GEN_2801) & _GEN_16215;
        rob_val_1_22 <= ~(_GEN_2309 | _GEN_2800) & _GEN_16214;
        rob_val_1_21 <= ~(_GEN_2308 | _GEN_2799) & _GEN_16213;
        rob_val_1_20 <= ~(_GEN_2307 | _GEN_2798) & _GEN_16212;
        rob_val_1_19 <= ~(_GEN_2306 | _GEN_2797) & _GEN_16211;
        rob_val_1_18 <= ~(_GEN_2305 | _GEN_2796) & _GEN_16210;
        rob_val_1_17 <= ~(_GEN_2304 | _GEN_2795) & _GEN_16209;
        rob_val_1_16 <= ~(_GEN_2303 | _GEN_2794) & _GEN_16208;
        rob_val_1_15 <= ~(_GEN_2302 | _GEN_2793) & _GEN_16207;
        rob_val_1_14 <= ~(_GEN_2301 | _GEN_2792) & _GEN_16206;
        rob_val_1_13 <= ~(_GEN_2300 | _GEN_2791) & _GEN_16205;
        rob_val_1_12 <= ~(_GEN_2299 | _GEN_2790) & _GEN_16204;
        rob_val_1_11 <= ~(_GEN_2298 | _GEN_2789) & _GEN_16203;
        rob_val_1_10 <= ~(_GEN_2297 | _GEN_2788) & _GEN_16202;
        rob_val_1_9 <= ~(_GEN_2296 | _GEN_2787) & _GEN_16201;
        rob_val_1_8 <= ~(_GEN_2295 | _GEN_2786) & _GEN_16200;
        rob_val_1_7 <= ~(_GEN_2294 | _GEN_2785) & _GEN_16199;
        rob_val_1_6 <= ~(_GEN_2293 | _GEN_2784) & _GEN_16198;
        rob_val_1_5 <= ~(_GEN_2292 | _GEN_2783) & _GEN_16197;
        rob_val_1_4 <= ~(_GEN_2291 | _GEN_2782) & _GEN_16196;
        rob_val_1_3 <= ~(_GEN_2290 | _GEN_2781) & _GEN_16195;
        rob_val_1_2 <= ~(_GEN_2289 | _GEN_2780) & _GEN_16194;
        rob_val_1_1 <= ~(_GEN_2288 | _GEN_2779) & _GEN_16193;
        rob_val_1_0 <= ~(_GEN_2318 | _GEN_2778) & _GEN_16192;
      end
      else begin
        rob_val_1_31 <= ~_GEN_2809 & _GEN_16223;
        rob_val_1_30 <= ~_GEN_2808 & _GEN_16222;
        rob_val_1_29 <= ~_GEN_2807 & _GEN_16221;
        rob_val_1_28 <= ~_GEN_2806 & _GEN_16220;
        rob_val_1_27 <= ~_GEN_2805 & _GEN_16219;
        rob_val_1_26 <= ~_GEN_2804 & _GEN_16218;
        rob_val_1_25 <= ~_GEN_2803 & _GEN_16217;
        rob_val_1_24 <= ~_GEN_2802 & _GEN_16216;
        rob_val_1_23 <= ~_GEN_2801 & _GEN_16215;
        rob_val_1_22 <= ~_GEN_2800 & _GEN_16214;
        rob_val_1_21 <= ~_GEN_2799 & _GEN_16213;
        rob_val_1_20 <= ~_GEN_2798 & _GEN_16212;
        rob_val_1_19 <= ~_GEN_2797 & _GEN_16211;
        rob_val_1_18 <= ~_GEN_2796 & _GEN_16210;
        rob_val_1_17 <= ~_GEN_2795 & _GEN_16209;
        rob_val_1_16 <= ~_GEN_2794 & _GEN_16208;
        rob_val_1_15 <= ~_GEN_2793 & _GEN_16207;
        rob_val_1_14 <= ~_GEN_2792 & _GEN_16206;
        rob_val_1_13 <= ~_GEN_2791 & _GEN_16205;
        rob_val_1_12 <= ~_GEN_2790 & _GEN_16204;
        rob_val_1_11 <= ~_GEN_2789 & _GEN_16203;
        rob_val_1_10 <= ~_GEN_2788 & _GEN_16202;
        rob_val_1_9 <= ~_GEN_2787 & _GEN_16201;
        rob_val_1_8 <= ~_GEN_2786 & _GEN_16200;
        rob_val_1_7 <= ~_GEN_2785 & _GEN_16199;
        rob_val_1_6 <= ~_GEN_2784 & _GEN_16198;
        rob_val_1_5 <= ~_GEN_2783 & _GEN_16197;
        rob_val_1_4 <= ~_GEN_2782 & _GEN_16196;
        rob_val_1_3 <= ~_GEN_2781 & _GEN_16195;
        rob_val_1_2 <= ~_GEN_2780 & _GEN_16194;
        rob_val_1_1 <= ~_GEN_2779 & _GEN_16193;
        rob_val_1_0 <= ~_GEN_2778 & _GEN_16192;
      end
      if (_io_commit_valids_2_output) begin
        rob_val_2_31 <= ~((&rob_head) | _GEN_2905) & _GEN_29587;
        rob_val_2_30 <= ~(_GEN_2317 | _GEN_2904) & _GEN_29586;
        rob_val_2_29 <= ~(_GEN_2316 | _GEN_2903) & _GEN_29585;
        rob_val_2_28 <= ~(_GEN_2315 | _GEN_2902) & _GEN_29584;
        rob_val_2_27 <= ~(_GEN_2314 | _GEN_2901) & _GEN_29583;
        rob_val_2_26 <= ~(_GEN_2313 | _GEN_2900) & _GEN_29582;
        rob_val_2_25 <= ~(_GEN_2312 | _GEN_2899) & _GEN_29581;
        rob_val_2_24 <= ~(_GEN_2311 | _GEN_2898) & _GEN_29580;
        rob_val_2_23 <= ~(_GEN_2310 | _GEN_2897) & _GEN_29579;
        rob_val_2_22 <= ~(_GEN_2309 | _GEN_2896) & _GEN_29578;
        rob_val_2_21 <= ~(_GEN_2308 | _GEN_2895) & _GEN_29577;
        rob_val_2_20 <= ~(_GEN_2307 | _GEN_2894) & _GEN_29576;
        rob_val_2_19 <= ~(_GEN_2306 | _GEN_2893) & _GEN_29575;
        rob_val_2_18 <= ~(_GEN_2305 | _GEN_2892) & _GEN_29574;
        rob_val_2_17 <= ~(_GEN_2304 | _GEN_2827) & _GEN_29573;
        rob_val_2_16 <= ~(_GEN_2303 | _GEN_2826) & _GEN_29572;
        rob_val_2_15 <= ~(_GEN_2302 | _GEN_2825) & _GEN_29571;
        rob_val_2_14 <= ~(_GEN_2301 | _GEN_2824) & _GEN_29570;
        rob_val_2_13 <= ~(_GEN_2300 | _GEN_2823) & _GEN_29569;
        rob_val_2_12 <= ~(_GEN_2299 | _GEN_2822) & _GEN_29568;
        rob_val_2_11 <= ~(_GEN_2298 | _GEN_2821) & _GEN_29567;
        rob_val_2_10 <= ~(_GEN_2297 | _GEN_2820) & _GEN_29566;
        rob_val_2_9 <= ~(_GEN_2296 | _GEN_2819) & _GEN_29565;
        rob_val_2_8 <= ~(_GEN_2295 | _GEN_2818) & _GEN_29564;
        rob_val_2_7 <= ~(_GEN_2294 | _GEN_2817) & _GEN_29563;
        rob_val_2_6 <= ~(_GEN_2293 | _GEN_2816) & _GEN_29562;
        rob_val_2_5 <= ~(_GEN_2292 | _GEN_2815) & _GEN_29561;
        rob_val_2_4 <= ~(_GEN_2291 | _GEN_2814) & _GEN_29560;
        rob_val_2_3 <= ~(_GEN_2290 | _GEN_2813) & _GEN_29559;
        rob_val_2_2 <= ~(_GEN_2289 | _GEN_2812) & _GEN_29558;
        rob_val_2_1 <= ~(_GEN_2288 | _GEN_2811) & _GEN_29557;
        rob_val_2_0 <= ~(_GEN_2318 | _GEN_2810) & _GEN_29556;
      end
      else begin
        rob_val_2_31 <= ~_GEN_2905 & _GEN_29587;
        rob_val_2_30 <= ~_GEN_2904 & _GEN_29586;
        rob_val_2_29 <= ~_GEN_2903 & _GEN_29585;
        rob_val_2_28 <= ~_GEN_2902 & _GEN_29584;
        rob_val_2_27 <= ~_GEN_2901 & _GEN_29583;
        rob_val_2_26 <= ~_GEN_2900 & _GEN_29582;
        rob_val_2_25 <= ~_GEN_2899 & _GEN_29581;
        rob_val_2_24 <= ~_GEN_2898 & _GEN_29580;
        rob_val_2_23 <= ~_GEN_2897 & _GEN_29579;
        rob_val_2_22 <= ~_GEN_2896 & _GEN_29578;
        rob_val_2_21 <= ~_GEN_2895 & _GEN_29577;
        rob_val_2_20 <= ~_GEN_2894 & _GEN_29576;
        rob_val_2_19 <= ~_GEN_2893 & _GEN_29575;
        rob_val_2_18 <= ~_GEN_2892 & _GEN_29574;
        rob_val_2_17 <= ~_GEN_2827 & _GEN_29573;
        rob_val_2_16 <= ~_GEN_2826 & _GEN_29572;
        rob_val_2_15 <= ~_GEN_2825 & _GEN_29571;
        rob_val_2_14 <= ~_GEN_2824 & _GEN_29570;
        rob_val_2_13 <= ~_GEN_2823 & _GEN_29569;
        rob_val_2_12 <= ~_GEN_2822 & _GEN_29568;
        rob_val_2_11 <= ~_GEN_2821 & _GEN_29567;
        rob_val_2_10 <= ~_GEN_2820 & _GEN_29566;
        rob_val_2_9 <= ~_GEN_2819 & _GEN_29565;
        rob_val_2_8 <= ~_GEN_2818 & _GEN_29564;
        rob_val_2_7 <= ~_GEN_2817 & _GEN_29563;
        rob_val_2_6 <= ~_GEN_2816 & _GEN_29562;
        rob_val_2_5 <= ~_GEN_2815 & _GEN_29561;
        rob_val_2_4 <= ~_GEN_2814 & _GEN_29560;
        rob_val_2_3 <= ~_GEN_2813 & _GEN_29559;
        rob_val_2_2 <= ~_GEN_2812 & _GEN_29558;
        rob_val_2_1 <= ~_GEN_2811 & _GEN_29557;
        rob_val_2_0 <= ~_GEN_2810 & _GEN_29556;
      end
      if (_io_commit_valids_3_output) begin
        rob_val_3_31 <= ~((&rob_head) | _GEN_2937) & _GEN_42951;
        rob_val_3_30 <= ~(_GEN_2317 | _GEN_2936) & _GEN_42950;
        rob_val_3_29 <= ~(_GEN_2316 | _GEN_2935) & _GEN_42949;
        rob_val_3_28 <= ~(_GEN_2315 | _GEN_2934) & _GEN_42948;
        rob_val_3_27 <= ~(_GEN_2314 | _GEN_2933) & _GEN_42947;
        rob_val_3_26 <= ~(_GEN_2313 | _GEN_2932) & _GEN_42946;
        rob_val_3_25 <= ~(_GEN_2312 | _GEN_2931) & _GEN_42945;
        rob_val_3_24 <= ~(_GEN_2311 | _GEN_2930) & _GEN_42944;
        rob_val_3_23 <= ~(_GEN_2310 | _GEN_2929) & _GEN_42943;
        rob_val_3_22 <= ~(_GEN_2309 | _GEN_2928) & _GEN_42942;
        rob_val_3_21 <= ~(_GEN_2308 | _GEN_2927) & _GEN_42941;
        rob_val_3_20 <= ~(_GEN_2307 | _GEN_2926) & _GEN_42940;
        rob_val_3_19 <= ~(_GEN_2306 | _GEN_2925) & _GEN_42939;
        rob_val_3_18 <= ~(_GEN_2305 | _GEN_2924) & _GEN_42938;
        rob_val_3_17 <= ~(_GEN_2304 | _GEN_2923) & _GEN_42937;
        rob_val_3_16 <= ~(_GEN_2303 | _GEN_2922) & _GEN_42936;
        rob_val_3_15 <= ~(_GEN_2302 | _GEN_2921) & _GEN_42935;
        rob_val_3_14 <= ~(_GEN_2301 | _GEN_2920) & _GEN_42934;
        rob_val_3_13 <= ~(_GEN_2300 | _GEN_2919) & _GEN_42933;
        rob_val_3_12 <= ~(_GEN_2299 | _GEN_2918) & _GEN_42932;
        rob_val_3_11 <= ~(_GEN_2298 | _GEN_2917) & _GEN_42931;
        rob_val_3_10 <= ~(_GEN_2297 | _GEN_2916) & _GEN_42930;
        rob_val_3_9 <= ~(_GEN_2296 | _GEN_2915) & _GEN_42929;
        rob_val_3_8 <= ~(_GEN_2295 | _GEN_2914) & _GEN_42928;
        rob_val_3_7 <= ~(_GEN_2294 | _GEN_2913) & _GEN_42927;
        rob_val_3_6 <= ~(_GEN_2293 | _GEN_2912) & _GEN_42926;
        rob_val_3_5 <= ~(_GEN_2292 | _GEN_2911) & _GEN_42925;
        rob_val_3_4 <= ~(_GEN_2291 | _GEN_2910) & _GEN_42924;
        rob_val_3_3 <= ~(_GEN_2290 | _GEN_2909) & _GEN_42923;
        rob_val_3_2 <= ~(_GEN_2289 | _GEN_2908) & _GEN_42922;
        rob_val_3_1 <= ~(_GEN_2288 | _GEN_2907) & _GEN_42921;
        rob_val_3_0 <= ~(_GEN_2318 | _GEN_2906) & _GEN_42920;
      end
      else begin
        rob_val_3_31 <= ~_GEN_2937 & _GEN_42951;
        rob_val_3_30 <= ~_GEN_2936 & _GEN_42950;
        rob_val_3_29 <= ~_GEN_2935 & _GEN_42949;
        rob_val_3_28 <= ~_GEN_2934 & _GEN_42948;
        rob_val_3_27 <= ~_GEN_2933 & _GEN_42947;
        rob_val_3_26 <= ~_GEN_2932 & _GEN_42946;
        rob_val_3_25 <= ~_GEN_2931 & _GEN_42945;
        rob_val_3_24 <= ~_GEN_2930 & _GEN_42944;
        rob_val_3_23 <= ~_GEN_2929 & _GEN_42943;
        rob_val_3_22 <= ~_GEN_2928 & _GEN_42942;
        rob_val_3_21 <= ~_GEN_2927 & _GEN_42941;
        rob_val_3_20 <= ~_GEN_2926 & _GEN_42940;
        rob_val_3_19 <= ~_GEN_2925 & _GEN_42939;
        rob_val_3_18 <= ~_GEN_2924 & _GEN_42938;
        rob_val_3_17 <= ~_GEN_2923 & _GEN_42937;
        rob_val_3_16 <= ~_GEN_2922 & _GEN_42936;
        rob_val_3_15 <= ~_GEN_2921 & _GEN_42935;
        rob_val_3_14 <= ~_GEN_2920 & _GEN_42934;
        rob_val_3_13 <= ~_GEN_2919 & _GEN_42933;
        rob_val_3_12 <= ~_GEN_2918 & _GEN_42932;
        rob_val_3_11 <= ~_GEN_2917 & _GEN_42931;
        rob_val_3_10 <= ~_GEN_2916 & _GEN_42930;
        rob_val_3_9 <= ~_GEN_2915 & _GEN_42929;
        rob_val_3_8 <= ~_GEN_2914 & _GEN_42928;
        rob_val_3_7 <= ~_GEN_2913 & _GEN_42927;
        rob_val_3_6 <= ~_GEN_2912 & _GEN_42926;
        rob_val_3_5 <= ~_GEN_2911 & _GEN_42925;
        rob_val_3_4 <= ~_GEN_2910 & _GEN_42924;
        rob_val_3_3 <= ~_GEN_2909 & _GEN_42923;
        rob_val_3_2 <= ~_GEN_2908 & _GEN_42922;
        rob_val_3_1 <= ~_GEN_2907 & _GEN_42921;
        rob_val_3_0 <= ~_GEN_2906 & _GEN_42920;
      end
      if (io_enq_valids_0 | io_enq_valids_1 | io_enq_valids_2 | io_enq_valids_3)
        r_partial_row <= io_enq_partial_stall;
    end
    r_xcpt_uop_br_mask <= next_xcpt_uop_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_2743) begin
      if (io_lxcpt_valid) begin
        if (_GEN_2744) begin
          r_xcpt_uop_rob_idx <= io_lxcpt_bits_uop_rob_idx;
          r_xcpt_uop_exc_cause <= {59'h0, io_lxcpt_bits_cause};
          r_xcpt_badvaddr <= io_lxcpt_bits_badvaddr;
        end
      end
      else if (_GEN_2745) begin
        r_xcpt_uop_rob_idx <= casez_tmp_93;
        r_xcpt_uop_exc_cause <= casez_tmp_94;
        r_xcpt_badvaddr <= {io_xcpt_fetch_pc[39:6], casez_tmp_92};
      end
    end
    rob_bsy__31 <= ~_GEN_896 & (_GEN_769 ? ~_GEN_832 & _GEN_7403 : ~_GEN_768 & _GEN_7403);
    rob_bsy__30 <= ~_GEN_895 & (_GEN_769 ? ~_GEN_831 & _GEN_7402 : ~_GEN_767 & _GEN_7402);
    rob_bsy__29 <= ~_GEN_894 & (_GEN_769 ? ~_GEN_829 & _GEN_7401 : ~_GEN_766 & _GEN_7401);
    rob_bsy__28 <= ~_GEN_893 & (_GEN_769 ? ~_GEN_827 & _GEN_7400 : ~_GEN_765 & _GEN_7400);
    rob_bsy__27 <= ~_GEN_892 & (_GEN_769 ? ~_GEN_825 & _GEN_7399 : ~_GEN_764 & _GEN_7399);
    rob_bsy__26 <= ~_GEN_891 & (_GEN_769 ? ~_GEN_823 & _GEN_7398 : ~_GEN_763 & _GEN_7398);
    rob_bsy__25 <= ~_GEN_890 & (_GEN_769 ? ~_GEN_821 & _GEN_7397 : ~_GEN_762 & _GEN_7397);
    rob_bsy__24 <= ~_GEN_889 & (_GEN_769 ? ~_GEN_819 & _GEN_7396 : ~_GEN_761 & _GEN_7396);
    rob_bsy__23 <= ~_GEN_888 & (_GEN_769 ? ~_GEN_817 & _GEN_7395 : ~_GEN_760 & _GEN_7395);
    rob_bsy__22 <= ~_GEN_887 & (_GEN_769 ? ~_GEN_815 & _GEN_7394 : ~_GEN_759 & _GEN_7394);
    rob_bsy__21 <= ~_GEN_886 & (_GEN_769 ? ~_GEN_813 & _GEN_7393 : ~_GEN_758 & _GEN_7393);
    rob_bsy__20 <= ~_GEN_885 & (_GEN_769 ? ~_GEN_811 & _GEN_7392 : ~_GEN_757 & _GEN_7392);
    rob_bsy__19 <= ~_GEN_884 & (_GEN_769 ? ~_GEN_809 & _GEN_7391 : ~_GEN_756 & _GEN_7391);
    rob_bsy__18 <= ~_GEN_883 & (_GEN_769 ? ~_GEN_807 & _GEN_7390 : ~_GEN_755 & _GEN_7390);
    rob_bsy__17 <= ~_GEN_882 & (_GEN_769 ? ~_GEN_805 & _GEN_7389 : ~_GEN_754 & _GEN_7389);
    rob_bsy__16 <= ~_GEN_881 & (_GEN_769 ? ~_GEN_803 & _GEN_7388 : ~_GEN_753 & _GEN_7388);
    rob_bsy__15 <= ~_GEN_880 & (_GEN_769 ? ~_GEN_801 & _GEN_7387 : ~_GEN_752 & _GEN_7387);
    rob_bsy__14 <= ~_GEN_879 & (_GEN_769 ? ~_GEN_799 & _GEN_7386 : ~_GEN_751 & _GEN_7386);
    rob_bsy__13 <= ~_GEN_878 & (_GEN_769 ? ~_GEN_797 & _GEN_7385 : ~_GEN_750 & _GEN_7385);
    rob_bsy__12 <= ~_GEN_877 & (_GEN_769 ? ~_GEN_795 & _GEN_7384 : ~_GEN_749 & _GEN_7384);
    rob_bsy__11 <= ~_GEN_876 & (_GEN_769 ? ~_GEN_793 & _GEN_7383 : ~_GEN_748 & _GEN_7383);
    rob_bsy__10 <= ~_GEN_875 & (_GEN_769 ? ~_GEN_791 & _GEN_7382 : ~_GEN_747 & _GEN_7382);
    rob_bsy__9 <= ~_GEN_874 & (_GEN_769 ? ~_GEN_789 & _GEN_7381 : ~_GEN_746 & _GEN_7381);
    rob_bsy__8 <= ~_GEN_873 & (_GEN_769 ? ~_GEN_787 & _GEN_7380 : ~_GEN_745 & _GEN_7380);
    rob_bsy__7 <= ~_GEN_872 & (_GEN_769 ? ~_GEN_785 & _GEN_7379 : ~_GEN_744 & _GEN_7379);
    rob_bsy__6 <= ~_GEN_871 & (_GEN_769 ? ~_GEN_783 & _GEN_7378 : ~_GEN_743 & _GEN_7378);
    rob_bsy__5 <= ~_GEN_870 & (_GEN_769 ? ~_GEN_781 & _GEN_7377 : ~_GEN_742 & _GEN_7377);
    rob_bsy__4 <= ~_GEN_869 & (_GEN_769 ? ~_GEN_779 & _GEN_7376 : ~_GEN_741 & _GEN_7376);
    rob_bsy__3 <= ~_GEN_868 & (_GEN_769 ? ~_GEN_777 & _GEN_7375 : ~_GEN_740 & _GEN_7375);
    rob_bsy__2 <= ~_GEN_867 & (_GEN_769 ? ~_GEN_775 & _GEN_7374 : ~_GEN_739 & _GEN_7374);
    rob_bsy__1 <= ~_GEN_866 & (_GEN_769 ? ~_GEN_773 & _GEN_7373 : ~_GEN_738 & _GEN_7373);
    rob_bsy__0 <= ~_GEN_865 & (_GEN_769 ? ~_GEN_771 & _GEN_7372 : ~_GEN_737 & _GEN_7372);
    rob_exception__31 <= ~_GEN_2509 & (_GEN_897 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_64 ? io_enq_uops_0_exception : rob_exception__31));
    rob_exception__30 <= ~_GEN_2508 & (_GEN_897 & _GEN_2446 | (_GEN_63 ? io_enq_uops_0_exception : rob_exception__30));
    rob_exception__29 <= ~_GEN_2507 & (_GEN_897 & _GEN_2445 | (_GEN_62 ? io_enq_uops_0_exception : rob_exception__29));
    rob_exception__28 <= ~_GEN_2506 & (_GEN_897 & _GEN_2444 | (_GEN_61 ? io_enq_uops_0_exception : rob_exception__28));
    rob_exception__27 <= ~_GEN_2505 & (_GEN_897 & _GEN_2443 | (_GEN_60 ? io_enq_uops_0_exception : rob_exception__27));
    rob_exception__26 <= ~_GEN_2504 & (_GEN_897 & _GEN_2442 | (_GEN_59 ? io_enq_uops_0_exception : rob_exception__26));
    rob_exception__25 <= ~_GEN_2503 & (_GEN_897 & _GEN_2441 | (_GEN_58 ? io_enq_uops_0_exception : rob_exception__25));
    rob_exception__24 <= ~_GEN_2502 & (_GEN_897 & _GEN_2440 | (_GEN_57 ? io_enq_uops_0_exception : rob_exception__24));
    rob_exception__23 <= ~_GEN_2501 & (_GEN_897 & _GEN_2439 | (_GEN_56 ? io_enq_uops_0_exception : rob_exception__23));
    rob_exception__22 <= ~_GEN_2500 & (_GEN_897 & _GEN_2438 | (_GEN_55 ? io_enq_uops_0_exception : rob_exception__22));
    rob_exception__21 <= ~_GEN_2499 & (_GEN_897 & _GEN_2437 | (_GEN_54 ? io_enq_uops_0_exception : rob_exception__21));
    rob_exception__20 <= ~_GEN_2498 & (_GEN_897 & _GEN_2436 | (_GEN_53 ? io_enq_uops_0_exception : rob_exception__20));
    rob_exception__19 <= ~_GEN_2497 & (_GEN_897 & _GEN_2435 | (_GEN_52 ? io_enq_uops_0_exception : rob_exception__19));
    rob_exception__18 <= ~_GEN_2496 & (_GEN_897 & _GEN_2434 | (_GEN_51 ? io_enq_uops_0_exception : rob_exception__18));
    rob_exception__17 <= ~_GEN_2495 & (_GEN_897 & _GEN_2433 | (_GEN_50 ? io_enq_uops_0_exception : rob_exception__17));
    rob_exception__16 <= ~_GEN_2494 & (_GEN_897 & _GEN_2432 | (_GEN_49 ? io_enq_uops_0_exception : rob_exception__16));
    rob_exception__15 <= ~_GEN_2493 & (_GEN_897 & _GEN_2431 | (_GEN_48 ? io_enq_uops_0_exception : rob_exception__15));
    rob_exception__14 <= ~_GEN_2492 & (_GEN_897 & _GEN_2430 | (_GEN_47 ? io_enq_uops_0_exception : rob_exception__14));
    rob_exception__13 <= ~_GEN_2491 & (_GEN_897 & _GEN_2429 | (_GEN_46 ? io_enq_uops_0_exception : rob_exception__13));
    rob_exception__12 <= ~_GEN_2490 & (_GEN_897 & _GEN_2428 | (_GEN_45 ? io_enq_uops_0_exception : rob_exception__12));
    rob_exception__11 <= ~_GEN_2489 & (_GEN_897 & _GEN_2427 | (_GEN_44 ? io_enq_uops_0_exception : rob_exception__11));
    rob_exception__10 <= ~_GEN_2488 & (_GEN_897 & _GEN_2426 | (_GEN_43 ? io_enq_uops_0_exception : rob_exception__10));
    rob_exception__9 <= ~_GEN_2487 & (_GEN_897 & _GEN_2425 | (_GEN_42 ? io_enq_uops_0_exception : rob_exception__9));
    rob_exception__8 <= ~_GEN_2486 & (_GEN_897 & _GEN_2424 | (_GEN_41 ? io_enq_uops_0_exception : rob_exception__8));
    rob_exception__7 <= ~_GEN_2485 & (_GEN_897 & _GEN_2423 | (_GEN_40 ? io_enq_uops_0_exception : rob_exception__7));
    rob_exception__6 <= ~_GEN_2484 & (_GEN_897 & _GEN_2422 | (_GEN_39 ? io_enq_uops_0_exception : rob_exception__6));
    rob_exception__5 <= ~_GEN_2483 & (_GEN_897 & _GEN_2421 | (_GEN_38 ? io_enq_uops_0_exception : rob_exception__5));
    rob_exception__4 <= ~_GEN_2482 & (_GEN_897 & _GEN_2420 | (_GEN_37 ? io_enq_uops_0_exception : rob_exception__4));
    rob_exception__3 <= ~_GEN_2481 & (_GEN_897 & _GEN_2419 | (_GEN_36 ? io_enq_uops_0_exception : rob_exception__3));
    rob_exception__2 <= ~_GEN_2480 & (_GEN_897 & _GEN_2418 | (_GEN_35 ? io_enq_uops_0_exception : rob_exception__2));
    rob_exception__1 <= ~_GEN_2479 & (_GEN_897 & _GEN_2417 | (_GEN_34 ? io_enq_uops_0_exception : rob_exception__1));
    rob_exception__0 <= ~_GEN_2478 & (_GEN_897 & _GEN_2416 | (_GEN_33 ? io_enq_uops_0_exception : rob_exception__0));
    block_commit_REG <= exception_thrown;
    block_commit_REG_2 <= block_commit_REG_1;
    rob_bsy_1_31 <= ~_GEN_1358 & (_GEN_1293 ? ~_GEN_1325 & _GEN_20767 : ~_GEN_1292 & _GEN_20767);
    rob_bsy_1_30 <= ~_GEN_1357 & (_GEN_1293 ? ~_GEN_1324 & _GEN_20766 : ~_GEN_1291 & _GEN_20766);
    rob_bsy_1_29 <= ~_GEN_1356 & (_GEN_1293 ? ~_GEN_1323 & _GEN_20765 : ~_GEN_1290 & _GEN_20765);
    rob_bsy_1_28 <= ~_GEN_1355 & (_GEN_1293 ? ~_GEN_1322 & _GEN_20764 : ~_GEN_1289 & _GEN_20764);
    rob_bsy_1_27 <= ~_GEN_1354 & (_GEN_1293 ? ~_GEN_1321 & _GEN_20763 : ~_GEN_1288 & _GEN_20763);
    rob_bsy_1_26 <= ~_GEN_1353 & (_GEN_1293 ? ~_GEN_1320 & _GEN_20762 : ~_GEN_1287 & _GEN_20762);
    rob_bsy_1_25 <= ~_GEN_1352 & (_GEN_1293 ? ~_GEN_1319 & _GEN_20761 : ~_GEN_1286 & _GEN_20761);
    rob_bsy_1_24 <= ~_GEN_1351 & (_GEN_1293 ? ~_GEN_1318 & _GEN_20760 : ~_GEN_1285 & _GEN_20760);
    rob_bsy_1_23 <= ~_GEN_1350 & (_GEN_1293 ? ~_GEN_1317 & _GEN_20759 : ~_GEN_1284 & _GEN_20759);
    rob_bsy_1_22 <= ~_GEN_1349 & (_GEN_1293 ? ~_GEN_1316 & _GEN_20758 : ~_GEN_1283 & _GEN_20758);
    rob_bsy_1_21 <= ~_GEN_1348 & (_GEN_1293 ? ~_GEN_1315 & _GEN_20757 : ~_GEN_1282 & _GEN_20757);
    rob_bsy_1_20 <= ~_GEN_1347 & (_GEN_1293 ? ~_GEN_1314 & _GEN_20756 : ~_GEN_1281 & _GEN_20756);
    rob_bsy_1_19 <= ~_GEN_1346 & (_GEN_1293 ? ~_GEN_1313 & _GEN_20755 : ~_GEN_1280 & _GEN_20755);
    rob_bsy_1_18 <= ~_GEN_1345 & (_GEN_1293 ? ~_GEN_1312 & _GEN_20754 : ~_GEN_1279 & _GEN_20754);
    rob_bsy_1_17 <= ~_GEN_1344 & (_GEN_1293 ? ~_GEN_1311 & _GEN_20753 : ~_GEN_1278 & _GEN_20753);
    rob_bsy_1_16 <= ~_GEN_1343 & (_GEN_1293 ? ~_GEN_1310 & _GEN_20752 : ~_GEN_1277 & _GEN_20752);
    rob_bsy_1_15 <= ~_GEN_1342 & (_GEN_1293 ? ~_GEN_1309 & _GEN_20751 : ~_GEN_1276 & _GEN_20751);
    rob_bsy_1_14 <= ~_GEN_1341 & (_GEN_1293 ? ~_GEN_1308 & _GEN_20750 : ~_GEN_1275 & _GEN_20750);
    rob_bsy_1_13 <= ~_GEN_1340 & (_GEN_1293 ? ~_GEN_1307 & _GEN_20749 : ~_GEN_1274 & _GEN_20749);
    rob_bsy_1_12 <= ~_GEN_1339 & (_GEN_1293 ? ~_GEN_1306 & _GEN_20748 : ~_GEN_1273 & _GEN_20748);
    rob_bsy_1_11 <= ~_GEN_1338 & (_GEN_1293 ? ~_GEN_1305 & _GEN_20747 : ~_GEN_1272 & _GEN_20747);
    rob_bsy_1_10 <= ~_GEN_1337 & (_GEN_1293 ? ~_GEN_1304 & _GEN_20746 : ~_GEN_1271 & _GEN_20746);
    rob_bsy_1_9 <= ~_GEN_1336 & (_GEN_1293 ? ~_GEN_1303 & _GEN_20745 : ~_GEN_1270 & _GEN_20745);
    rob_bsy_1_8 <= ~_GEN_1335 & (_GEN_1293 ? ~_GEN_1302 & _GEN_20744 : ~_GEN_1269 & _GEN_20744);
    rob_bsy_1_7 <= ~_GEN_1334 & (_GEN_1293 ? ~_GEN_1301 & _GEN_20743 : ~_GEN_1268 & _GEN_20743);
    rob_bsy_1_6 <= ~_GEN_1333 & (_GEN_1293 ? ~_GEN_1300 & _GEN_20742 : ~_GEN_1267 & _GEN_20742);
    rob_bsy_1_5 <= ~_GEN_1332 & (_GEN_1293 ? ~_GEN_1299 & _GEN_20741 : ~_GEN_1266 & _GEN_20741);
    rob_bsy_1_4 <= ~_GEN_1331 & (_GEN_1293 ? ~_GEN_1298 & _GEN_20740 : ~_GEN_1265 & _GEN_20740);
    rob_bsy_1_3 <= ~_GEN_1330 & (_GEN_1293 ? ~_GEN_1297 & _GEN_20739 : ~_GEN_1264 & _GEN_20739);
    rob_bsy_1_2 <= ~_GEN_1329 & (_GEN_1293 ? ~_GEN_1296 & _GEN_20738 : ~_GEN_1263 & _GEN_20738);
    rob_bsy_1_1 <= ~_GEN_1328 & (_GEN_1293 ? ~_GEN_1295 & _GEN_20737 : ~_GEN_1262 & _GEN_20737);
    rob_bsy_1_0 <= ~_GEN_1327 & (_GEN_1293 ? ~_GEN_1294 & _GEN_20736 : ~_GEN_1261 & _GEN_20736);
    rob_exception_1_31 <= ~_GEN_2576 & (_GEN_1359 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_929 ? io_enq_uops_1_exception : rob_exception_1_31));
    rob_exception_1_30 <= ~_GEN_2575 & (_GEN_1359 & _GEN_2446 | (_GEN_928 ? io_enq_uops_1_exception : rob_exception_1_30));
    rob_exception_1_29 <= ~_GEN_2574 & (_GEN_1359 & _GEN_2445 | (_GEN_927 ? io_enq_uops_1_exception : rob_exception_1_29));
    rob_exception_1_28 <= ~_GEN_2573 & (_GEN_1359 & _GEN_2444 | (_GEN_926 ? io_enq_uops_1_exception : rob_exception_1_28));
    rob_exception_1_27 <= ~_GEN_2572 & (_GEN_1359 & _GEN_2443 | (_GEN_925 ? io_enq_uops_1_exception : rob_exception_1_27));
    rob_exception_1_26 <= ~_GEN_2571 & (_GEN_1359 & _GEN_2442 | (_GEN_924 ? io_enq_uops_1_exception : rob_exception_1_26));
    rob_exception_1_25 <= ~_GEN_2570 & (_GEN_1359 & _GEN_2441 | (_GEN_923 ? io_enq_uops_1_exception : rob_exception_1_25));
    rob_exception_1_24 <= ~_GEN_2569 & (_GEN_1359 & _GEN_2440 | (_GEN_922 ? io_enq_uops_1_exception : rob_exception_1_24));
    rob_exception_1_23 <= ~_GEN_2568 & (_GEN_1359 & _GEN_2439 | (_GEN_921 ? io_enq_uops_1_exception : rob_exception_1_23));
    rob_exception_1_22 <= ~_GEN_2567 & (_GEN_1359 & _GEN_2438 | (_GEN_920 ? io_enq_uops_1_exception : rob_exception_1_22));
    rob_exception_1_21 <= ~_GEN_2566 & (_GEN_1359 & _GEN_2437 | (_GEN_919 ? io_enq_uops_1_exception : rob_exception_1_21));
    rob_exception_1_20 <= ~_GEN_2565 & (_GEN_1359 & _GEN_2436 | (_GEN_918 ? io_enq_uops_1_exception : rob_exception_1_20));
    rob_exception_1_19 <= ~_GEN_2564 & (_GEN_1359 & _GEN_2435 | (_GEN_917 ? io_enq_uops_1_exception : rob_exception_1_19));
    rob_exception_1_18 <= ~_GEN_2563 & (_GEN_1359 & _GEN_2434 | (_GEN_916 ? io_enq_uops_1_exception : rob_exception_1_18));
    rob_exception_1_17 <= ~_GEN_2562 & (_GEN_1359 & _GEN_2433 | (_GEN_915 ? io_enq_uops_1_exception : rob_exception_1_17));
    rob_exception_1_16 <= ~_GEN_2561 & (_GEN_1359 & _GEN_2432 | (_GEN_914 ? io_enq_uops_1_exception : rob_exception_1_16));
    rob_exception_1_15 <= ~_GEN_2560 & (_GEN_1359 & _GEN_2431 | (_GEN_913 ? io_enq_uops_1_exception : rob_exception_1_15));
    rob_exception_1_14 <= ~_GEN_2559 & (_GEN_1359 & _GEN_2430 | (_GEN_912 ? io_enq_uops_1_exception : rob_exception_1_14));
    rob_exception_1_13 <= ~_GEN_2558 & (_GEN_1359 & _GEN_2429 | (_GEN_911 ? io_enq_uops_1_exception : rob_exception_1_13));
    rob_exception_1_12 <= ~_GEN_2557 & (_GEN_1359 & _GEN_2428 | (_GEN_910 ? io_enq_uops_1_exception : rob_exception_1_12));
    rob_exception_1_11 <= ~_GEN_2556 & (_GEN_1359 & _GEN_2427 | (_GEN_909 ? io_enq_uops_1_exception : rob_exception_1_11));
    rob_exception_1_10 <= ~_GEN_2555 & (_GEN_1359 & _GEN_2426 | (_GEN_908 ? io_enq_uops_1_exception : rob_exception_1_10));
    rob_exception_1_9 <= ~_GEN_2554 & (_GEN_1359 & _GEN_2425 | (_GEN_907 ? io_enq_uops_1_exception : rob_exception_1_9));
    rob_exception_1_8 <= ~_GEN_2553 & (_GEN_1359 & _GEN_2424 | (_GEN_906 ? io_enq_uops_1_exception : rob_exception_1_8));
    rob_exception_1_7 <= ~_GEN_2552 & (_GEN_1359 & _GEN_2423 | (_GEN_905 ? io_enq_uops_1_exception : rob_exception_1_7));
    rob_exception_1_6 <= ~_GEN_2551 & (_GEN_1359 & _GEN_2422 | (_GEN_904 ? io_enq_uops_1_exception : rob_exception_1_6));
    rob_exception_1_5 <= ~_GEN_2550 & (_GEN_1359 & _GEN_2421 | (_GEN_903 ? io_enq_uops_1_exception : rob_exception_1_5));
    rob_exception_1_4 <= ~_GEN_2549 & (_GEN_1359 & _GEN_2420 | (_GEN_902 ? io_enq_uops_1_exception : rob_exception_1_4));
    rob_exception_1_3 <= ~_GEN_2548 & (_GEN_1359 & _GEN_2419 | (_GEN_901 ? io_enq_uops_1_exception : rob_exception_1_3));
    rob_exception_1_2 <= ~_GEN_2547 & (_GEN_1359 & _GEN_2418 | (_GEN_900 ? io_enq_uops_1_exception : rob_exception_1_2));
    rob_exception_1_1 <= ~_GEN_2546 & (_GEN_1359 & _GEN_2417 | (_GEN_899 ? io_enq_uops_1_exception : rob_exception_1_1));
    rob_exception_1_0 <= ~_GEN_2545 & (_GEN_1359 & _GEN_2416 | (_GEN_898 ? io_enq_uops_1_exception : rob_exception_1_0));
    rob_bsy_2_31 <= ~_GEN_1820 & (_GEN_1755 ? ~_GEN_1787 & _GEN_34131 : ~_GEN_1754 & _GEN_34131);
    rob_bsy_2_30 <= ~_GEN_1819 & (_GEN_1755 ? ~_GEN_1786 & _GEN_34130 : ~_GEN_1753 & _GEN_34130);
    rob_bsy_2_29 <= ~_GEN_1818 & (_GEN_1755 ? ~_GEN_1785 & _GEN_34129 : ~_GEN_1752 & _GEN_34129);
    rob_bsy_2_28 <= ~_GEN_1817 & (_GEN_1755 ? ~_GEN_1784 & _GEN_34128 : ~_GEN_1751 & _GEN_34128);
    rob_bsy_2_27 <= ~_GEN_1816 & (_GEN_1755 ? ~_GEN_1783 & _GEN_34127 : ~_GEN_1750 & _GEN_34127);
    rob_bsy_2_26 <= ~_GEN_1815 & (_GEN_1755 ? ~_GEN_1782 & _GEN_34126 : ~_GEN_1749 & _GEN_34126);
    rob_bsy_2_25 <= ~_GEN_1814 & (_GEN_1755 ? ~_GEN_1781 & _GEN_34125 : ~_GEN_1748 & _GEN_34125);
    rob_bsy_2_24 <= ~_GEN_1813 & (_GEN_1755 ? ~_GEN_1780 & _GEN_34124 : ~_GEN_1747 & _GEN_34124);
    rob_bsy_2_23 <= ~_GEN_1812 & (_GEN_1755 ? ~_GEN_1779 & _GEN_34123 : ~_GEN_1746 & _GEN_34123);
    rob_bsy_2_22 <= ~_GEN_1811 & (_GEN_1755 ? ~_GEN_1778 & _GEN_34122 : ~_GEN_1745 & _GEN_34122);
    rob_bsy_2_21 <= ~_GEN_1810 & (_GEN_1755 ? ~_GEN_1777 & _GEN_34121 : ~_GEN_1744 & _GEN_34121);
    rob_bsy_2_20 <= ~_GEN_1809 & (_GEN_1755 ? ~_GEN_1776 & _GEN_34120 : ~_GEN_1743 & _GEN_34120);
    rob_bsy_2_19 <= ~_GEN_1808 & (_GEN_1755 ? ~_GEN_1775 & _GEN_34119 : ~_GEN_1742 & _GEN_34119);
    rob_bsy_2_18 <= ~_GEN_1807 & (_GEN_1755 ? ~_GEN_1774 & _GEN_34118 : ~_GEN_1741 & _GEN_34118);
    rob_bsy_2_17 <= ~_GEN_1806 & (_GEN_1755 ? ~_GEN_1773 & _GEN_34117 : ~_GEN_1740 & _GEN_34117);
    rob_bsy_2_16 <= ~_GEN_1805 & (_GEN_1755 ? ~_GEN_1772 & _GEN_34116 : ~_GEN_1739 & _GEN_34116);
    rob_bsy_2_15 <= ~_GEN_1804 & (_GEN_1755 ? ~_GEN_1771 & _GEN_34115 : ~_GEN_1738 & _GEN_34115);
    rob_bsy_2_14 <= ~_GEN_1803 & (_GEN_1755 ? ~_GEN_1770 & _GEN_34114 : ~_GEN_1737 & _GEN_34114);
    rob_bsy_2_13 <= ~_GEN_1802 & (_GEN_1755 ? ~_GEN_1769 & _GEN_34113 : ~_GEN_1736 & _GEN_34113);
    rob_bsy_2_12 <= ~_GEN_1801 & (_GEN_1755 ? ~_GEN_1768 & _GEN_34112 : ~_GEN_1735 & _GEN_34112);
    rob_bsy_2_11 <= ~_GEN_1800 & (_GEN_1755 ? ~_GEN_1767 & _GEN_34111 : ~_GEN_1734 & _GEN_34111);
    rob_bsy_2_10 <= ~_GEN_1799 & (_GEN_1755 ? ~_GEN_1766 & _GEN_34110 : ~_GEN_1733 & _GEN_34110);
    rob_bsy_2_9 <= ~_GEN_1798 & (_GEN_1755 ? ~_GEN_1765 & _GEN_34109 : ~_GEN_1732 & _GEN_34109);
    rob_bsy_2_8 <= ~_GEN_1797 & (_GEN_1755 ? ~_GEN_1764 & _GEN_34108 : ~_GEN_1731 & _GEN_34108);
    rob_bsy_2_7 <= ~_GEN_1796 & (_GEN_1755 ? ~_GEN_1763 & _GEN_34107 : ~_GEN_1730 & _GEN_34107);
    rob_bsy_2_6 <= ~_GEN_1795 & (_GEN_1755 ? ~_GEN_1762 & _GEN_34106 : ~_GEN_1729 & _GEN_34106);
    rob_bsy_2_5 <= ~_GEN_1794 & (_GEN_1755 ? ~_GEN_1761 & _GEN_34105 : ~_GEN_1728 & _GEN_34105);
    rob_bsy_2_4 <= ~_GEN_1793 & (_GEN_1755 ? ~_GEN_1760 & _GEN_34104 : ~_GEN_1727 & _GEN_34104);
    rob_bsy_2_3 <= ~_GEN_1792 & (_GEN_1755 ? ~_GEN_1759 & _GEN_34103 : ~_GEN_1726 & _GEN_34103);
    rob_bsy_2_2 <= ~_GEN_1791 & (_GEN_1755 ? ~_GEN_1758 & _GEN_34102 : ~_GEN_1725 & _GEN_34102);
    rob_bsy_2_1 <= ~_GEN_1790 & (_GEN_1755 ? ~_GEN_1757 & _GEN_34101 : ~_GEN_1724 & _GEN_34101);
    rob_bsy_2_0 <= ~_GEN_1789 & (_GEN_1755 ? ~_GEN_1756 & _GEN_34100 : ~_GEN_1723 & _GEN_34100);
    rob_exception_2_31 <= ~_GEN_2643 & (_GEN_1821 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_1391 ? io_enq_uops_2_exception : rob_exception_2_31));
    rob_exception_2_30 <= ~_GEN_2642 & (_GEN_1821 & _GEN_2446 | (_GEN_1390 ? io_enq_uops_2_exception : rob_exception_2_30));
    rob_exception_2_29 <= ~_GEN_2641 & (_GEN_1821 & _GEN_2445 | (_GEN_1389 ? io_enq_uops_2_exception : rob_exception_2_29));
    rob_exception_2_28 <= ~_GEN_2640 & (_GEN_1821 & _GEN_2444 | (_GEN_1388 ? io_enq_uops_2_exception : rob_exception_2_28));
    rob_exception_2_27 <= ~_GEN_2639 & (_GEN_1821 & _GEN_2443 | (_GEN_1387 ? io_enq_uops_2_exception : rob_exception_2_27));
    rob_exception_2_26 <= ~_GEN_2638 & (_GEN_1821 & _GEN_2442 | (_GEN_1386 ? io_enq_uops_2_exception : rob_exception_2_26));
    rob_exception_2_25 <= ~_GEN_2637 & (_GEN_1821 & _GEN_2441 | (_GEN_1385 ? io_enq_uops_2_exception : rob_exception_2_25));
    rob_exception_2_24 <= ~_GEN_2636 & (_GEN_1821 & _GEN_2440 | (_GEN_1384 ? io_enq_uops_2_exception : rob_exception_2_24));
    rob_exception_2_23 <= ~_GEN_2635 & (_GEN_1821 & _GEN_2439 | (_GEN_1383 ? io_enq_uops_2_exception : rob_exception_2_23));
    rob_exception_2_22 <= ~_GEN_2634 & (_GEN_1821 & _GEN_2438 | (_GEN_1382 ? io_enq_uops_2_exception : rob_exception_2_22));
    rob_exception_2_21 <= ~_GEN_2633 & (_GEN_1821 & _GEN_2437 | (_GEN_1381 ? io_enq_uops_2_exception : rob_exception_2_21));
    rob_exception_2_20 <= ~_GEN_2632 & (_GEN_1821 & _GEN_2436 | (_GEN_1380 ? io_enq_uops_2_exception : rob_exception_2_20));
    rob_exception_2_19 <= ~_GEN_2631 & (_GEN_1821 & _GEN_2435 | (_GEN_1379 ? io_enq_uops_2_exception : rob_exception_2_19));
    rob_exception_2_18 <= ~_GEN_2630 & (_GEN_1821 & _GEN_2434 | (_GEN_1378 ? io_enq_uops_2_exception : rob_exception_2_18));
    rob_exception_2_17 <= ~_GEN_2629 & (_GEN_1821 & _GEN_2433 | (_GEN_1377 ? io_enq_uops_2_exception : rob_exception_2_17));
    rob_exception_2_16 <= ~_GEN_2628 & (_GEN_1821 & _GEN_2432 | (_GEN_1376 ? io_enq_uops_2_exception : rob_exception_2_16));
    rob_exception_2_15 <= ~_GEN_2627 & (_GEN_1821 & _GEN_2431 | (_GEN_1375 ? io_enq_uops_2_exception : rob_exception_2_15));
    rob_exception_2_14 <= ~_GEN_2626 & (_GEN_1821 & _GEN_2430 | (_GEN_1374 ? io_enq_uops_2_exception : rob_exception_2_14));
    rob_exception_2_13 <= ~_GEN_2625 & (_GEN_1821 & _GEN_2429 | (_GEN_1373 ? io_enq_uops_2_exception : rob_exception_2_13));
    rob_exception_2_12 <= ~_GEN_2624 & (_GEN_1821 & _GEN_2428 | (_GEN_1372 ? io_enq_uops_2_exception : rob_exception_2_12));
    rob_exception_2_11 <= ~_GEN_2623 & (_GEN_1821 & _GEN_2427 | (_GEN_1371 ? io_enq_uops_2_exception : rob_exception_2_11));
    rob_exception_2_10 <= ~_GEN_2622 & (_GEN_1821 & _GEN_2426 | (_GEN_1370 ? io_enq_uops_2_exception : rob_exception_2_10));
    rob_exception_2_9 <= ~_GEN_2621 & (_GEN_1821 & _GEN_2425 | (_GEN_1369 ? io_enq_uops_2_exception : rob_exception_2_9));
    rob_exception_2_8 <= ~_GEN_2620 & (_GEN_1821 & _GEN_2424 | (_GEN_1368 ? io_enq_uops_2_exception : rob_exception_2_8));
    rob_exception_2_7 <= ~_GEN_2619 & (_GEN_1821 & _GEN_2423 | (_GEN_1367 ? io_enq_uops_2_exception : rob_exception_2_7));
    rob_exception_2_6 <= ~_GEN_2618 & (_GEN_1821 & _GEN_2422 | (_GEN_1366 ? io_enq_uops_2_exception : rob_exception_2_6));
    rob_exception_2_5 <= ~_GEN_2617 & (_GEN_1821 & _GEN_2421 | (_GEN_1365 ? io_enq_uops_2_exception : rob_exception_2_5));
    rob_exception_2_4 <= ~_GEN_2616 & (_GEN_1821 & _GEN_2420 | (_GEN_1364 ? io_enq_uops_2_exception : rob_exception_2_4));
    rob_exception_2_3 <= ~_GEN_2615 & (_GEN_1821 & _GEN_2419 | (_GEN_1363 ? io_enq_uops_2_exception : rob_exception_2_3));
    rob_exception_2_2 <= ~_GEN_2614 & (_GEN_1821 & _GEN_2418 | (_GEN_1362 ? io_enq_uops_2_exception : rob_exception_2_2));
    rob_exception_2_1 <= ~_GEN_2613 & (_GEN_1821 & _GEN_2417 | (_GEN_1361 ? io_enq_uops_2_exception : rob_exception_2_1));
    rob_exception_2_0 <= ~_GEN_2612 & (_GEN_1821 & _GEN_2416 | (_GEN_1360 ? io_enq_uops_2_exception : rob_exception_2_0));
    rob_bsy_3_31 <= ~_GEN_2282 & (_GEN_2217 ? ~_GEN_2249 & _GEN_47495 : ~_GEN_2216 & _GEN_47495);
    rob_bsy_3_30 <= ~_GEN_2281 & (_GEN_2217 ? ~_GEN_2248 & _GEN_47494 : ~_GEN_2215 & _GEN_47494);
    rob_bsy_3_29 <= ~_GEN_2280 & (_GEN_2217 ? ~_GEN_2247 & _GEN_47493 : ~_GEN_2214 & _GEN_47493);
    rob_bsy_3_28 <= ~_GEN_2279 & (_GEN_2217 ? ~_GEN_2246 & _GEN_47492 : ~_GEN_2213 & _GEN_47492);
    rob_bsy_3_27 <= ~_GEN_2278 & (_GEN_2217 ? ~_GEN_2245 & _GEN_47491 : ~_GEN_2212 & _GEN_47491);
    rob_bsy_3_26 <= ~_GEN_2277 & (_GEN_2217 ? ~_GEN_2244 & _GEN_47490 : ~_GEN_2211 & _GEN_47490);
    rob_bsy_3_25 <= ~_GEN_2276 & (_GEN_2217 ? ~_GEN_2243 & _GEN_47489 : ~_GEN_2210 & _GEN_47489);
    rob_bsy_3_24 <= ~_GEN_2275 & (_GEN_2217 ? ~_GEN_2242 & _GEN_47488 : ~_GEN_2209 & _GEN_47488);
    rob_bsy_3_23 <= ~_GEN_2274 & (_GEN_2217 ? ~_GEN_2241 & _GEN_47487 : ~_GEN_2208 & _GEN_47487);
    rob_bsy_3_22 <= ~_GEN_2273 & (_GEN_2217 ? ~_GEN_2240 & _GEN_47486 : ~_GEN_2207 & _GEN_47486);
    rob_bsy_3_21 <= ~_GEN_2272 & (_GEN_2217 ? ~_GEN_2239 & _GEN_47485 : ~_GEN_2206 & _GEN_47485);
    rob_bsy_3_20 <= ~_GEN_2271 & (_GEN_2217 ? ~_GEN_2238 & _GEN_47484 : ~_GEN_2205 & _GEN_47484);
    rob_bsy_3_19 <= ~_GEN_2270 & (_GEN_2217 ? ~_GEN_2237 & _GEN_47483 : ~_GEN_2204 & _GEN_47483);
    rob_bsy_3_18 <= ~_GEN_2269 & (_GEN_2217 ? ~_GEN_2236 & _GEN_47482 : ~_GEN_2203 & _GEN_47482);
    rob_bsy_3_17 <= ~_GEN_2268 & (_GEN_2217 ? ~_GEN_2235 & _GEN_47481 : ~_GEN_2202 & _GEN_47481);
    rob_bsy_3_16 <= ~_GEN_2267 & (_GEN_2217 ? ~_GEN_2234 & _GEN_47480 : ~_GEN_2201 & _GEN_47480);
    rob_bsy_3_15 <= ~_GEN_2266 & (_GEN_2217 ? ~_GEN_2233 & _GEN_47479 : ~_GEN_2200 & _GEN_47479);
    rob_bsy_3_14 <= ~_GEN_2265 & (_GEN_2217 ? ~_GEN_2232 & _GEN_47478 : ~_GEN_2199 & _GEN_47478);
    rob_bsy_3_13 <= ~_GEN_2264 & (_GEN_2217 ? ~_GEN_2231 & _GEN_47477 : ~_GEN_2198 & _GEN_47477);
    rob_bsy_3_12 <= ~_GEN_2263 & (_GEN_2217 ? ~_GEN_2230 & _GEN_47476 : ~_GEN_2197 & _GEN_47476);
    rob_bsy_3_11 <= ~_GEN_2262 & (_GEN_2217 ? ~_GEN_2229 & _GEN_47475 : ~_GEN_2196 & _GEN_47475);
    rob_bsy_3_10 <= ~_GEN_2261 & (_GEN_2217 ? ~_GEN_2228 & _GEN_47474 : ~_GEN_2195 & _GEN_47474);
    rob_bsy_3_9 <= ~_GEN_2260 & (_GEN_2217 ? ~_GEN_2227 & _GEN_47473 : ~_GEN_2194 & _GEN_47473);
    rob_bsy_3_8 <= ~_GEN_2259 & (_GEN_2217 ? ~_GEN_2226 & _GEN_47472 : ~_GEN_2193 & _GEN_47472);
    rob_bsy_3_7 <= ~_GEN_2258 & (_GEN_2217 ? ~_GEN_2225 & _GEN_47471 : ~_GEN_2192 & _GEN_47471);
    rob_bsy_3_6 <= ~_GEN_2257 & (_GEN_2217 ? ~_GEN_2224 & _GEN_47470 : ~_GEN_2191 & _GEN_47470);
    rob_bsy_3_5 <= ~_GEN_2256 & (_GEN_2217 ? ~_GEN_2223 & _GEN_47469 : ~_GEN_2190 & _GEN_47469);
    rob_bsy_3_4 <= ~_GEN_2255 & (_GEN_2217 ? ~_GEN_2222 & _GEN_47468 : ~_GEN_2189 & _GEN_47468);
    rob_bsy_3_3 <= ~_GEN_2254 & (_GEN_2217 ? ~_GEN_2221 & _GEN_47467 : ~_GEN_2188 & _GEN_47467);
    rob_bsy_3_2 <= ~_GEN_2253 & (_GEN_2217 ? ~_GEN_2220 & _GEN_47466 : ~_GEN_2187 & _GEN_47466);
    rob_bsy_3_1 <= ~_GEN_2252 & (_GEN_2217 ? ~_GEN_2219 & _GEN_47465 : ~_GEN_2186 & _GEN_47465);
    rob_bsy_3_0 <= ~_GEN_2251 & (_GEN_2217 ? ~_GEN_2218 & _GEN_47464 : ~_GEN_2185 & _GEN_47464);
    rob_exception_3_31 <= ~_GEN_2710 & (_GEN_2283 & (&(io_lxcpt_bits_uop_rob_idx[6:2])) | (_GEN_1853 ? io_enq_uops_3_exception : rob_exception_3_31));
    rob_exception_3_30 <= ~_GEN_2709 & (_GEN_2283 & _GEN_2446 | (_GEN_1852 ? io_enq_uops_3_exception : rob_exception_3_30));
    rob_exception_3_29 <= ~_GEN_2708 & (_GEN_2283 & _GEN_2445 | (_GEN_1851 ? io_enq_uops_3_exception : rob_exception_3_29));
    rob_exception_3_28 <= ~_GEN_2707 & (_GEN_2283 & _GEN_2444 | (_GEN_1850 ? io_enq_uops_3_exception : rob_exception_3_28));
    rob_exception_3_27 <= ~_GEN_2706 & (_GEN_2283 & _GEN_2443 | (_GEN_1849 ? io_enq_uops_3_exception : rob_exception_3_27));
    rob_exception_3_26 <= ~_GEN_2705 & (_GEN_2283 & _GEN_2442 | (_GEN_1848 ? io_enq_uops_3_exception : rob_exception_3_26));
    rob_exception_3_25 <= ~_GEN_2704 & (_GEN_2283 & _GEN_2441 | (_GEN_1847 ? io_enq_uops_3_exception : rob_exception_3_25));
    rob_exception_3_24 <= ~_GEN_2703 & (_GEN_2283 & _GEN_2440 | (_GEN_1846 ? io_enq_uops_3_exception : rob_exception_3_24));
    rob_exception_3_23 <= ~_GEN_2702 & (_GEN_2283 & _GEN_2439 | (_GEN_1845 ? io_enq_uops_3_exception : rob_exception_3_23));
    rob_exception_3_22 <= ~_GEN_2701 & (_GEN_2283 & _GEN_2438 | (_GEN_1844 ? io_enq_uops_3_exception : rob_exception_3_22));
    rob_exception_3_21 <= ~_GEN_2700 & (_GEN_2283 & _GEN_2437 | (_GEN_1843 ? io_enq_uops_3_exception : rob_exception_3_21));
    rob_exception_3_20 <= ~_GEN_2699 & (_GEN_2283 & _GEN_2436 | (_GEN_1842 ? io_enq_uops_3_exception : rob_exception_3_20));
    rob_exception_3_19 <= ~_GEN_2698 & (_GEN_2283 & _GEN_2435 | (_GEN_1841 ? io_enq_uops_3_exception : rob_exception_3_19));
    rob_exception_3_18 <= ~_GEN_2697 & (_GEN_2283 & _GEN_2434 | (_GEN_1840 ? io_enq_uops_3_exception : rob_exception_3_18));
    rob_exception_3_17 <= ~_GEN_2696 & (_GEN_2283 & _GEN_2433 | (_GEN_1839 ? io_enq_uops_3_exception : rob_exception_3_17));
    rob_exception_3_16 <= ~_GEN_2695 & (_GEN_2283 & _GEN_2432 | (_GEN_1838 ? io_enq_uops_3_exception : rob_exception_3_16));
    rob_exception_3_15 <= ~_GEN_2694 & (_GEN_2283 & _GEN_2431 | (_GEN_1837 ? io_enq_uops_3_exception : rob_exception_3_15));
    rob_exception_3_14 <= ~_GEN_2693 & (_GEN_2283 & _GEN_2430 | (_GEN_1836 ? io_enq_uops_3_exception : rob_exception_3_14));
    rob_exception_3_13 <= ~_GEN_2692 & (_GEN_2283 & _GEN_2429 | (_GEN_1835 ? io_enq_uops_3_exception : rob_exception_3_13));
    rob_exception_3_12 <= ~_GEN_2691 & (_GEN_2283 & _GEN_2428 | (_GEN_1834 ? io_enq_uops_3_exception : rob_exception_3_12));
    rob_exception_3_11 <= ~_GEN_2690 & (_GEN_2283 & _GEN_2427 | (_GEN_1833 ? io_enq_uops_3_exception : rob_exception_3_11));
    rob_exception_3_10 <= ~_GEN_2689 & (_GEN_2283 & _GEN_2426 | (_GEN_1832 ? io_enq_uops_3_exception : rob_exception_3_10));
    rob_exception_3_9 <= ~_GEN_2688 & (_GEN_2283 & _GEN_2425 | (_GEN_1831 ? io_enq_uops_3_exception : rob_exception_3_9));
    rob_exception_3_8 <= ~_GEN_2687 & (_GEN_2283 & _GEN_2424 | (_GEN_1830 ? io_enq_uops_3_exception : rob_exception_3_8));
    rob_exception_3_7 <= ~_GEN_2686 & (_GEN_2283 & _GEN_2423 | (_GEN_1829 ? io_enq_uops_3_exception : rob_exception_3_7));
    rob_exception_3_6 <= ~_GEN_2685 & (_GEN_2283 & _GEN_2422 | (_GEN_1828 ? io_enq_uops_3_exception : rob_exception_3_6));
    rob_exception_3_5 <= ~_GEN_2684 & (_GEN_2283 & _GEN_2421 | (_GEN_1827 ? io_enq_uops_3_exception : rob_exception_3_5));
    rob_exception_3_4 <= ~_GEN_2683 & (_GEN_2283 & _GEN_2420 | (_GEN_1826 ? io_enq_uops_3_exception : rob_exception_3_4));
    rob_exception_3_3 <= ~_GEN_2682 & (_GEN_2283 & _GEN_2419 | (_GEN_1825 ? io_enq_uops_3_exception : rob_exception_3_3));
    rob_exception_3_2 <= ~_GEN_2681 & (_GEN_2283 & _GEN_2418 | (_GEN_1824 ? io_enq_uops_3_exception : rob_exception_3_2));
    rob_exception_3_1 <= ~_GEN_2680 & (_GEN_2283 & _GEN_2417 | (_GEN_1823 ? io_enq_uops_3_exception : rob_exception_3_1));
    rob_exception_3_0 <= ~_GEN_2679 & (_GEN_2283 & _GEN_2416 | (_GEN_1822 ? io_enq_uops_3_exception : rob_exception_3_0));
    if (_GEN_2384 & _GEN_2385)
      rob_fflags_0_0 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2353)
      rob_fflags_0_0 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2321)
      rob_fflags_0_0 <= io_fflags_0_bits_flags;
    else if (_GEN_33)
      rob_fflags_0_0 <= 5'h0;
    if (_GEN_2384 & _GEN_2386)
      rob_fflags_0_1 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2354)
      rob_fflags_0_1 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2322)
      rob_fflags_0_1 <= io_fflags_0_bits_flags;
    else if (_GEN_34)
      rob_fflags_0_1 <= 5'h0;
    if (_GEN_2384 & _GEN_2387)
      rob_fflags_0_2 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2355)
      rob_fflags_0_2 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2323)
      rob_fflags_0_2 <= io_fflags_0_bits_flags;
    else if (_GEN_35)
      rob_fflags_0_2 <= 5'h0;
    if (_GEN_2384 & _GEN_2388)
      rob_fflags_0_3 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2356)
      rob_fflags_0_3 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2324)
      rob_fflags_0_3 <= io_fflags_0_bits_flags;
    else if (_GEN_36)
      rob_fflags_0_3 <= 5'h0;
    if (_GEN_2384 & _GEN_2389)
      rob_fflags_0_4 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2357)
      rob_fflags_0_4 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2325)
      rob_fflags_0_4 <= io_fflags_0_bits_flags;
    else if (_GEN_37)
      rob_fflags_0_4 <= 5'h0;
    if (_GEN_2384 & _GEN_2390)
      rob_fflags_0_5 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2358)
      rob_fflags_0_5 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2326)
      rob_fflags_0_5 <= io_fflags_0_bits_flags;
    else if (_GEN_38)
      rob_fflags_0_5 <= 5'h0;
    if (_GEN_2384 & _GEN_2391)
      rob_fflags_0_6 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2359)
      rob_fflags_0_6 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2327)
      rob_fflags_0_6 <= io_fflags_0_bits_flags;
    else if (_GEN_39)
      rob_fflags_0_6 <= 5'h0;
    if (_GEN_2384 & _GEN_2392)
      rob_fflags_0_7 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2360)
      rob_fflags_0_7 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2328)
      rob_fflags_0_7 <= io_fflags_0_bits_flags;
    else if (_GEN_40)
      rob_fflags_0_7 <= 5'h0;
    if (_GEN_2384 & _GEN_2393)
      rob_fflags_0_8 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2361)
      rob_fflags_0_8 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2329)
      rob_fflags_0_8 <= io_fflags_0_bits_flags;
    else if (_GEN_41)
      rob_fflags_0_8 <= 5'h0;
    if (_GEN_2384 & _GEN_2394)
      rob_fflags_0_9 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2362)
      rob_fflags_0_9 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2330)
      rob_fflags_0_9 <= io_fflags_0_bits_flags;
    else if (_GEN_42)
      rob_fflags_0_9 <= 5'h0;
    if (_GEN_2384 & _GEN_2395)
      rob_fflags_0_10 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2363)
      rob_fflags_0_10 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2331)
      rob_fflags_0_10 <= io_fflags_0_bits_flags;
    else if (_GEN_43)
      rob_fflags_0_10 <= 5'h0;
    if (_GEN_2384 & _GEN_2396)
      rob_fflags_0_11 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2364)
      rob_fflags_0_11 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2332)
      rob_fflags_0_11 <= io_fflags_0_bits_flags;
    else if (_GEN_44)
      rob_fflags_0_11 <= 5'h0;
    if (_GEN_2384 & _GEN_2397)
      rob_fflags_0_12 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2365)
      rob_fflags_0_12 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2333)
      rob_fflags_0_12 <= io_fflags_0_bits_flags;
    else if (_GEN_45)
      rob_fflags_0_12 <= 5'h0;
    if (_GEN_2384 & _GEN_2398)
      rob_fflags_0_13 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2366)
      rob_fflags_0_13 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2334)
      rob_fflags_0_13 <= io_fflags_0_bits_flags;
    else if (_GEN_46)
      rob_fflags_0_13 <= 5'h0;
    if (_GEN_2384 & _GEN_2399)
      rob_fflags_0_14 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2367)
      rob_fflags_0_14 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2335)
      rob_fflags_0_14 <= io_fflags_0_bits_flags;
    else if (_GEN_47)
      rob_fflags_0_14 <= 5'h0;
    if (_GEN_2384 & _GEN_2400)
      rob_fflags_0_15 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2368)
      rob_fflags_0_15 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2336)
      rob_fflags_0_15 <= io_fflags_0_bits_flags;
    else if (_GEN_48)
      rob_fflags_0_15 <= 5'h0;
    if (_GEN_2384 & _GEN_2401)
      rob_fflags_0_16 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2369)
      rob_fflags_0_16 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2337)
      rob_fflags_0_16 <= io_fflags_0_bits_flags;
    else if (_GEN_49)
      rob_fflags_0_16 <= 5'h0;
    if (_GEN_2384 & _GEN_2402)
      rob_fflags_0_17 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2370)
      rob_fflags_0_17 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2338)
      rob_fflags_0_17 <= io_fflags_0_bits_flags;
    else if (_GEN_50)
      rob_fflags_0_17 <= 5'h0;
    if (_GEN_2384 & _GEN_2403)
      rob_fflags_0_18 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2371)
      rob_fflags_0_18 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2339)
      rob_fflags_0_18 <= io_fflags_0_bits_flags;
    else if (_GEN_51)
      rob_fflags_0_18 <= 5'h0;
    if (_GEN_2384 & _GEN_2404)
      rob_fflags_0_19 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2372)
      rob_fflags_0_19 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2340)
      rob_fflags_0_19 <= io_fflags_0_bits_flags;
    else if (_GEN_52)
      rob_fflags_0_19 <= 5'h0;
    if (_GEN_2384 & _GEN_2405)
      rob_fflags_0_20 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2373)
      rob_fflags_0_20 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2341)
      rob_fflags_0_20 <= io_fflags_0_bits_flags;
    else if (_GEN_53)
      rob_fflags_0_20 <= 5'h0;
    if (_GEN_2384 & _GEN_2406)
      rob_fflags_0_21 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2374)
      rob_fflags_0_21 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2342)
      rob_fflags_0_21 <= io_fflags_0_bits_flags;
    else if (_GEN_54)
      rob_fflags_0_21 <= 5'h0;
    if (_GEN_2384 & _GEN_2407)
      rob_fflags_0_22 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2375)
      rob_fflags_0_22 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2343)
      rob_fflags_0_22 <= io_fflags_0_bits_flags;
    else if (_GEN_55)
      rob_fflags_0_22 <= 5'h0;
    if (_GEN_2384 & _GEN_2408)
      rob_fflags_0_23 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2376)
      rob_fflags_0_23 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2344)
      rob_fflags_0_23 <= io_fflags_0_bits_flags;
    else if (_GEN_56)
      rob_fflags_0_23 <= 5'h0;
    if (_GEN_2384 & _GEN_2409)
      rob_fflags_0_24 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2377)
      rob_fflags_0_24 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2345)
      rob_fflags_0_24 <= io_fflags_0_bits_flags;
    else if (_GEN_57)
      rob_fflags_0_24 <= 5'h0;
    if (_GEN_2384 & _GEN_2410)
      rob_fflags_0_25 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2378)
      rob_fflags_0_25 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2346)
      rob_fflags_0_25 <= io_fflags_0_bits_flags;
    else if (_GEN_58)
      rob_fflags_0_25 <= 5'h0;
    if (_GEN_2384 & _GEN_2411)
      rob_fflags_0_26 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2379)
      rob_fflags_0_26 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2347)
      rob_fflags_0_26 <= io_fflags_0_bits_flags;
    else if (_GEN_59)
      rob_fflags_0_26 <= 5'h0;
    if (_GEN_2384 & _GEN_2412)
      rob_fflags_0_27 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2380)
      rob_fflags_0_27 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2348)
      rob_fflags_0_27 <= io_fflags_0_bits_flags;
    else if (_GEN_60)
      rob_fflags_0_27 <= 5'h0;
    if (_GEN_2384 & _GEN_2413)
      rob_fflags_0_28 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2381)
      rob_fflags_0_28 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2349)
      rob_fflags_0_28 <= io_fflags_0_bits_flags;
    else if (_GEN_61)
      rob_fflags_0_28 <= 5'h0;
    if (_GEN_2384 & _GEN_2414)
      rob_fflags_0_29 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2382)
      rob_fflags_0_29 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2350)
      rob_fflags_0_29 <= io_fflags_0_bits_flags;
    else if (_GEN_62)
      rob_fflags_0_29 <= 5'h0;
    if (_GEN_2384 & _GEN_2415)
      rob_fflags_0_30 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & _GEN_2383)
      rob_fflags_0_30 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & _GEN_2351)
      rob_fflags_0_30 <= io_fflags_0_bits_flags;
    else if (_GEN_63)
      rob_fflags_0_30 <= 5'h0;
    if (_GEN_2384 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_0_31 <= io_fflags_3_bits_flags;
    else if (_GEN_2352 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_0_31 <= io_fflags_2_bits_flags;
    else if (_GEN_2320 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_0_31 <= io_fflags_0_bits_flags;
    else if (_GEN_64)
      rob_fflags_0_31 <= 5'h0;
    if (_GEN_2544 & _GEN_2385)
      rob_fflags_1_0 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2353)
      rob_fflags_1_0 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2321)
      rob_fflags_1_0 <= io_fflags_0_bits_flags;
    else if (_GEN_898)
      rob_fflags_1_0 <= 5'h0;
    if (_GEN_2544 & _GEN_2386)
      rob_fflags_1_1 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2354)
      rob_fflags_1_1 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2322)
      rob_fflags_1_1 <= io_fflags_0_bits_flags;
    else if (_GEN_899)
      rob_fflags_1_1 <= 5'h0;
    if (_GEN_2544 & _GEN_2387)
      rob_fflags_1_2 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2355)
      rob_fflags_1_2 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2323)
      rob_fflags_1_2 <= io_fflags_0_bits_flags;
    else if (_GEN_900)
      rob_fflags_1_2 <= 5'h0;
    if (_GEN_2544 & _GEN_2388)
      rob_fflags_1_3 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2356)
      rob_fflags_1_3 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2324)
      rob_fflags_1_3 <= io_fflags_0_bits_flags;
    else if (_GEN_901)
      rob_fflags_1_3 <= 5'h0;
    if (_GEN_2544 & _GEN_2389)
      rob_fflags_1_4 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2357)
      rob_fflags_1_4 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2325)
      rob_fflags_1_4 <= io_fflags_0_bits_flags;
    else if (_GEN_902)
      rob_fflags_1_4 <= 5'h0;
    if (_GEN_2544 & _GEN_2390)
      rob_fflags_1_5 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2358)
      rob_fflags_1_5 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2326)
      rob_fflags_1_5 <= io_fflags_0_bits_flags;
    else if (_GEN_903)
      rob_fflags_1_5 <= 5'h0;
    if (_GEN_2544 & _GEN_2391)
      rob_fflags_1_6 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2359)
      rob_fflags_1_6 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2327)
      rob_fflags_1_6 <= io_fflags_0_bits_flags;
    else if (_GEN_904)
      rob_fflags_1_6 <= 5'h0;
    if (_GEN_2544 & _GEN_2392)
      rob_fflags_1_7 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2360)
      rob_fflags_1_7 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2328)
      rob_fflags_1_7 <= io_fflags_0_bits_flags;
    else if (_GEN_905)
      rob_fflags_1_7 <= 5'h0;
    if (_GEN_2544 & _GEN_2393)
      rob_fflags_1_8 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2361)
      rob_fflags_1_8 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2329)
      rob_fflags_1_8 <= io_fflags_0_bits_flags;
    else if (_GEN_906)
      rob_fflags_1_8 <= 5'h0;
    if (_GEN_2544 & _GEN_2394)
      rob_fflags_1_9 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2362)
      rob_fflags_1_9 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2330)
      rob_fflags_1_9 <= io_fflags_0_bits_flags;
    else if (_GEN_907)
      rob_fflags_1_9 <= 5'h0;
    if (_GEN_2544 & _GEN_2395)
      rob_fflags_1_10 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2363)
      rob_fflags_1_10 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2331)
      rob_fflags_1_10 <= io_fflags_0_bits_flags;
    else if (_GEN_908)
      rob_fflags_1_10 <= 5'h0;
    if (_GEN_2544 & _GEN_2396)
      rob_fflags_1_11 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2364)
      rob_fflags_1_11 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2332)
      rob_fflags_1_11 <= io_fflags_0_bits_flags;
    else if (_GEN_909)
      rob_fflags_1_11 <= 5'h0;
    if (_GEN_2544 & _GEN_2397)
      rob_fflags_1_12 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2365)
      rob_fflags_1_12 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2333)
      rob_fflags_1_12 <= io_fflags_0_bits_flags;
    else if (_GEN_910)
      rob_fflags_1_12 <= 5'h0;
    if (_GEN_2544 & _GEN_2398)
      rob_fflags_1_13 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2366)
      rob_fflags_1_13 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2334)
      rob_fflags_1_13 <= io_fflags_0_bits_flags;
    else if (_GEN_911)
      rob_fflags_1_13 <= 5'h0;
    if (_GEN_2544 & _GEN_2399)
      rob_fflags_1_14 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2367)
      rob_fflags_1_14 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2335)
      rob_fflags_1_14 <= io_fflags_0_bits_flags;
    else if (_GEN_912)
      rob_fflags_1_14 <= 5'h0;
    if (_GEN_2544 & _GEN_2400)
      rob_fflags_1_15 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2368)
      rob_fflags_1_15 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2336)
      rob_fflags_1_15 <= io_fflags_0_bits_flags;
    else if (_GEN_913)
      rob_fflags_1_15 <= 5'h0;
    if (_GEN_2544 & _GEN_2401)
      rob_fflags_1_16 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2369)
      rob_fflags_1_16 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2337)
      rob_fflags_1_16 <= io_fflags_0_bits_flags;
    else if (_GEN_914)
      rob_fflags_1_16 <= 5'h0;
    if (_GEN_2544 & _GEN_2402)
      rob_fflags_1_17 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2370)
      rob_fflags_1_17 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2338)
      rob_fflags_1_17 <= io_fflags_0_bits_flags;
    else if (_GEN_915)
      rob_fflags_1_17 <= 5'h0;
    if (_GEN_2544 & _GEN_2403)
      rob_fflags_1_18 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2371)
      rob_fflags_1_18 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2339)
      rob_fflags_1_18 <= io_fflags_0_bits_flags;
    else if (_GEN_916)
      rob_fflags_1_18 <= 5'h0;
    if (_GEN_2544 & _GEN_2404)
      rob_fflags_1_19 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2372)
      rob_fflags_1_19 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2340)
      rob_fflags_1_19 <= io_fflags_0_bits_flags;
    else if (_GEN_917)
      rob_fflags_1_19 <= 5'h0;
    if (_GEN_2544 & _GEN_2405)
      rob_fflags_1_20 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2373)
      rob_fflags_1_20 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2341)
      rob_fflags_1_20 <= io_fflags_0_bits_flags;
    else if (_GEN_918)
      rob_fflags_1_20 <= 5'h0;
    if (_GEN_2544 & _GEN_2406)
      rob_fflags_1_21 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2374)
      rob_fflags_1_21 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2342)
      rob_fflags_1_21 <= io_fflags_0_bits_flags;
    else if (_GEN_919)
      rob_fflags_1_21 <= 5'h0;
    if (_GEN_2544 & _GEN_2407)
      rob_fflags_1_22 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2375)
      rob_fflags_1_22 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2343)
      rob_fflags_1_22 <= io_fflags_0_bits_flags;
    else if (_GEN_920)
      rob_fflags_1_22 <= 5'h0;
    if (_GEN_2544 & _GEN_2408)
      rob_fflags_1_23 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2376)
      rob_fflags_1_23 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2344)
      rob_fflags_1_23 <= io_fflags_0_bits_flags;
    else if (_GEN_921)
      rob_fflags_1_23 <= 5'h0;
    if (_GEN_2544 & _GEN_2409)
      rob_fflags_1_24 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2377)
      rob_fflags_1_24 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2345)
      rob_fflags_1_24 <= io_fflags_0_bits_flags;
    else if (_GEN_922)
      rob_fflags_1_24 <= 5'h0;
    if (_GEN_2544 & _GEN_2410)
      rob_fflags_1_25 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2378)
      rob_fflags_1_25 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2346)
      rob_fflags_1_25 <= io_fflags_0_bits_flags;
    else if (_GEN_923)
      rob_fflags_1_25 <= 5'h0;
    if (_GEN_2544 & _GEN_2411)
      rob_fflags_1_26 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2379)
      rob_fflags_1_26 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2347)
      rob_fflags_1_26 <= io_fflags_0_bits_flags;
    else if (_GEN_924)
      rob_fflags_1_26 <= 5'h0;
    if (_GEN_2544 & _GEN_2412)
      rob_fflags_1_27 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2380)
      rob_fflags_1_27 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2348)
      rob_fflags_1_27 <= io_fflags_0_bits_flags;
    else if (_GEN_925)
      rob_fflags_1_27 <= 5'h0;
    if (_GEN_2544 & _GEN_2413)
      rob_fflags_1_28 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2381)
      rob_fflags_1_28 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2349)
      rob_fflags_1_28 <= io_fflags_0_bits_flags;
    else if (_GEN_926)
      rob_fflags_1_28 <= 5'h0;
    if (_GEN_2544 & _GEN_2414)
      rob_fflags_1_29 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2382)
      rob_fflags_1_29 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2350)
      rob_fflags_1_29 <= io_fflags_0_bits_flags;
    else if (_GEN_927)
      rob_fflags_1_29 <= 5'h0;
    if (_GEN_2544 & _GEN_2415)
      rob_fflags_1_30 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & _GEN_2383)
      rob_fflags_1_30 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & _GEN_2351)
      rob_fflags_1_30 <= io_fflags_0_bits_flags;
    else if (_GEN_928)
      rob_fflags_1_30 <= 5'h0;
    if (_GEN_2544 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_1_31 <= io_fflags_3_bits_flags;
    else if (_GEN_2543 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_1_31 <= io_fflags_2_bits_flags;
    else if (_GEN_2542 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_1_31 <= io_fflags_0_bits_flags;
    else if (_GEN_929)
      rob_fflags_1_31 <= 5'h0;
    if (_GEN_2611 & _GEN_2385)
      rob_fflags_2_0 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2353)
      rob_fflags_2_0 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2321)
      rob_fflags_2_0 <= io_fflags_0_bits_flags;
    else if (_GEN_1360)
      rob_fflags_2_0 <= 5'h0;
    if (_GEN_2611 & _GEN_2386)
      rob_fflags_2_1 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2354)
      rob_fflags_2_1 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2322)
      rob_fflags_2_1 <= io_fflags_0_bits_flags;
    else if (_GEN_1361)
      rob_fflags_2_1 <= 5'h0;
    if (_GEN_2611 & _GEN_2387)
      rob_fflags_2_2 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2355)
      rob_fflags_2_2 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2323)
      rob_fflags_2_2 <= io_fflags_0_bits_flags;
    else if (_GEN_1362)
      rob_fflags_2_2 <= 5'h0;
    if (_GEN_2611 & _GEN_2388)
      rob_fflags_2_3 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2356)
      rob_fflags_2_3 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2324)
      rob_fflags_2_3 <= io_fflags_0_bits_flags;
    else if (_GEN_1363)
      rob_fflags_2_3 <= 5'h0;
    if (_GEN_2611 & _GEN_2389)
      rob_fflags_2_4 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2357)
      rob_fflags_2_4 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2325)
      rob_fflags_2_4 <= io_fflags_0_bits_flags;
    else if (_GEN_1364)
      rob_fflags_2_4 <= 5'h0;
    if (_GEN_2611 & _GEN_2390)
      rob_fflags_2_5 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2358)
      rob_fflags_2_5 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2326)
      rob_fflags_2_5 <= io_fflags_0_bits_flags;
    else if (_GEN_1365)
      rob_fflags_2_5 <= 5'h0;
    if (_GEN_2611 & _GEN_2391)
      rob_fflags_2_6 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2359)
      rob_fflags_2_6 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2327)
      rob_fflags_2_6 <= io_fflags_0_bits_flags;
    else if (_GEN_1366)
      rob_fflags_2_6 <= 5'h0;
    if (_GEN_2611 & _GEN_2392)
      rob_fflags_2_7 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2360)
      rob_fflags_2_7 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2328)
      rob_fflags_2_7 <= io_fflags_0_bits_flags;
    else if (_GEN_1367)
      rob_fflags_2_7 <= 5'h0;
    if (_GEN_2611 & _GEN_2393)
      rob_fflags_2_8 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2361)
      rob_fflags_2_8 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2329)
      rob_fflags_2_8 <= io_fflags_0_bits_flags;
    else if (_GEN_1368)
      rob_fflags_2_8 <= 5'h0;
    if (_GEN_2611 & _GEN_2394)
      rob_fflags_2_9 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2362)
      rob_fflags_2_9 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2330)
      rob_fflags_2_9 <= io_fflags_0_bits_flags;
    else if (_GEN_1369)
      rob_fflags_2_9 <= 5'h0;
    if (_GEN_2611 & _GEN_2395)
      rob_fflags_2_10 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2363)
      rob_fflags_2_10 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2331)
      rob_fflags_2_10 <= io_fflags_0_bits_flags;
    else if (_GEN_1370)
      rob_fflags_2_10 <= 5'h0;
    if (_GEN_2611 & _GEN_2396)
      rob_fflags_2_11 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2364)
      rob_fflags_2_11 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2332)
      rob_fflags_2_11 <= io_fflags_0_bits_flags;
    else if (_GEN_1371)
      rob_fflags_2_11 <= 5'h0;
    if (_GEN_2611 & _GEN_2397)
      rob_fflags_2_12 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2365)
      rob_fflags_2_12 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2333)
      rob_fflags_2_12 <= io_fflags_0_bits_flags;
    else if (_GEN_1372)
      rob_fflags_2_12 <= 5'h0;
    if (_GEN_2611 & _GEN_2398)
      rob_fflags_2_13 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2366)
      rob_fflags_2_13 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2334)
      rob_fflags_2_13 <= io_fflags_0_bits_flags;
    else if (_GEN_1373)
      rob_fflags_2_13 <= 5'h0;
    if (_GEN_2611 & _GEN_2399)
      rob_fflags_2_14 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2367)
      rob_fflags_2_14 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2335)
      rob_fflags_2_14 <= io_fflags_0_bits_flags;
    else if (_GEN_1374)
      rob_fflags_2_14 <= 5'h0;
    if (_GEN_2611 & _GEN_2400)
      rob_fflags_2_15 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2368)
      rob_fflags_2_15 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2336)
      rob_fflags_2_15 <= io_fflags_0_bits_flags;
    else if (_GEN_1375)
      rob_fflags_2_15 <= 5'h0;
    if (_GEN_2611 & _GEN_2401)
      rob_fflags_2_16 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2369)
      rob_fflags_2_16 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2337)
      rob_fflags_2_16 <= io_fflags_0_bits_flags;
    else if (_GEN_1376)
      rob_fflags_2_16 <= 5'h0;
    if (_GEN_2611 & _GEN_2402)
      rob_fflags_2_17 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2370)
      rob_fflags_2_17 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2338)
      rob_fflags_2_17 <= io_fflags_0_bits_flags;
    else if (_GEN_1377)
      rob_fflags_2_17 <= 5'h0;
    if (_GEN_2611 & _GEN_2403)
      rob_fflags_2_18 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2371)
      rob_fflags_2_18 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2339)
      rob_fflags_2_18 <= io_fflags_0_bits_flags;
    else if (_GEN_1378)
      rob_fflags_2_18 <= 5'h0;
    if (_GEN_2611 & _GEN_2404)
      rob_fflags_2_19 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2372)
      rob_fflags_2_19 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2340)
      rob_fflags_2_19 <= io_fflags_0_bits_flags;
    else if (_GEN_1379)
      rob_fflags_2_19 <= 5'h0;
    if (_GEN_2611 & _GEN_2405)
      rob_fflags_2_20 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2373)
      rob_fflags_2_20 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2341)
      rob_fflags_2_20 <= io_fflags_0_bits_flags;
    else if (_GEN_1380)
      rob_fflags_2_20 <= 5'h0;
    if (_GEN_2611 & _GEN_2406)
      rob_fflags_2_21 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2374)
      rob_fflags_2_21 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2342)
      rob_fflags_2_21 <= io_fflags_0_bits_flags;
    else if (_GEN_1381)
      rob_fflags_2_21 <= 5'h0;
    if (_GEN_2611 & _GEN_2407)
      rob_fflags_2_22 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2375)
      rob_fflags_2_22 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2343)
      rob_fflags_2_22 <= io_fflags_0_bits_flags;
    else if (_GEN_1382)
      rob_fflags_2_22 <= 5'h0;
    if (_GEN_2611 & _GEN_2408)
      rob_fflags_2_23 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2376)
      rob_fflags_2_23 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2344)
      rob_fflags_2_23 <= io_fflags_0_bits_flags;
    else if (_GEN_1383)
      rob_fflags_2_23 <= 5'h0;
    if (_GEN_2611 & _GEN_2409)
      rob_fflags_2_24 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2377)
      rob_fflags_2_24 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2345)
      rob_fflags_2_24 <= io_fflags_0_bits_flags;
    else if (_GEN_1384)
      rob_fflags_2_24 <= 5'h0;
    if (_GEN_2611 & _GEN_2410)
      rob_fflags_2_25 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2378)
      rob_fflags_2_25 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2346)
      rob_fflags_2_25 <= io_fflags_0_bits_flags;
    else if (_GEN_1385)
      rob_fflags_2_25 <= 5'h0;
    if (_GEN_2611 & _GEN_2411)
      rob_fflags_2_26 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2379)
      rob_fflags_2_26 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2347)
      rob_fflags_2_26 <= io_fflags_0_bits_flags;
    else if (_GEN_1386)
      rob_fflags_2_26 <= 5'h0;
    if (_GEN_2611 & _GEN_2412)
      rob_fflags_2_27 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2380)
      rob_fflags_2_27 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2348)
      rob_fflags_2_27 <= io_fflags_0_bits_flags;
    else if (_GEN_1387)
      rob_fflags_2_27 <= 5'h0;
    if (_GEN_2611 & _GEN_2413)
      rob_fflags_2_28 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2381)
      rob_fflags_2_28 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2349)
      rob_fflags_2_28 <= io_fflags_0_bits_flags;
    else if (_GEN_1388)
      rob_fflags_2_28 <= 5'h0;
    if (_GEN_2611 & _GEN_2414)
      rob_fflags_2_29 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2382)
      rob_fflags_2_29 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2350)
      rob_fflags_2_29 <= io_fflags_0_bits_flags;
    else if (_GEN_1389)
      rob_fflags_2_29 <= 5'h0;
    if (_GEN_2611 & _GEN_2415)
      rob_fflags_2_30 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & _GEN_2383)
      rob_fflags_2_30 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & _GEN_2351)
      rob_fflags_2_30 <= io_fflags_0_bits_flags;
    else if (_GEN_1390)
      rob_fflags_2_30 <= 5'h0;
    if (_GEN_2611 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_2_31 <= io_fflags_3_bits_flags;
    else if (_GEN_2610 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_2_31 <= io_fflags_2_bits_flags;
    else if (_GEN_2609 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_2_31 <= io_fflags_0_bits_flags;
    else if (_GEN_1391)
      rob_fflags_2_31 <= 5'h0;
    if (_GEN_2678 & _GEN_2385)
      rob_fflags_3_0 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2353)
      rob_fflags_3_0 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2321)
      rob_fflags_3_0 <= io_fflags_0_bits_flags;
    else if (_GEN_1822)
      rob_fflags_3_0 <= 5'h0;
    if (_GEN_2678 & _GEN_2386)
      rob_fflags_3_1 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2354)
      rob_fflags_3_1 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2322)
      rob_fflags_3_1 <= io_fflags_0_bits_flags;
    else if (_GEN_1823)
      rob_fflags_3_1 <= 5'h0;
    if (_GEN_2678 & _GEN_2387)
      rob_fflags_3_2 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2355)
      rob_fflags_3_2 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2323)
      rob_fflags_3_2 <= io_fflags_0_bits_flags;
    else if (_GEN_1824)
      rob_fflags_3_2 <= 5'h0;
    if (_GEN_2678 & _GEN_2388)
      rob_fflags_3_3 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2356)
      rob_fflags_3_3 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2324)
      rob_fflags_3_3 <= io_fflags_0_bits_flags;
    else if (_GEN_1825)
      rob_fflags_3_3 <= 5'h0;
    if (_GEN_2678 & _GEN_2389)
      rob_fflags_3_4 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2357)
      rob_fflags_3_4 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2325)
      rob_fflags_3_4 <= io_fflags_0_bits_flags;
    else if (_GEN_1826)
      rob_fflags_3_4 <= 5'h0;
    if (_GEN_2678 & _GEN_2390)
      rob_fflags_3_5 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2358)
      rob_fflags_3_5 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2326)
      rob_fflags_3_5 <= io_fflags_0_bits_flags;
    else if (_GEN_1827)
      rob_fflags_3_5 <= 5'h0;
    if (_GEN_2678 & _GEN_2391)
      rob_fflags_3_6 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2359)
      rob_fflags_3_6 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2327)
      rob_fflags_3_6 <= io_fflags_0_bits_flags;
    else if (_GEN_1828)
      rob_fflags_3_6 <= 5'h0;
    if (_GEN_2678 & _GEN_2392)
      rob_fflags_3_7 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2360)
      rob_fflags_3_7 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2328)
      rob_fflags_3_7 <= io_fflags_0_bits_flags;
    else if (_GEN_1829)
      rob_fflags_3_7 <= 5'h0;
    if (_GEN_2678 & _GEN_2393)
      rob_fflags_3_8 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2361)
      rob_fflags_3_8 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2329)
      rob_fflags_3_8 <= io_fflags_0_bits_flags;
    else if (_GEN_1830)
      rob_fflags_3_8 <= 5'h0;
    if (_GEN_2678 & _GEN_2394)
      rob_fflags_3_9 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2362)
      rob_fflags_3_9 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2330)
      rob_fflags_3_9 <= io_fflags_0_bits_flags;
    else if (_GEN_1831)
      rob_fflags_3_9 <= 5'h0;
    if (_GEN_2678 & _GEN_2395)
      rob_fflags_3_10 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2363)
      rob_fflags_3_10 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2331)
      rob_fflags_3_10 <= io_fflags_0_bits_flags;
    else if (_GEN_1832)
      rob_fflags_3_10 <= 5'h0;
    if (_GEN_2678 & _GEN_2396)
      rob_fflags_3_11 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2364)
      rob_fflags_3_11 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2332)
      rob_fflags_3_11 <= io_fflags_0_bits_flags;
    else if (_GEN_1833)
      rob_fflags_3_11 <= 5'h0;
    if (_GEN_2678 & _GEN_2397)
      rob_fflags_3_12 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2365)
      rob_fflags_3_12 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2333)
      rob_fflags_3_12 <= io_fflags_0_bits_flags;
    else if (_GEN_1834)
      rob_fflags_3_12 <= 5'h0;
    if (_GEN_2678 & _GEN_2398)
      rob_fflags_3_13 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2366)
      rob_fflags_3_13 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2334)
      rob_fflags_3_13 <= io_fflags_0_bits_flags;
    else if (_GEN_1835)
      rob_fflags_3_13 <= 5'h0;
    if (_GEN_2678 & _GEN_2399)
      rob_fflags_3_14 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2367)
      rob_fflags_3_14 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2335)
      rob_fflags_3_14 <= io_fflags_0_bits_flags;
    else if (_GEN_1836)
      rob_fflags_3_14 <= 5'h0;
    if (_GEN_2678 & _GEN_2400)
      rob_fflags_3_15 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2368)
      rob_fflags_3_15 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2336)
      rob_fflags_3_15 <= io_fflags_0_bits_flags;
    else if (_GEN_1837)
      rob_fflags_3_15 <= 5'h0;
    if (_GEN_2678 & _GEN_2401)
      rob_fflags_3_16 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2369)
      rob_fflags_3_16 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2337)
      rob_fflags_3_16 <= io_fflags_0_bits_flags;
    else if (_GEN_1838)
      rob_fflags_3_16 <= 5'h0;
    if (_GEN_2678 & _GEN_2402)
      rob_fflags_3_17 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2370)
      rob_fflags_3_17 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2338)
      rob_fflags_3_17 <= io_fflags_0_bits_flags;
    else if (_GEN_1839)
      rob_fflags_3_17 <= 5'h0;
    if (_GEN_2678 & _GEN_2403)
      rob_fflags_3_18 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2371)
      rob_fflags_3_18 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2339)
      rob_fflags_3_18 <= io_fflags_0_bits_flags;
    else if (_GEN_1840)
      rob_fflags_3_18 <= 5'h0;
    if (_GEN_2678 & _GEN_2404)
      rob_fflags_3_19 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2372)
      rob_fflags_3_19 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2340)
      rob_fflags_3_19 <= io_fflags_0_bits_flags;
    else if (_GEN_1841)
      rob_fflags_3_19 <= 5'h0;
    if (_GEN_2678 & _GEN_2405)
      rob_fflags_3_20 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2373)
      rob_fflags_3_20 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2341)
      rob_fflags_3_20 <= io_fflags_0_bits_flags;
    else if (_GEN_1842)
      rob_fflags_3_20 <= 5'h0;
    if (_GEN_2678 & _GEN_2406)
      rob_fflags_3_21 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2374)
      rob_fflags_3_21 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2342)
      rob_fflags_3_21 <= io_fflags_0_bits_flags;
    else if (_GEN_1843)
      rob_fflags_3_21 <= 5'h0;
    if (_GEN_2678 & _GEN_2407)
      rob_fflags_3_22 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2375)
      rob_fflags_3_22 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2343)
      rob_fflags_3_22 <= io_fflags_0_bits_flags;
    else if (_GEN_1844)
      rob_fflags_3_22 <= 5'h0;
    if (_GEN_2678 & _GEN_2408)
      rob_fflags_3_23 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2376)
      rob_fflags_3_23 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2344)
      rob_fflags_3_23 <= io_fflags_0_bits_flags;
    else if (_GEN_1845)
      rob_fflags_3_23 <= 5'h0;
    if (_GEN_2678 & _GEN_2409)
      rob_fflags_3_24 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2377)
      rob_fflags_3_24 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2345)
      rob_fflags_3_24 <= io_fflags_0_bits_flags;
    else if (_GEN_1846)
      rob_fflags_3_24 <= 5'h0;
    if (_GEN_2678 & _GEN_2410)
      rob_fflags_3_25 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2378)
      rob_fflags_3_25 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2346)
      rob_fflags_3_25 <= io_fflags_0_bits_flags;
    else if (_GEN_1847)
      rob_fflags_3_25 <= 5'h0;
    if (_GEN_2678 & _GEN_2411)
      rob_fflags_3_26 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2379)
      rob_fflags_3_26 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2347)
      rob_fflags_3_26 <= io_fflags_0_bits_flags;
    else if (_GEN_1848)
      rob_fflags_3_26 <= 5'h0;
    if (_GEN_2678 & _GEN_2412)
      rob_fflags_3_27 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2380)
      rob_fflags_3_27 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2348)
      rob_fflags_3_27 <= io_fflags_0_bits_flags;
    else if (_GEN_1849)
      rob_fflags_3_27 <= 5'h0;
    if (_GEN_2678 & _GEN_2413)
      rob_fflags_3_28 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2381)
      rob_fflags_3_28 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2349)
      rob_fflags_3_28 <= io_fflags_0_bits_flags;
    else if (_GEN_1850)
      rob_fflags_3_28 <= 5'h0;
    if (_GEN_2678 & _GEN_2414)
      rob_fflags_3_29 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2382)
      rob_fflags_3_29 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2350)
      rob_fflags_3_29 <= io_fflags_0_bits_flags;
    else if (_GEN_1851)
      rob_fflags_3_29 <= 5'h0;
    if (_GEN_2678 & _GEN_2415)
      rob_fflags_3_30 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & _GEN_2383)
      rob_fflags_3_30 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & _GEN_2351)
      rob_fflags_3_30 <= io_fflags_0_bits_flags;
    else if (_GEN_1852)
      rob_fflags_3_30 <= 5'h0;
    if (_GEN_2678 & (&(io_fflags_3_bits_uop_rob_idx[6:2])))
      rob_fflags_3_31 <= io_fflags_3_bits_flags;
    else if (_GEN_2677 & (&(io_fflags_2_bits_uop_rob_idx[6:2])))
      rob_fflags_3_31 <= io_fflags_2_bits_flags;
    else if (_GEN_2676 & (&(io_fflags_0_bits_uop_rob_idx[6:2])))
      rob_fflags_3_31 <= io_fflags_0_bits_flags;
    else if (_GEN_1853)
      rob_fflags_3_31 <= 5'h0;
    if (_GEN_33) begin
      rob_uop__0_uopc <= io_enq_uops_0_uopc;
      rob_uop__0_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__0_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__0_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__0_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__0_pdst <= io_enq_uops_0_pdst;
      rob_uop__0_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__0_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__0_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__0_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__0_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__0_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__0_ldst <= io_enq_uops_0_ldst;
      rob_uop__0_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__0_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__0_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2510) | ~rob_val__0) begin
      if (_GEN_33)
        rob_uop__0_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__0_br_mask <= rob_uop__0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_34) begin
      rob_uop__1_uopc <= io_enq_uops_0_uopc;
      rob_uop__1_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__1_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__1_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__1_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__1_pdst <= io_enq_uops_0_pdst;
      rob_uop__1_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__1_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__1_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__1_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__1_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__1_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__1_ldst <= io_enq_uops_0_ldst;
      rob_uop__1_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__1_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__1_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2511) | ~rob_val__1) begin
      if (_GEN_34)
        rob_uop__1_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__1_br_mask <= rob_uop__1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_35) begin
      rob_uop__2_uopc <= io_enq_uops_0_uopc;
      rob_uop__2_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__2_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__2_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__2_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__2_pdst <= io_enq_uops_0_pdst;
      rob_uop__2_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__2_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__2_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__2_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__2_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__2_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__2_ldst <= io_enq_uops_0_ldst;
      rob_uop__2_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__2_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__2_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2512) | ~rob_val__2) begin
      if (_GEN_35)
        rob_uop__2_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__2_br_mask <= rob_uop__2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_36) begin
      rob_uop__3_uopc <= io_enq_uops_0_uopc;
      rob_uop__3_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__3_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__3_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__3_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__3_pdst <= io_enq_uops_0_pdst;
      rob_uop__3_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__3_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__3_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__3_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__3_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__3_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__3_ldst <= io_enq_uops_0_ldst;
      rob_uop__3_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__3_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__3_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2513) | ~rob_val__3) begin
      if (_GEN_36)
        rob_uop__3_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__3_br_mask <= rob_uop__3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_37) begin
      rob_uop__4_uopc <= io_enq_uops_0_uopc;
      rob_uop__4_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__4_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__4_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__4_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__4_pdst <= io_enq_uops_0_pdst;
      rob_uop__4_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__4_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__4_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__4_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__4_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__4_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__4_ldst <= io_enq_uops_0_ldst;
      rob_uop__4_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__4_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__4_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2514) | ~rob_val__4) begin
      if (_GEN_37)
        rob_uop__4_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__4_br_mask <= rob_uop__4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_38) begin
      rob_uop__5_uopc <= io_enq_uops_0_uopc;
      rob_uop__5_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__5_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__5_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__5_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__5_pdst <= io_enq_uops_0_pdst;
      rob_uop__5_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__5_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__5_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__5_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__5_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__5_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__5_ldst <= io_enq_uops_0_ldst;
      rob_uop__5_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__5_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__5_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2515) | ~rob_val__5) begin
      if (_GEN_38)
        rob_uop__5_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__5_br_mask <= rob_uop__5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_39) begin
      rob_uop__6_uopc <= io_enq_uops_0_uopc;
      rob_uop__6_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__6_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__6_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__6_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__6_pdst <= io_enq_uops_0_pdst;
      rob_uop__6_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__6_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__6_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__6_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__6_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__6_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__6_ldst <= io_enq_uops_0_ldst;
      rob_uop__6_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__6_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__6_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2516) | ~rob_val__6) begin
      if (_GEN_39)
        rob_uop__6_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__6_br_mask <= rob_uop__6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_40) begin
      rob_uop__7_uopc <= io_enq_uops_0_uopc;
      rob_uop__7_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__7_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__7_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__7_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__7_pdst <= io_enq_uops_0_pdst;
      rob_uop__7_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__7_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__7_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__7_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__7_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__7_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__7_ldst <= io_enq_uops_0_ldst;
      rob_uop__7_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__7_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__7_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2517) | ~rob_val__7) begin
      if (_GEN_40)
        rob_uop__7_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__7_br_mask <= rob_uop__7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_41) begin
      rob_uop__8_uopc <= io_enq_uops_0_uopc;
      rob_uop__8_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__8_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__8_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__8_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__8_pdst <= io_enq_uops_0_pdst;
      rob_uop__8_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__8_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__8_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__8_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__8_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__8_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__8_ldst <= io_enq_uops_0_ldst;
      rob_uop__8_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__8_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__8_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2518) | ~rob_val__8) begin
      if (_GEN_41)
        rob_uop__8_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__8_br_mask <= rob_uop__8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_42) begin
      rob_uop__9_uopc <= io_enq_uops_0_uopc;
      rob_uop__9_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__9_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__9_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__9_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__9_pdst <= io_enq_uops_0_pdst;
      rob_uop__9_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__9_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__9_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__9_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__9_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__9_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__9_ldst <= io_enq_uops_0_ldst;
      rob_uop__9_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__9_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__9_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2519) | ~rob_val__9) begin
      if (_GEN_42)
        rob_uop__9_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__9_br_mask <= rob_uop__9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_43) begin
      rob_uop__10_uopc <= io_enq_uops_0_uopc;
      rob_uop__10_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__10_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__10_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__10_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__10_pdst <= io_enq_uops_0_pdst;
      rob_uop__10_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__10_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__10_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__10_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__10_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__10_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__10_ldst <= io_enq_uops_0_ldst;
      rob_uop__10_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__10_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__10_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2520) | ~rob_val__10) begin
      if (_GEN_43)
        rob_uop__10_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__10_br_mask <= rob_uop__10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_44) begin
      rob_uop__11_uopc <= io_enq_uops_0_uopc;
      rob_uop__11_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__11_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__11_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__11_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__11_pdst <= io_enq_uops_0_pdst;
      rob_uop__11_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__11_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__11_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__11_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__11_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__11_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__11_ldst <= io_enq_uops_0_ldst;
      rob_uop__11_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__11_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__11_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2521) | ~rob_val__11) begin
      if (_GEN_44)
        rob_uop__11_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__11_br_mask <= rob_uop__11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_45) begin
      rob_uop__12_uopc <= io_enq_uops_0_uopc;
      rob_uop__12_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__12_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__12_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__12_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__12_pdst <= io_enq_uops_0_pdst;
      rob_uop__12_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__12_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__12_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__12_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__12_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__12_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__12_ldst <= io_enq_uops_0_ldst;
      rob_uop__12_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__12_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__12_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2522) | ~rob_val__12) begin
      if (_GEN_45)
        rob_uop__12_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__12_br_mask <= rob_uop__12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_46) begin
      rob_uop__13_uopc <= io_enq_uops_0_uopc;
      rob_uop__13_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__13_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__13_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__13_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__13_pdst <= io_enq_uops_0_pdst;
      rob_uop__13_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__13_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__13_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__13_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__13_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__13_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__13_ldst <= io_enq_uops_0_ldst;
      rob_uop__13_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__13_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__13_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2523) | ~rob_val__13) begin
      if (_GEN_46)
        rob_uop__13_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__13_br_mask <= rob_uop__13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_47) begin
      rob_uop__14_uopc <= io_enq_uops_0_uopc;
      rob_uop__14_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__14_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__14_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__14_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__14_pdst <= io_enq_uops_0_pdst;
      rob_uop__14_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__14_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__14_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__14_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__14_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__14_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__14_ldst <= io_enq_uops_0_ldst;
      rob_uop__14_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__14_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__14_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2524) | ~rob_val__14) begin
      if (_GEN_47)
        rob_uop__14_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__14_br_mask <= rob_uop__14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_48) begin
      rob_uop__15_uopc <= io_enq_uops_0_uopc;
      rob_uop__15_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__15_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__15_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__15_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__15_pdst <= io_enq_uops_0_pdst;
      rob_uop__15_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__15_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__15_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__15_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__15_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__15_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__15_ldst <= io_enq_uops_0_ldst;
      rob_uop__15_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__15_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__15_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2525) | ~rob_val__15) begin
      if (_GEN_48)
        rob_uop__15_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__15_br_mask <= rob_uop__15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_49) begin
      rob_uop__16_uopc <= io_enq_uops_0_uopc;
      rob_uop__16_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__16_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__16_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__16_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__16_pdst <= io_enq_uops_0_pdst;
      rob_uop__16_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__16_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__16_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__16_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__16_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__16_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__16_ldst <= io_enq_uops_0_ldst;
      rob_uop__16_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__16_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__16_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2526) | ~rob_val__16) begin
      if (_GEN_49)
        rob_uop__16_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__16_br_mask <= rob_uop__16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_50) begin
      rob_uop__17_uopc <= io_enq_uops_0_uopc;
      rob_uop__17_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__17_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__17_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__17_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__17_pdst <= io_enq_uops_0_pdst;
      rob_uop__17_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__17_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__17_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__17_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__17_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__17_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__17_ldst <= io_enq_uops_0_ldst;
      rob_uop__17_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__17_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__17_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2527) | ~rob_val__17) begin
      if (_GEN_50)
        rob_uop__17_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__17_br_mask <= rob_uop__17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_51) begin
      rob_uop__18_uopc <= io_enq_uops_0_uopc;
      rob_uop__18_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__18_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__18_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__18_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__18_pdst <= io_enq_uops_0_pdst;
      rob_uop__18_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__18_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__18_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__18_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__18_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__18_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__18_ldst <= io_enq_uops_0_ldst;
      rob_uop__18_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__18_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__18_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2528) | ~rob_val__18) begin
      if (_GEN_51)
        rob_uop__18_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__18_br_mask <= rob_uop__18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_52) begin
      rob_uop__19_uopc <= io_enq_uops_0_uopc;
      rob_uop__19_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__19_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__19_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__19_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__19_pdst <= io_enq_uops_0_pdst;
      rob_uop__19_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__19_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__19_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__19_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__19_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__19_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__19_ldst <= io_enq_uops_0_ldst;
      rob_uop__19_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__19_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__19_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2529) | ~rob_val__19) begin
      if (_GEN_52)
        rob_uop__19_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__19_br_mask <= rob_uop__19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_53) begin
      rob_uop__20_uopc <= io_enq_uops_0_uopc;
      rob_uop__20_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__20_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__20_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__20_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__20_pdst <= io_enq_uops_0_pdst;
      rob_uop__20_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__20_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__20_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__20_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__20_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__20_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__20_ldst <= io_enq_uops_0_ldst;
      rob_uop__20_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__20_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__20_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2530) | ~rob_val__20) begin
      if (_GEN_53)
        rob_uop__20_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__20_br_mask <= rob_uop__20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_54) begin
      rob_uop__21_uopc <= io_enq_uops_0_uopc;
      rob_uop__21_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__21_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__21_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__21_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__21_pdst <= io_enq_uops_0_pdst;
      rob_uop__21_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__21_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__21_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__21_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__21_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__21_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__21_ldst <= io_enq_uops_0_ldst;
      rob_uop__21_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__21_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__21_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2531) | ~rob_val__21) begin
      if (_GEN_54)
        rob_uop__21_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__21_br_mask <= rob_uop__21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_55) begin
      rob_uop__22_uopc <= io_enq_uops_0_uopc;
      rob_uop__22_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__22_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__22_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__22_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__22_pdst <= io_enq_uops_0_pdst;
      rob_uop__22_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__22_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__22_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__22_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__22_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__22_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__22_ldst <= io_enq_uops_0_ldst;
      rob_uop__22_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__22_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__22_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2532) | ~rob_val__22) begin
      if (_GEN_55)
        rob_uop__22_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__22_br_mask <= rob_uop__22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_56) begin
      rob_uop__23_uopc <= io_enq_uops_0_uopc;
      rob_uop__23_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__23_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__23_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__23_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__23_pdst <= io_enq_uops_0_pdst;
      rob_uop__23_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__23_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__23_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__23_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__23_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__23_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__23_ldst <= io_enq_uops_0_ldst;
      rob_uop__23_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__23_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__23_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2533) | ~rob_val__23) begin
      if (_GEN_56)
        rob_uop__23_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__23_br_mask <= rob_uop__23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_57) begin
      rob_uop__24_uopc <= io_enq_uops_0_uopc;
      rob_uop__24_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__24_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__24_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__24_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__24_pdst <= io_enq_uops_0_pdst;
      rob_uop__24_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__24_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__24_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__24_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__24_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__24_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__24_ldst <= io_enq_uops_0_ldst;
      rob_uop__24_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__24_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__24_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2534) | ~rob_val__24) begin
      if (_GEN_57)
        rob_uop__24_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__24_br_mask <= rob_uop__24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_58) begin
      rob_uop__25_uopc <= io_enq_uops_0_uopc;
      rob_uop__25_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__25_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__25_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__25_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__25_pdst <= io_enq_uops_0_pdst;
      rob_uop__25_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__25_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__25_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__25_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__25_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__25_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__25_ldst <= io_enq_uops_0_ldst;
      rob_uop__25_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__25_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__25_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2535) | ~rob_val__25) begin
      if (_GEN_58)
        rob_uop__25_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__25_br_mask <= rob_uop__25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_59) begin
      rob_uop__26_uopc <= io_enq_uops_0_uopc;
      rob_uop__26_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__26_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__26_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__26_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__26_pdst <= io_enq_uops_0_pdst;
      rob_uop__26_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__26_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__26_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__26_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__26_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__26_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__26_ldst <= io_enq_uops_0_ldst;
      rob_uop__26_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__26_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__26_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2536) | ~rob_val__26) begin
      if (_GEN_59)
        rob_uop__26_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__26_br_mask <= rob_uop__26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_60) begin
      rob_uop__27_uopc <= io_enq_uops_0_uopc;
      rob_uop__27_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__27_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__27_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__27_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__27_pdst <= io_enq_uops_0_pdst;
      rob_uop__27_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__27_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__27_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__27_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__27_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__27_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__27_ldst <= io_enq_uops_0_ldst;
      rob_uop__27_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__27_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__27_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2537) | ~rob_val__27) begin
      if (_GEN_60)
        rob_uop__27_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__27_br_mask <= rob_uop__27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_61) begin
      rob_uop__28_uopc <= io_enq_uops_0_uopc;
      rob_uop__28_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__28_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__28_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__28_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__28_pdst <= io_enq_uops_0_pdst;
      rob_uop__28_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__28_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__28_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__28_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__28_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__28_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__28_ldst <= io_enq_uops_0_ldst;
      rob_uop__28_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__28_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__28_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2538) | ~rob_val__28) begin
      if (_GEN_61)
        rob_uop__28_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__28_br_mask <= rob_uop__28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_62) begin
      rob_uop__29_uopc <= io_enq_uops_0_uopc;
      rob_uop__29_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__29_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__29_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__29_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__29_pdst <= io_enq_uops_0_pdst;
      rob_uop__29_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__29_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__29_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__29_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__29_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__29_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__29_ldst <= io_enq_uops_0_ldst;
      rob_uop__29_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__29_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__29_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2539) | ~rob_val__29) begin
      if (_GEN_62)
        rob_uop__29_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__29_br_mask <= rob_uop__29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_63) begin
      rob_uop__30_uopc <= io_enq_uops_0_uopc;
      rob_uop__30_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__30_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__30_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__30_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__30_pdst <= io_enq_uops_0_pdst;
      rob_uop__30_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__30_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__30_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__30_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__30_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__30_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__30_ldst <= io_enq_uops_0_ldst;
      rob_uop__30_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__30_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__30_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2540) | ~rob_val__30) begin
      if (_GEN_63)
        rob_uop__30_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__30_br_mask <= rob_uop__30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_64) begin
      rob_uop__31_uopc <= io_enq_uops_0_uopc;
      rob_uop__31_is_rvc <= io_enq_uops_0_is_rvc;
      rob_uop__31_ftq_idx <= io_enq_uops_0_ftq_idx;
      rob_uop__31_edge_inst <= io_enq_uops_0_edge_inst;
      rob_uop__31_pc_lob <= io_enq_uops_0_pc_lob;
      rob_uop__31_pdst <= io_enq_uops_0_pdst;
      rob_uop__31_stale_pdst <= io_enq_uops_0_stale_pdst;
      rob_uop__31_is_fencei <= io_enq_uops_0_is_fencei;
      rob_uop__31_uses_ldq <= io_enq_uops_0_uses_ldq;
      rob_uop__31_uses_stq <= io_enq_uops_0_uses_stq;
      rob_uop__31_is_sys_pc2epc <= io_enq_uops_0_is_sys_pc2epc;
      rob_uop__31_flush_on_commit <= io_enq_uops_0_flush_on_commit;
      rob_uop__31_ldst <= io_enq_uops_0_ldst;
      rob_uop__31_ldst_val <= io_enq_uops_0_ldst_val;
      rob_uop__31_dst_rtype <= io_enq_uops_0_dst_rtype;
      rob_uop__31_fp_val <= io_enq_uops_0_fp_val;
    end
    if ((|_GEN_2541) | ~rob_val__31) begin
      if (_GEN_64)
        rob_uop__31_br_mask <= io_enq_uops_0_br_mask;
    end
    else
      rob_uop__31_br_mask <= rob_uop__31_br_mask & ~io_brupdate_b1_resolve_mask;
    rob_predicated__0 <= ~(_GEN_641 & _GEN_642 | _GEN_609 | _GEN_513 & _GEN_514) & (_GEN_481 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_386 | _GEN_353 | _GEN_257 & _GEN_258 | _GEN_225 | _GEN_129 & _GEN_130) & (_GEN_97 ? io_wb_resps_0_bits_predicated : ~_GEN_33 & rob_predicated__0));
    rob_predicated__1 <= ~(_GEN_641 & _GEN_644 | _GEN_610 | _GEN_513 & _GEN_516) & (_GEN_482 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_388 | _GEN_354 | _GEN_257 & _GEN_260 | _GEN_226 | _GEN_129 & _GEN_132) & (_GEN_98 ? io_wb_resps_0_bits_predicated : ~_GEN_34 & rob_predicated__1));
    rob_predicated__2 <= ~(_GEN_641 & _GEN_646 | _GEN_611 | _GEN_513 & _GEN_518) & (_GEN_483 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_390 | _GEN_355 | _GEN_257 & _GEN_262 | _GEN_227 | _GEN_129 & _GEN_134) & (_GEN_99 ? io_wb_resps_0_bits_predicated : ~_GEN_35 & rob_predicated__2));
    rob_predicated__3 <= ~(_GEN_641 & _GEN_648 | _GEN_612 | _GEN_513 & _GEN_520) & (_GEN_484 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_392 | _GEN_356 | _GEN_257 & _GEN_264 | _GEN_228 | _GEN_129 & _GEN_136) & (_GEN_100 ? io_wb_resps_0_bits_predicated : ~_GEN_36 & rob_predicated__3));
    rob_predicated__4 <= ~(_GEN_641 & _GEN_650 | _GEN_613 | _GEN_513 & _GEN_522) & (_GEN_485 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_394 | _GEN_357 | _GEN_257 & _GEN_266 | _GEN_229 | _GEN_129 & _GEN_138) & (_GEN_101 ? io_wb_resps_0_bits_predicated : ~_GEN_37 & rob_predicated__4));
    rob_predicated__5 <= ~(_GEN_641 & _GEN_652 | _GEN_614 | _GEN_513 & _GEN_524) & (_GEN_486 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_396 | _GEN_358 | _GEN_257 & _GEN_268 | _GEN_230 | _GEN_129 & _GEN_140) & (_GEN_102 ? io_wb_resps_0_bits_predicated : ~_GEN_38 & rob_predicated__5));
    rob_predicated__6 <= ~(_GEN_641 & _GEN_654 | _GEN_615 | _GEN_513 & _GEN_526) & (_GEN_487 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_398 | _GEN_359 | _GEN_257 & _GEN_270 | _GEN_231 | _GEN_129 & _GEN_142) & (_GEN_103 ? io_wb_resps_0_bits_predicated : ~_GEN_39 & rob_predicated__6));
    rob_predicated__7 <= ~(_GEN_641 & _GEN_656 | _GEN_616 | _GEN_513 & _GEN_528) & (_GEN_488 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_400 | _GEN_360 | _GEN_257 & _GEN_272 | _GEN_232 | _GEN_129 & _GEN_144) & (_GEN_104 ? io_wb_resps_0_bits_predicated : ~_GEN_40 & rob_predicated__7));
    rob_predicated__8 <= ~(_GEN_641 & _GEN_658 | _GEN_617 | _GEN_513 & _GEN_530) & (_GEN_489 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_402 | _GEN_361 | _GEN_257 & _GEN_274 | _GEN_233 | _GEN_129 & _GEN_146) & (_GEN_105 ? io_wb_resps_0_bits_predicated : ~_GEN_41 & rob_predicated__8));
    rob_predicated__9 <= ~(_GEN_641 & _GEN_660 | _GEN_618 | _GEN_513 & _GEN_532) & (_GEN_490 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_404 | _GEN_362 | _GEN_257 & _GEN_276 | _GEN_234 | _GEN_129 & _GEN_148) & (_GEN_106 ? io_wb_resps_0_bits_predicated : ~_GEN_42 & rob_predicated__9));
    rob_predicated__10 <= ~(_GEN_641 & _GEN_662 | _GEN_619 | _GEN_513 & _GEN_534) & (_GEN_491 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_406 | _GEN_363 | _GEN_257 & _GEN_278 | _GEN_235 | _GEN_129 & _GEN_150) & (_GEN_107 ? io_wb_resps_0_bits_predicated : ~_GEN_43 & rob_predicated__10));
    rob_predicated__11 <= ~(_GEN_641 & _GEN_664 | _GEN_620 | _GEN_513 & _GEN_536) & (_GEN_492 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_408 | _GEN_364 | _GEN_257 & _GEN_280 | _GEN_236 | _GEN_129 & _GEN_152) & (_GEN_108 ? io_wb_resps_0_bits_predicated : ~_GEN_44 & rob_predicated__11));
    rob_predicated__12 <= ~(_GEN_641 & _GEN_666 | _GEN_621 | _GEN_513 & _GEN_538) & (_GEN_493 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_410 | _GEN_365 | _GEN_257 & _GEN_282 | _GEN_237 | _GEN_129 & _GEN_154) & (_GEN_109 ? io_wb_resps_0_bits_predicated : ~_GEN_45 & rob_predicated__12));
    rob_predicated__13 <= ~(_GEN_641 & _GEN_668 | _GEN_622 | _GEN_513 & _GEN_540) & (_GEN_494 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_412 | _GEN_366 | _GEN_257 & _GEN_284 | _GEN_238 | _GEN_129 & _GEN_156) & (_GEN_110 ? io_wb_resps_0_bits_predicated : ~_GEN_46 & rob_predicated__13));
    rob_predicated__14 <= ~(_GEN_641 & _GEN_670 | _GEN_623 | _GEN_513 & _GEN_542) & (_GEN_495 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_414 | _GEN_367 | _GEN_257 & _GEN_286 | _GEN_239 | _GEN_129 & _GEN_158) & (_GEN_111 ? io_wb_resps_0_bits_predicated : ~_GEN_47 & rob_predicated__14));
    rob_predicated__15 <= ~(_GEN_641 & _GEN_672 | _GEN_624 | _GEN_513 & _GEN_544) & (_GEN_496 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_416 | _GEN_368 | _GEN_257 & _GEN_288 | _GEN_240 | _GEN_129 & _GEN_160) & (_GEN_112 ? io_wb_resps_0_bits_predicated : ~_GEN_48 & rob_predicated__15));
    rob_predicated__16 <= ~(_GEN_641 & _GEN_674 | _GEN_625 | _GEN_513 & _GEN_546) & (_GEN_497 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_418 | _GEN_369 | _GEN_257 & _GEN_290 | _GEN_241 | _GEN_129 & _GEN_162) & (_GEN_113 ? io_wb_resps_0_bits_predicated : ~_GEN_49 & rob_predicated__16));
    rob_predicated__17 <= ~(_GEN_641 & _GEN_676 | _GEN_626 | _GEN_513 & _GEN_548) & (_GEN_498 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_420 | _GEN_370 | _GEN_257 & _GEN_292 | _GEN_242 | _GEN_129 & _GEN_164) & (_GEN_114 ? io_wb_resps_0_bits_predicated : ~_GEN_50 & rob_predicated__17));
    rob_predicated__18 <= ~(_GEN_641 & _GEN_678 | _GEN_627 | _GEN_513 & _GEN_550) & (_GEN_499 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_422 | _GEN_371 | _GEN_257 & _GEN_294 | _GEN_243 | _GEN_129 & _GEN_166) & (_GEN_115 ? io_wb_resps_0_bits_predicated : ~_GEN_51 & rob_predicated__18));
    rob_predicated__19 <= ~(_GEN_641 & _GEN_680 | _GEN_628 | _GEN_513 & _GEN_552) & (_GEN_500 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_424 | _GEN_372 | _GEN_257 & _GEN_296 | _GEN_244 | _GEN_129 & _GEN_168) & (_GEN_116 ? io_wb_resps_0_bits_predicated : ~_GEN_52 & rob_predicated__19));
    rob_predicated__20 <= ~(_GEN_641 & _GEN_682 | _GEN_629 | _GEN_513 & _GEN_554) & (_GEN_501 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_426 | _GEN_373 | _GEN_257 & _GEN_298 | _GEN_245 | _GEN_129 & _GEN_170) & (_GEN_117 ? io_wb_resps_0_bits_predicated : ~_GEN_53 & rob_predicated__20));
    rob_predicated__21 <= ~(_GEN_641 & _GEN_684 | _GEN_630 | _GEN_513 & _GEN_556) & (_GEN_502 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_428 | _GEN_374 | _GEN_257 & _GEN_300 | _GEN_246 | _GEN_129 & _GEN_172) & (_GEN_118 ? io_wb_resps_0_bits_predicated : ~_GEN_54 & rob_predicated__21));
    rob_predicated__22 <= ~(_GEN_641 & _GEN_686 | _GEN_631 | _GEN_513 & _GEN_558) & (_GEN_503 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_430 | _GEN_375 | _GEN_257 & _GEN_302 | _GEN_247 | _GEN_129 & _GEN_174) & (_GEN_119 ? io_wb_resps_0_bits_predicated : ~_GEN_55 & rob_predicated__22));
    rob_predicated__23 <= ~(_GEN_641 & _GEN_688 | _GEN_632 | _GEN_513 & _GEN_560) & (_GEN_504 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_432 | _GEN_376 | _GEN_257 & _GEN_304 | _GEN_248 | _GEN_129 & _GEN_176) & (_GEN_120 ? io_wb_resps_0_bits_predicated : ~_GEN_56 & rob_predicated__23));
    rob_predicated__24 <= ~(_GEN_641 & _GEN_690 | _GEN_633 | _GEN_513 & _GEN_562) & (_GEN_505 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_434 | _GEN_377 | _GEN_257 & _GEN_306 | _GEN_249 | _GEN_129 & _GEN_178) & (_GEN_121 ? io_wb_resps_0_bits_predicated : ~_GEN_57 & rob_predicated__24));
    rob_predicated__25 <= ~(_GEN_641 & _GEN_692 | _GEN_634 | _GEN_513 & _GEN_564) & (_GEN_506 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_436 | _GEN_378 | _GEN_257 & _GEN_308 | _GEN_250 | _GEN_129 & _GEN_180) & (_GEN_122 ? io_wb_resps_0_bits_predicated : ~_GEN_58 & rob_predicated__25));
    rob_predicated__26 <= ~(_GEN_641 & _GEN_694 | _GEN_635 | _GEN_513 & _GEN_566) & (_GEN_507 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_438 | _GEN_379 | _GEN_257 & _GEN_310 | _GEN_251 | _GEN_129 & _GEN_182) & (_GEN_123 ? io_wb_resps_0_bits_predicated : ~_GEN_59 & rob_predicated__26));
    rob_predicated__27 <= ~(_GEN_641 & _GEN_696 | _GEN_636 | _GEN_513 & _GEN_568) & (_GEN_508 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_440 | _GEN_380 | _GEN_257 & _GEN_312 | _GEN_252 | _GEN_129 & _GEN_184) & (_GEN_124 ? io_wb_resps_0_bits_predicated : ~_GEN_60 & rob_predicated__27));
    rob_predicated__28 <= ~(_GEN_641 & _GEN_698 | _GEN_637 | _GEN_513 & _GEN_570) & (_GEN_509 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_442 | _GEN_381 | _GEN_257 & _GEN_314 | _GEN_253 | _GEN_129 & _GEN_186) & (_GEN_125 ? io_wb_resps_0_bits_predicated : ~_GEN_61 & rob_predicated__28));
    rob_predicated__29 <= ~(_GEN_641 & _GEN_700 | _GEN_638 | _GEN_513 & _GEN_572) & (_GEN_510 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_444 | _GEN_382 | _GEN_257 & _GEN_316 | _GEN_254 | _GEN_129 & _GEN_188) & (_GEN_126 ? io_wb_resps_0_bits_predicated : ~_GEN_62 & rob_predicated__29));
    rob_predicated__30 <= ~(_GEN_641 & _GEN_702 | _GEN_639 | _GEN_513 & _GEN_574) & (_GEN_511 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & _GEN_446 | _GEN_383 | _GEN_257 & _GEN_318 | _GEN_255 | _GEN_129 & _GEN_190) & (_GEN_127 ? io_wb_resps_0_bits_predicated : ~_GEN_63 & rob_predicated__30));
    rob_predicated__31 <= ~(_GEN_641 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_640 | _GEN_513 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_512 ? io_wb_resps_6_bits_predicated : ~(_GEN_385 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_384 | _GEN_257 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_256 | _GEN_129 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_128 ? io_wb_resps_0_bits_predicated : ~_GEN_64 & rob_predicated__31));
    if (_GEN_898) begin
      rob_uop_1_0_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_0_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_0_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_0_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_0_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_0_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_0_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_0_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_0_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_0_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_0_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_0_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_0_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_0_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_0_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_0_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2577) | ~rob_val_1_0) begin
      if (_GEN_898)
        rob_uop_1_0_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_0_br_mask <= rob_uop_1_0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_899) begin
      rob_uop_1_1_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_1_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_1_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_1_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_1_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_1_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_1_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_1_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_1_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_1_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_1_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_1_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_1_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_1_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_1_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_1_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2578) | ~rob_val_1_1) begin
      if (_GEN_899)
        rob_uop_1_1_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_1_br_mask <= rob_uop_1_1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_900) begin
      rob_uop_1_2_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_2_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_2_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_2_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_2_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_2_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_2_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_2_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_2_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_2_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_2_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_2_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_2_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_2_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_2_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_2_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2579) | ~rob_val_1_2) begin
      if (_GEN_900)
        rob_uop_1_2_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_2_br_mask <= rob_uop_1_2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_901) begin
      rob_uop_1_3_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_3_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_3_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_3_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_3_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_3_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_3_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_3_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_3_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_3_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_3_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_3_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_3_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_3_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_3_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_3_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2580) | ~rob_val_1_3) begin
      if (_GEN_901)
        rob_uop_1_3_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_3_br_mask <= rob_uop_1_3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_902) begin
      rob_uop_1_4_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_4_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_4_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_4_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_4_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_4_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_4_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_4_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_4_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_4_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_4_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_4_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_4_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_4_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_4_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_4_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2581) | ~rob_val_1_4) begin
      if (_GEN_902)
        rob_uop_1_4_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_4_br_mask <= rob_uop_1_4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_903) begin
      rob_uop_1_5_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_5_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_5_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_5_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_5_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_5_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_5_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_5_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_5_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_5_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_5_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_5_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_5_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_5_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_5_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_5_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2582) | ~rob_val_1_5) begin
      if (_GEN_903)
        rob_uop_1_5_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_5_br_mask <= rob_uop_1_5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_904) begin
      rob_uop_1_6_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_6_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_6_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_6_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_6_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_6_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_6_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_6_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_6_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_6_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_6_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_6_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_6_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_6_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_6_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_6_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2583) | ~rob_val_1_6) begin
      if (_GEN_904)
        rob_uop_1_6_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_6_br_mask <= rob_uop_1_6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_905) begin
      rob_uop_1_7_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_7_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_7_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_7_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_7_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_7_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_7_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_7_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_7_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_7_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_7_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_7_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_7_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_7_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_7_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_7_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2584) | ~rob_val_1_7) begin
      if (_GEN_905)
        rob_uop_1_7_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_7_br_mask <= rob_uop_1_7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_906) begin
      rob_uop_1_8_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_8_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_8_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_8_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_8_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_8_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_8_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_8_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_8_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_8_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_8_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_8_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_8_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_8_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_8_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_8_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2585) | ~rob_val_1_8) begin
      if (_GEN_906)
        rob_uop_1_8_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_8_br_mask <= rob_uop_1_8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_907) begin
      rob_uop_1_9_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_9_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_9_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_9_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_9_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_9_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_9_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_9_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_9_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_9_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_9_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_9_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_9_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_9_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_9_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_9_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2586) | ~rob_val_1_9) begin
      if (_GEN_907)
        rob_uop_1_9_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_9_br_mask <= rob_uop_1_9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_908) begin
      rob_uop_1_10_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_10_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_10_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_10_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_10_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_10_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_10_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_10_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_10_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_10_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_10_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_10_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_10_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_10_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_10_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_10_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2587) | ~rob_val_1_10) begin
      if (_GEN_908)
        rob_uop_1_10_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_10_br_mask <= rob_uop_1_10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_909) begin
      rob_uop_1_11_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_11_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_11_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_11_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_11_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_11_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_11_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_11_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_11_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_11_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_11_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_11_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_11_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_11_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_11_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_11_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2588) | ~rob_val_1_11) begin
      if (_GEN_909)
        rob_uop_1_11_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_11_br_mask <= rob_uop_1_11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_910) begin
      rob_uop_1_12_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_12_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_12_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_12_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_12_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_12_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_12_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_12_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_12_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_12_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_12_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_12_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_12_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_12_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_12_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_12_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2589) | ~rob_val_1_12) begin
      if (_GEN_910)
        rob_uop_1_12_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_12_br_mask <= rob_uop_1_12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_911) begin
      rob_uop_1_13_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_13_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_13_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_13_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_13_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_13_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_13_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_13_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_13_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_13_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_13_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_13_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_13_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_13_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_13_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_13_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2590) | ~rob_val_1_13) begin
      if (_GEN_911)
        rob_uop_1_13_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_13_br_mask <= rob_uop_1_13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_912) begin
      rob_uop_1_14_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_14_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_14_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_14_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_14_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_14_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_14_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_14_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_14_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_14_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_14_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_14_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_14_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_14_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_14_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_14_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2591) | ~rob_val_1_14) begin
      if (_GEN_912)
        rob_uop_1_14_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_14_br_mask <= rob_uop_1_14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_913) begin
      rob_uop_1_15_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_15_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_15_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_15_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_15_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_15_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_15_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_15_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_15_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_15_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_15_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_15_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_15_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_15_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_15_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_15_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2592) | ~rob_val_1_15) begin
      if (_GEN_913)
        rob_uop_1_15_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_15_br_mask <= rob_uop_1_15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_914) begin
      rob_uop_1_16_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_16_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_16_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_16_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_16_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_16_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_16_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_16_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_16_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_16_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_16_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_16_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_16_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_16_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_16_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_16_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2593) | ~rob_val_1_16) begin
      if (_GEN_914)
        rob_uop_1_16_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_16_br_mask <= rob_uop_1_16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_915) begin
      rob_uop_1_17_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_17_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_17_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_17_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_17_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_17_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_17_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_17_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_17_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_17_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_17_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_17_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_17_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_17_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_17_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_17_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2594) | ~rob_val_1_17) begin
      if (_GEN_915)
        rob_uop_1_17_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_17_br_mask <= rob_uop_1_17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_916) begin
      rob_uop_1_18_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_18_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_18_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_18_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_18_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_18_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_18_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_18_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_18_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_18_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_18_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_18_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_18_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_18_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_18_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_18_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2595) | ~rob_val_1_18) begin
      if (_GEN_916)
        rob_uop_1_18_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_18_br_mask <= rob_uop_1_18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_917) begin
      rob_uop_1_19_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_19_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_19_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_19_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_19_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_19_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_19_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_19_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_19_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_19_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_19_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_19_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_19_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_19_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_19_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_19_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2596) | ~rob_val_1_19) begin
      if (_GEN_917)
        rob_uop_1_19_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_19_br_mask <= rob_uop_1_19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_918) begin
      rob_uop_1_20_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_20_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_20_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_20_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_20_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_20_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_20_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_20_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_20_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_20_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_20_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_20_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_20_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_20_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_20_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_20_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2597) | ~rob_val_1_20) begin
      if (_GEN_918)
        rob_uop_1_20_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_20_br_mask <= rob_uop_1_20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_919) begin
      rob_uop_1_21_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_21_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_21_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_21_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_21_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_21_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_21_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_21_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_21_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_21_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_21_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_21_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_21_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_21_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_21_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_21_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2598) | ~rob_val_1_21) begin
      if (_GEN_919)
        rob_uop_1_21_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_21_br_mask <= rob_uop_1_21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_920) begin
      rob_uop_1_22_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_22_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_22_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_22_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_22_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_22_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_22_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_22_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_22_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_22_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_22_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_22_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_22_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_22_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_22_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_22_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2599) | ~rob_val_1_22) begin
      if (_GEN_920)
        rob_uop_1_22_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_22_br_mask <= rob_uop_1_22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_921) begin
      rob_uop_1_23_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_23_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_23_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_23_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_23_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_23_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_23_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_23_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_23_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_23_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_23_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_23_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_23_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_23_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_23_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_23_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2600) | ~rob_val_1_23) begin
      if (_GEN_921)
        rob_uop_1_23_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_23_br_mask <= rob_uop_1_23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_922) begin
      rob_uop_1_24_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_24_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_24_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_24_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_24_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_24_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_24_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_24_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_24_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_24_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_24_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_24_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_24_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_24_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_24_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_24_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2601) | ~rob_val_1_24) begin
      if (_GEN_922)
        rob_uop_1_24_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_24_br_mask <= rob_uop_1_24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_923) begin
      rob_uop_1_25_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_25_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_25_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_25_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_25_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_25_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_25_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_25_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_25_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_25_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_25_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_25_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_25_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_25_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_25_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_25_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2602) | ~rob_val_1_25) begin
      if (_GEN_923)
        rob_uop_1_25_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_25_br_mask <= rob_uop_1_25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_924) begin
      rob_uop_1_26_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_26_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_26_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_26_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_26_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_26_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_26_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_26_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_26_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_26_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_26_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_26_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_26_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_26_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_26_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_26_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2603) | ~rob_val_1_26) begin
      if (_GEN_924)
        rob_uop_1_26_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_26_br_mask <= rob_uop_1_26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_925) begin
      rob_uop_1_27_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_27_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_27_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_27_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_27_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_27_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_27_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_27_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_27_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_27_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_27_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_27_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_27_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_27_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_27_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_27_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2604) | ~rob_val_1_27) begin
      if (_GEN_925)
        rob_uop_1_27_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_27_br_mask <= rob_uop_1_27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_926) begin
      rob_uop_1_28_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_28_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_28_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_28_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_28_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_28_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_28_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_28_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_28_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_28_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_28_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_28_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_28_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_28_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_28_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_28_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2605) | ~rob_val_1_28) begin
      if (_GEN_926)
        rob_uop_1_28_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_28_br_mask <= rob_uop_1_28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_927) begin
      rob_uop_1_29_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_29_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_29_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_29_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_29_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_29_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_29_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_29_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_29_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_29_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_29_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_29_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_29_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_29_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_29_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_29_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2606) | ~rob_val_1_29) begin
      if (_GEN_927)
        rob_uop_1_29_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_29_br_mask <= rob_uop_1_29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_928) begin
      rob_uop_1_30_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_30_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_30_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_30_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_30_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_30_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_30_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_30_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_30_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_30_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_30_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_30_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_30_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_30_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_30_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_30_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2607) | ~rob_val_1_30) begin
      if (_GEN_928)
        rob_uop_1_30_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_30_br_mask <= rob_uop_1_30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_929) begin
      rob_uop_1_31_uopc <= io_enq_uops_1_uopc;
      rob_uop_1_31_is_rvc <= io_enq_uops_1_is_rvc;
      rob_uop_1_31_ftq_idx <= io_enq_uops_1_ftq_idx;
      rob_uop_1_31_edge_inst <= io_enq_uops_1_edge_inst;
      rob_uop_1_31_pc_lob <= io_enq_uops_1_pc_lob;
      rob_uop_1_31_pdst <= io_enq_uops_1_pdst;
      rob_uop_1_31_stale_pdst <= io_enq_uops_1_stale_pdst;
      rob_uop_1_31_is_fencei <= io_enq_uops_1_is_fencei;
      rob_uop_1_31_uses_ldq <= io_enq_uops_1_uses_ldq;
      rob_uop_1_31_uses_stq <= io_enq_uops_1_uses_stq;
      rob_uop_1_31_is_sys_pc2epc <= io_enq_uops_1_is_sys_pc2epc;
      rob_uop_1_31_flush_on_commit <= io_enq_uops_1_flush_on_commit;
      rob_uop_1_31_ldst <= io_enq_uops_1_ldst;
      rob_uop_1_31_ldst_val <= io_enq_uops_1_ldst_val;
      rob_uop_1_31_dst_rtype <= io_enq_uops_1_dst_rtype;
      rob_uop_1_31_fp_val <= io_enq_uops_1_fp_val;
    end
    if ((|_GEN_2608) | ~rob_val_1_31) begin
      if (_GEN_929)
        rob_uop_1_31_br_mask <= io_enq_uops_1_br_mask;
    end
    else
      rob_uop_1_31_br_mask <= rob_uop_1_31_br_mask & ~io_brupdate_b1_resolve_mask;
    rob_predicated_1_0 <= ~(_GEN_1227 & _GEN_642 | _GEN_1195 | _GEN_1161 & _GEN_514) & (_GEN_1129 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_386 | _GEN_1063 | _GEN_1029 & _GEN_258 | _GEN_997 | _GEN_963 & _GEN_130) & (_GEN_931 ? io_wb_resps_0_bits_predicated : ~_GEN_898 & rob_predicated_1_0));
    rob_predicated_1_1 <= ~(_GEN_1227 & _GEN_644 | _GEN_1196 | _GEN_1161 & _GEN_516) & (_GEN_1130 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_388 | _GEN_1064 | _GEN_1029 & _GEN_260 | _GEN_998 | _GEN_963 & _GEN_132) & (_GEN_932 ? io_wb_resps_0_bits_predicated : ~_GEN_899 & rob_predicated_1_1));
    rob_predicated_1_2 <= ~(_GEN_1227 & _GEN_646 | _GEN_1197 | _GEN_1161 & _GEN_518) & (_GEN_1131 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_390 | _GEN_1065 | _GEN_1029 & _GEN_262 | _GEN_999 | _GEN_963 & _GEN_134) & (_GEN_933 ? io_wb_resps_0_bits_predicated : ~_GEN_900 & rob_predicated_1_2));
    rob_predicated_1_3 <= ~(_GEN_1227 & _GEN_648 | _GEN_1198 | _GEN_1161 & _GEN_520) & (_GEN_1132 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_392 | _GEN_1066 | _GEN_1029 & _GEN_264 | _GEN_1000 | _GEN_963 & _GEN_136) & (_GEN_934 ? io_wb_resps_0_bits_predicated : ~_GEN_901 & rob_predicated_1_3));
    rob_predicated_1_4 <= ~(_GEN_1227 & _GEN_650 | _GEN_1199 | _GEN_1161 & _GEN_522) & (_GEN_1133 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_394 | _GEN_1067 | _GEN_1029 & _GEN_266 | _GEN_1001 | _GEN_963 & _GEN_138) & (_GEN_935 ? io_wb_resps_0_bits_predicated : ~_GEN_902 & rob_predicated_1_4));
    rob_predicated_1_5 <= ~(_GEN_1227 & _GEN_652 | _GEN_1200 | _GEN_1161 & _GEN_524) & (_GEN_1134 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_396 | _GEN_1068 | _GEN_1029 & _GEN_268 | _GEN_1002 | _GEN_963 & _GEN_140) & (_GEN_936 ? io_wb_resps_0_bits_predicated : ~_GEN_903 & rob_predicated_1_5));
    rob_predicated_1_6 <= ~(_GEN_1227 & _GEN_654 | _GEN_1201 | _GEN_1161 & _GEN_526) & (_GEN_1135 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_398 | _GEN_1069 | _GEN_1029 & _GEN_270 | _GEN_1003 | _GEN_963 & _GEN_142) & (_GEN_937 ? io_wb_resps_0_bits_predicated : ~_GEN_904 & rob_predicated_1_6));
    rob_predicated_1_7 <= ~(_GEN_1227 & _GEN_656 | _GEN_1202 | _GEN_1161 & _GEN_528) & (_GEN_1136 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_400 | _GEN_1070 | _GEN_1029 & _GEN_272 | _GEN_1004 | _GEN_963 & _GEN_144) & (_GEN_938 ? io_wb_resps_0_bits_predicated : ~_GEN_905 & rob_predicated_1_7));
    rob_predicated_1_8 <= ~(_GEN_1227 & _GEN_658 | _GEN_1203 | _GEN_1161 & _GEN_530) & (_GEN_1137 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_402 | _GEN_1071 | _GEN_1029 & _GEN_274 | _GEN_1005 | _GEN_963 & _GEN_146) & (_GEN_939 ? io_wb_resps_0_bits_predicated : ~_GEN_906 & rob_predicated_1_8));
    rob_predicated_1_9 <= ~(_GEN_1227 & _GEN_660 | _GEN_1204 | _GEN_1161 & _GEN_532) & (_GEN_1138 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_404 | _GEN_1072 | _GEN_1029 & _GEN_276 | _GEN_1006 | _GEN_963 & _GEN_148) & (_GEN_940 ? io_wb_resps_0_bits_predicated : ~_GEN_907 & rob_predicated_1_9));
    rob_predicated_1_10 <= ~(_GEN_1227 & _GEN_662 | _GEN_1205 | _GEN_1161 & _GEN_534) & (_GEN_1139 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_406 | _GEN_1073 | _GEN_1029 & _GEN_278 | _GEN_1007 | _GEN_963 & _GEN_150) & (_GEN_941 ? io_wb_resps_0_bits_predicated : ~_GEN_908 & rob_predicated_1_10));
    rob_predicated_1_11 <= ~(_GEN_1227 & _GEN_664 | _GEN_1206 | _GEN_1161 & _GEN_536) & (_GEN_1140 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_408 | _GEN_1074 | _GEN_1029 & _GEN_280 | _GEN_1008 | _GEN_963 & _GEN_152) & (_GEN_942 ? io_wb_resps_0_bits_predicated : ~_GEN_909 & rob_predicated_1_11));
    rob_predicated_1_12 <= ~(_GEN_1227 & _GEN_666 | _GEN_1207 | _GEN_1161 & _GEN_538) & (_GEN_1141 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_410 | _GEN_1075 | _GEN_1029 & _GEN_282 | _GEN_1009 | _GEN_963 & _GEN_154) & (_GEN_943 ? io_wb_resps_0_bits_predicated : ~_GEN_910 & rob_predicated_1_12));
    rob_predicated_1_13 <= ~(_GEN_1227 & _GEN_668 | _GEN_1208 | _GEN_1161 & _GEN_540) & (_GEN_1142 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_412 | _GEN_1076 | _GEN_1029 & _GEN_284 | _GEN_1010 | _GEN_963 & _GEN_156) & (_GEN_944 ? io_wb_resps_0_bits_predicated : ~_GEN_911 & rob_predicated_1_13));
    rob_predicated_1_14 <= ~(_GEN_1227 & _GEN_670 | _GEN_1209 | _GEN_1161 & _GEN_542) & (_GEN_1143 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_414 | _GEN_1077 | _GEN_1029 & _GEN_286 | _GEN_1011 | _GEN_963 & _GEN_158) & (_GEN_945 ? io_wb_resps_0_bits_predicated : ~_GEN_912 & rob_predicated_1_14));
    rob_predicated_1_15 <= ~(_GEN_1227 & _GEN_672 | _GEN_1210 | _GEN_1161 & _GEN_544) & (_GEN_1144 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_416 | _GEN_1078 | _GEN_1029 & _GEN_288 | _GEN_1012 | _GEN_963 & _GEN_160) & (_GEN_946 ? io_wb_resps_0_bits_predicated : ~_GEN_913 & rob_predicated_1_15));
    rob_predicated_1_16 <= ~(_GEN_1227 & _GEN_674 | _GEN_1211 | _GEN_1161 & _GEN_546) & (_GEN_1145 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_418 | _GEN_1079 | _GEN_1029 & _GEN_290 | _GEN_1013 | _GEN_963 & _GEN_162) & (_GEN_947 ? io_wb_resps_0_bits_predicated : ~_GEN_914 & rob_predicated_1_16));
    rob_predicated_1_17 <= ~(_GEN_1227 & _GEN_676 | _GEN_1212 | _GEN_1161 & _GEN_548) & (_GEN_1146 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_420 | _GEN_1080 | _GEN_1029 & _GEN_292 | _GEN_1014 | _GEN_963 & _GEN_164) & (_GEN_948 ? io_wb_resps_0_bits_predicated : ~_GEN_915 & rob_predicated_1_17));
    rob_predicated_1_18 <= ~(_GEN_1227 & _GEN_678 | _GEN_1213 | _GEN_1161 & _GEN_550) & (_GEN_1147 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_422 | _GEN_1081 | _GEN_1029 & _GEN_294 | _GEN_1015 | _GEN_963 & _GEN_166) & (_GEN_949 ? io_wb_resps_0_bits_predicated : ~_GEN_916 & rob_predicated_1_18));
    rob_predicated_1_19 <= ~(_GEN_1227 & _GEN_680 | _GEN_1214 | _GEN_1161 & _GEN_552) & (_GEN_1148 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_424 | _GEN_1082 | _GEN_1029 & _GEN_296 | _GEN_1016 | _GEN_963 & _GEN_168) & (_GEN_950 ? io_wb_resps_0_bits_predicated : ~_GEN_917 & rob_predicated_1_19));
    rob_predicated_1_20 <= ~(_GEN_1227 & _GEN_682 | _GEN_1215 | _GEN_1161 & _GEN_554) & (_GEN_1149 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_426 | _GEN_1083 | _GEN_1029 & _GEN_298 | _GEN_1017 | _GEN_963 & _GEN_170) & (_GEN_951 ? io_wb_resps_0_bits_predicated : ~_GEN_918 & rob_predicated_1_20));
    rob_predicated_1_21 <= ~(_GEN_1227 & _GEN_684 | _GEN_1216 | _GEN_1161 & _GEN_556) & (_GEN_1150 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_428 | _GEN_1084 | _GEN_1029 & _GEN_300 | _GEN_1018 | _GEN_963 & _GEN_172) & (_GEN_952 ? io_wb_resps_0_bits_predicated : ~_GEN_919 & rob_predicated_1_21));
    rob_predicated_1_22 <= ~(_GEN_1227 & _GEN_686 | _GEN_1217 | _GEN_1161 & _GEN_558) & (_GEN_1151 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_430 | _GEN_1085 | _GEN_1029 & _GEN_302 | _GEN_1019 | _GEN_963 & _GEN_174) & (_GEN_953 ? io_wb_resps_0_bits_predicated : ~_GEN_920 & rob_predicated_1_22));
    rob_predicated_1_23 <= ~(_GEN_1227 & _GEN_688 | _GEN_1218 | _GEN_1161 & _GEN_560) & (_GEN_1152 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_432 | _GEN_1086 | _GEN_1029 & _GEN_304 | _GEN_1020 | _GEN_963 & _GEN_176) & (_GEN_954 ? io_wb_resps_0_bits_predicated : ~_GEN_921 & rob_predicated_1_23));
    rob_predicated_1_24 <= ~(_GEN_1227 & _GEN_690 | _GEN_1219 | _GEN_1161 & _GEN_562) & (_GEN_1153 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_434 | _GEN_1087 | _GEN_1029 & _GEN_306 | _GEN_1021 | _GEN_963 & _GEN_178) & (_GEN_955 ? io_wb_resps_0_bits_predicated : ~_GEN_922 & rob_predicated_1_24));
    rob_predicated_1_25 <= ~(_GEN_1227 & _GEN_692 | _GEN_1220 | _GEN_1161 & _GEN_564) & (_GEN_1154 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_436 | _GEN_1088 | _GEN_1029 & _GEN_308 | _GEN_1022 | _GEN_963 & _GEN_180) & (_GEN_956 ? io_wb_resps_0_bits_predicated : ~_GEN_923 & rob_predicated_1_25));
    rob_predicated_1_26 <= ~(_GEN_1227 & _GEN_694 | _GEN_1221 | _GEN_1161 & _GEN_566) & (_GEN_1155 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_438 | _GEN_1089 | _GEN_1029 & _GEN_310 | _GEN_1023 | _GEN_963 & _GEN_182) & (_GEN_957 ? io_wb_resps_0_bits_predicated : ~_GEN_924 & rob_predicated_1_26));
    rob_predicated_1_27 <= ~(_GEN_1227 & _GEN_696 | _GEN_1222 | _GEN_1161 & _GEN_568) & (_GEN_1156 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_440 | _GEN_1090 | _GEN_1029 & _GEN_312 | _GEN_1024 | _GEN_963 & _GEN_184) & (_GEN_958 ? io_wb_resps_0_bits_predicated : ~_GEN_925 & rob_predicated_1_27));
    rob_predicated_1_28 <= ~(_GEN_1227 & _GEN_698 | _GEN_1223 | _GEN_1161 & _GEN_570) & (_GEN_1157 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_442 | _GEN_1091 | _GEN_1029 & _GEN_314 | _GEN_1025 | _GEN_963 & _GEN_186) & (_GEN_959 ? io_wb_resps_0_bits_predicated : ~_GEN_926 & rob_predicated_1_28));
    rob_predicated_1_29 <= ~(_GEN_1227 & _GEN_700 | _GEN_1224 | _GEN_1161 & _GEN_572) & (_GEN_1158 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_444 | _GEN_1092 | _GEN_1029 & _GEN_316 | _GEN_1026 | _GEN_963 & _GEN_188) & (_GEN_960 ? io_wb_resps_0_bits_predicated : ~_GEN_927 & rob_predicated_1_29));
    rob_predicated_1_30 <= ~(_GEN_1227 & _GEN_702 | _GEN_1225 | _GEN_1161 & _GEN_574) & (_GEN_1159 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & _GEN_446 | _GEN_1093 | _GEN_1029 & _GEN_318 | _GEN_1027 | _GEN_963 & _GEN_190) & (_GEN_961 ? io_wb_resps_0_bits_predicated : ~_GEN_928 & rob_predicated_1_30));
    rob_predicated_1_31 <= ~(_GEN_1227 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1226 | _GEN_1161 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_1160 ? io_wb_resps_6_bits_predicated : ~(_GEN_1095 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1094 | _GEN_1029 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1028 | _GEN_963 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_962 ? io_wb_resps_0_bits_predicated : ~_GEN_929 & rob_predicated_1_31));
    if (_GEN_1360) begin
      rob_uop_2_0_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_0_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_0_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_0_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_0_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_0_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_0_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_0_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_0_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_0_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_0_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_0_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_0_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_0_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_0_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_0_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2644) | ~rob_val_2_0) begin
      if (_GEN_1360)
        rob_uop_2_0_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_0_br_mask <= rob_uop_2_0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1361) begin
      rob_uop_2_1_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_1_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_1_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_1_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_1_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_1_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_1_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_1_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_1_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_1_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_1_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_1_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_1_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_1_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_1_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_1_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2645) | ~rob_val_2_1) begin
      if (_GEN_1361)
        rob_uop_2_1_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_1_br_mask <= rob_uop_2_1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1362) begin
      rob_uop_2_2_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_2_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_2_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_2_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_2_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_2_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_2_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_2_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_2_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_2_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_2_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_2_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_2_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_2_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_2_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_2_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2646) | ~rob_val_2_2) begin
      if (_GEN_1362)
        rob_uop_2_2_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_2_br_mask <= rob_uop_2_2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1363) begin
      rob_uop_2_3_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_3_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_3_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_3_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_3_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_3_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_3_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_3_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_3_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_3_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_3_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_3_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_3_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_3_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_3_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_3_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2647) | ~rob_val_2_3) begin
      if (_GEN_1363)
        rob_uop_2_3_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_3_br_mask <= rob_uop_2_3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1364) begin
      rob_uop_2_4_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_4_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_4_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_4_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_4_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_4_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_4_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_4_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_4_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_4_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_4_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_4_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_4_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_4_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_4_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_4_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2648) | ~rob_val_2_4) begin
      if (_GEN_1364)
        rob_uop_2_4_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_4_br_mask <= rob_uop_2_4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1365) begin
      rob_uop_2_5_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_5_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_5_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_5_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_5_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_5_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_5_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_5_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_5_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_5_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_5_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_5_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_5_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_5_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_5_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_5_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2649) | ~rob_val_2_5) begin
      if (_GEN_1365)
        rob_uop_2_5_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_5_br_mask <= rob_uop_2_5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1366) begin
      rob_uop_2_6_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_6_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_6_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_6_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_6_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_6_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_6_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_6_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_6_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_6_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_6_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_6_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_6_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_6_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_6_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_6_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2650) | ~rob_val_2_6) begin
      if (_GEN_1366)
        rob_uop_2_6_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_6_br_mask <= rob_uop_2_6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1367) begin
      rob_uop_2_7_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_7_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_7_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_7_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_7_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_7_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_7_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_7_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_7_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_7_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_7_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_7_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_7_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_7_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_7_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_7_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2651) | ~rob_val_2_7) begin
      if (_GEN_1367)
        rob_uop_2_7_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_7_br_mask <= rob_uop_2_7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1368) begin
      rob_uop_2_8_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_8_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_8_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_8_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_8_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_8_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_8_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_8_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_8_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_8_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_8_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_8_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_8_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_8_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_8_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_8_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2652) | ~rob_val_2_8) begin
      if (_GEN_1368)
        rob_uop_2_8_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_8_br_mask <= rob_uop_2_8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1369) begin
      rob_uop_2_9_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_9_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_9_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_9_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_9_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_9_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_9_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_9_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_9_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_9_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_9_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_9_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_9_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_9_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_9_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_9_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2653) | ~rob_val_2_9) begin
      if (_GEN_1369)
        rob_uop_2_9_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_9_br_mask <= rob_uop_2_9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1370) begin
      rob_uop_2_10_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_10_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_10_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_10_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_10_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_10_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_10_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_10_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_10_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_10_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_10_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_10_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_10_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_10_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_10_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_10_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2654) | ~rob_val_2_10) begin
      if (_GEN_1370)
        rob_uop_2_10_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_10_br_mask <= rob_uop_2_10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1371) begin
      rob_uop_2_11_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_11_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_11_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_11_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_11_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_11_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_11_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_11_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_11_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_11_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_11_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_11_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_11_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_11_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_11_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_11_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2655) | ~rob_val_2_11) begin
      if (_GEN_1371)
        rob_uop_2_11_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_11_br_mask <= rob_uop_2_11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1372) begin
      rob_uop_2_12_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_12_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_12_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_12_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_12_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_12_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_12_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_12_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_12_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_12_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_12_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_12_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_12_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_12_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_12_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_12_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2656) | ~rob_val_2_12) begin
      if (_GEN_1372)
        rob_uop_2_12_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_12_br_mask <= rob_uop_2_12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1373) begin
      rob_uop_2_13_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_13_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_13_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_13_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_13_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_13_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_13_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_13_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_13_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_13_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_13_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_13_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_13_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_13_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_13_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_13_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2657) | ~rob_val_2_13) begin
      if (_GEN_1373)
        rob_uop_2_13_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_13_br_mask <= rob_uop_2_13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1374) begin
      rob_uop_2_14_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_14_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_14_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_14_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_14_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_14_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_14_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_14_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_14_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_14_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_14_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_14_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_14_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_14_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_14_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_14_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2658) | ~rob_val_2_14) begin
      if (_GEN_1374)
        rob_uop_2_14_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_14_br_mask <= rob_uop_2_14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1375) begin
      rob_uop_2_15_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_15_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_15_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_15_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_15_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_15_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_15_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_15_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_15_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_15_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_15_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_15_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_15_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_15_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_15_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_15_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2659) | ~rob_val_2_15) begin
      if (_GEN_1375)
        rob_uop_2_15_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_15_br_mask <= rob_uop_2_15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1376) begin
      rob_uop_2_16_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_16_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_16_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_16_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_16_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_16_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_16_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_16_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_16_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_16_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_16_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_16_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_16_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_16_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_16_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_16_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2660) | ~rob_val_2_16) begin
      if (_GEN_1376)
        rob_uop_2_16_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_16_br_mask <= rob_uop_2_16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1377) begin
      rob_uop_2_17_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_17_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_17_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_17_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_17_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_17_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_17_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_17_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_17_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_17_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_17_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_17_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_17_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_17_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_17_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_17_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2661) | ~rob_val_2_17) begin
      if (_GEN_1377)
        rob_uop_2_17_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_17_br_mask <= rob_uop_2_17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1378) begin
      rob_uop_2_18_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_18_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_18_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_18_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_18_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_18_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_18_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_18_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_18_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_18_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_18_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_18_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_18_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_18_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_18_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_18_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2662) | ~rob_val_2_18) begin
      if (_GEN_1378)
        rob_uop_2_18_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_18_br_mask <= rob_uop_2_18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1379) begin
      rob_uop_2_19_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_19_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_19_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_19_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_19_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_19_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_19_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_19_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_19_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_19_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_19_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_19_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_19_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_19_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_19_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_19_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2663) | ~rob_val_2_19) begin
      if (_GEN_1379)
        rob_uop_2_19_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_19_br_mask <= rob_uop_2_19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1380) begin
      rob_uop_2_20_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_20_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_20_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_20_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_20_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_20_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_20_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_20_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_20_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_20_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_20_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_20_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_20_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_20_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_20_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_20_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2664) | ~rob_val_2_20) begin
      if (_GEN_1380)
        rob_uop_2_20_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_20_br_mask <= rob_uop_2_20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1381) begin
      rob_uop_2_21_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_21_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_21_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_21_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_21_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_21_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_21_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_21_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_21_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_21_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_21_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_21_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_21_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_21_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_21_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_21_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2665) | ~rob_val_2_21) begin
      if (_GEN_1381)
        rob_uop_2_21_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_21_br_mask <= rob_uop_2_21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1382) begin
      rob_uop_2_22_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_22_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_22_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_22_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_22_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_22_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_22_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_22_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_22_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_22_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_22_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_22_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_22_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_22_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_22_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_22_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2666) | ~rob_val_2_22) begin
      if (_GEN_1382)
        rob_uop_2_22_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_22_br_mask <= rob_uop_2_22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1383) begin
      rob_uop_2_23_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_23_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_23_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_23_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_23_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_23_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_23_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_23_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_23_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_23_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_23_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_23_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_23_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_23_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_23_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_23_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2667) | ~rob_val_2_23) begin
      if (_GEN_1383)
        rob_uop_2_23_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_23_br_mask <= rob_uop_2_23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1384) begin
      rob_uop_2_24_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_24_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_24_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_24_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_24_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_24_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_24_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_24_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_24_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_24_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_24_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_24_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_24_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_24_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_24_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_24_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2668) | ~rob_val_2_24) begin
      if (_GEN_1384)
        rob_uop_2_24_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_24_br_mask <= rob_uop_2_24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1385) begin
      rob_uop_2_25_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_25_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_25_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_25_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_25_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_25_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_25_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_25_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_25_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_25_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_25_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_25_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_25_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_25_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_25_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_25_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2669) | ~rob_val_2_25) begin
      if (_GEN_1385)
        rob_uop_2_25_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_25_br_mask <= rob_uop_2_25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1386) begin
      rob_uop_2_26_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_26_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_26_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_26_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_26_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_26_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_26_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_26_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_26_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_26_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_26_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_26_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_26_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_26_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_26_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_26_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2670) | ~rob_val_2_26) begin
      if (_GEN_1386)
        rob_uop_2_26_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_26_br_mask <= rob_uop_2_26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1387) begin
      rob_uop_2_27_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_27_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_27_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_27_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_27_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_27_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_27_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_27_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_27_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_27_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_27_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_27_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_27_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_27_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_27_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_27_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2671) | ~rob_val_2_27) begin
      if (_GEN_1387)
        rob_uop_2_27_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_27_br_mask <= rob_uop_2_27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1388) begin
      rob_uop_2_28_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_28_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_28_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_28_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_28_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_28_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_28_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_28_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_28_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_28_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_28_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_28_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_28_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_28_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_28_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_28_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2672) | ~rob_val_2_28) begin
      if (_GEN_1388)
        rob_uop_2_28_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_28_br_mask <= rob_uop_2_28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1389) begin
      rob_uop_2_29_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_29_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_29_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_29_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_29_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_29_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_29_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_29_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_29_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_29_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_29_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_29_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_29_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_29_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_29_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_29_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2673) | ~rob_val_2_29) begin
      if (_GEN_1389)
        rob_uop_2_29_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_29_br_mask <= rob_uop_2_29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1390) begin
      rob_uop_2_30_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_30_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_30_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_30_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_30_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_30_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_30_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_30_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_30_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_30_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_30_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_30_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_30_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_30_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_30_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_30_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2674) | ~rob_val_2_30) begin
      if (_GEN_1390)
        rob_uop_2_30_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_30_br_mask <= rob_uop_2_30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1391) begin
      rob_uop_2_31_uopc <= io_enq_uops_2_uopc;
      rob_uop_2_31_is_rvc <= io_enq_uops_2_is_rvc;
      rob_uop_2_31_ftq_idx <= io_enq_uops_2_ftq_idx;
      rob_uop_2_31_edge_inst <= io_enq_uops_2_edge_inst;
      rob_uop_2_31_pc_lob <= io_enq_uops_2_pc_lob;
      rob_uop_2_31_pdst <= io_enq_uops_2_pdst;
      rob_uop_2_31_stale_pdst <= io_enq_uops_2_stale_pdst;
      rob_uop_2_31_is_fencei <= io_enq_uops_2_is_fencei;
      rob_uop_2_31_uses_ldq <= io_enq_uops_2_uses_ldq;
      rob_uop_2_31_uses_stq <= io_enq_uops_2_uses_stq;
      rob_uop_2_31_is_sys_pc2epc <= io_enq_uops_2_is_sys_pc2epc;
      rob_uop_2_31_flush_on_commit <= io_enq_uops_2_flush_on_commit;
      rob_uop_2_31_ldst <= io_enq_uops_2_ldst;
      rob_uop_2_31_ldst_val <= io_enq_uops_2_ldst_val;
      rob_uop_2_31_dst_rtype <= io_enq_uops_2_dst_rtype;
      rob_uop_2_31_fp_val <= io_enq_uops_2_fp_val;
    end
    if ((|_GEN_2675) | ~rob_val_2_31) begin
      if (_GEN_1391)
        rob_uop_2_31_br_mask <= io_enq_uops_2_br_mask;
    end
    else
      rob_uop_2_31_br_mask <= rob_uop_2_31_br_mask & ~io_brupdate_b1_resolve_mask;
    rob_predicated_2_0 <= ~(_GEN_1689 & _GEN_642 | _GEN_1657 | _GEN_1623 & _GEN_514) & (_GEN_1591 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_386 | _GEN_1525 | _GEN_1491 & _GEN_258 | _GEN_1459 | _GEN_1425 & _GEN_130) & (_GEN_1393 ? io_wb_resps_0_bits_predicated : ~_GEN_1360 & rob_predicated_2_0));
    rob_predicated_2_1 <= ~(_GEN_1689 & _GEN_644 | _GEN_1658 | _GEN_1623 & _GEN_516) & (_GEN_1592 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_388 | _GEN_1526 | _GEN_1491 & _GEN_260 | _GEN_1460 | _GEN_1425 & _GEN_132) & (_GEN_1394 ? io_wb_resps_0_bits_predicated : ~_GEN_1361 & rob_predicated_2_1));
    rob_predicated_2_2 <= ~(_GEN_1689 & _GEN_646 | _GEN_1659 | _GEN_1623 & _GEN_518) & (_GEN_1593 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_390 | _GEN_1527 | _GEN_1491 & _GEN_262 | _GEN_1461 | _GEN_1425 & _GEN_134) & (_GEN_1395 ? io_wb_resps_0_bits_predicated : ~_GEN_1362 & rob_predicated_2_2));
    rob_predicated_2_3 <= ~(_GEN_1689 & _GEN_648 | _GEN_1660 | _GEN_1623 & _GEN_520) & (_GEN_1594 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_392 | _GEN_1528 | _GEN_1491 & _GEN_264 | _GEN_1462 | _GEN_1425 & _GEN_136) & (_GEN_1396 ? io_wb_resps_0_bits_predicated : ~_GEN_1363 & rob_predicated_2_3));
    rob_predicated_2_4 <= ~(_GEN_1689 & _GEN_650 | _GEN_1661 | _GEN_1623 & _GEN_522) & (_GEN_1595 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_394 | _GEN_1529 | _GEN_1491 & _GEN_266 | _GEN_1463 | _GEN_1425 & _GEN_138) & (_GEN_1397 ? io_wb_resps_0_bits_predicated : ~_GEN_1364 & rob_predicated_2_4));
    rob_predicated_2_5 <= ~(_GEN_1689 & _GEN_652 | _GEN_1662 | _GEN_1623 & _GEN_524) & (_GEN_1596 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_396 | _GEN_1530 | _GEN_1491 & _GEN_268 | _GEN_1464 | _GEN_1425 & _GEN_140) & (_GEN_1398 ? io_wb_resps_0_bits_predicated : ~_GEN_1365 & rob_predicated_2_5));
    rob_predicated_2_6 <= ~(_GEN_1689 & _GEN_654 | _GEN_1663 | _GEN_1623 & _GEN_526) & (_GEN_1597 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_398 | _GEN_1531 | _GEN_1491 & _GEN_270 | _GEN_1465 | _GEN_1425 & _GEN_142) & (_GEN_1399 ? io_wb_resps_0_bits_predicated : ~_GEN_1366 & rob_predicated_2_6));
    rob_predicated_2_7 <= ~(_GEN_1689 & _GEN_656 | _GEN_1664 | _GEN_1623 & _GEN_528) & (_GEN_1598 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_400 | _GEN_1532 | _GEN_1491 & _GEN_272 | _GEN_1466 | _GEN_1425 & _GEN_144) & (_GEN_1400 ? io_wb_resps_0_bits_predicated : ~_GEN_1367 & rob_predicated_2_7));
    rob_predicated_2_8 <= ~(_GEN_1689 & _GEN_658 | _GEN_1665 | _GEN_1623 & _GEN_530) & (_GEN_1599 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_402 | _GEN_1533 | _GEN_1491 & _GEN_274 | _GEN_1467 | _GEN_1425 & _GEN_146) & (_GEN_1401 ? io_wb_resps_0_bits_predicated : ~_GEN_1368 & rob_predicated_2_8));
    rob_predicated_2_9 <= ~(_GEN_1689 & _GEN_660 | _GEN_1666 | _GEN_1623 & _GEN_532) & (_GEN_1600 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_404 | _GEN_1534 | _GEN_1491 & _GEN_276 | _GEN_1468 | _GEN_1425 & _GEN_148) & (_GEN_1402 ? io_wb_resps_0_bits_predicated : ~_GEN_1369 & rob_predicated_2_9));
    rob_predicated_2_10 <= ~(_GEN_1689 & _GEN_662 | _GEN_1667 | _GEN_1623 & _GEN_534) & (_GEN_1601 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_406 | _GEN_1535 | _GEN_1491 & _GEN_278 | _GEN_1469 | _GEN_1425 & _GEN_150) & (_GEN_1403 ? io_wb_resps_0_bits_predicated : ~_GEN_1370 & rob_predicated_2_10));
    rob_predicated_2_11 <= ~(_GEN_1689 & _GEN_664 | _GEN_1668 | _GEN_1623 & _GEN_536) & (_GEN_1602 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_408 | _GEN_1536 | _GEN_1491 & _GEN_280 | _GEN_1470 | _GEN_1425 & _GEN_152) & (_GEN_1404 ? io_wb_resps_0_bits_predicated : ~_GEN_1371 & rob_predicated_2_11));
    rob_predicated_2_12 <= ~(_GEN_1689 & _GEN_666 | _GEN_1669 | _GEN_1623 & _GEN_538) & (_GEN_1603 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_410 | _GEN_1537 | _GEN_1491 & _GEN_282 | _GEN_1471 | _GEN_1425 & _GEN_154) & (_GEN_1405 ? io_wb_resps_0_bits_predicated : ~_GEN_1372 & rob_predicated_2_12));
    rob_predicated_2_13 <= ~(_GEN_1689 & _GEN_668 | _GEN_1670 | _GEN_1623 & _GEN_540) & (_GEN_1604 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_412 | _GEN_1538 | _GEN_1491 & _GEN_284 | _GEN_1472 | _GEN_1425 & _GEN_156) & (_GEN_1406 ? io_wb_resps_0_bits_predicated : ~_GEN_1373 & rob_predicated_2_13));
    rob_predicated_2_14 <= ~(_GEN_1689 & _GEN_670 | _GEN_1671 | _GEN_1623 & _GEN_542) & (_GEN_1605 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_414 | _GEN_1539 | _GEN_1491 & _GEN_286 | _GEN_1473 | _GEN_1425 & _GEN_158) & (_GEN_1407 ? io_wb_resps_0_bits_predicated : ~_GEN_1374 & rob_predicated_2_14));
    rob_predicated_2_15 <= ~(_GEN_1689 & _GEN_672 | _GEN_1672 | _GEN_1623 & _GEN_544) & (_GEN_1606 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_416 | _GEN_1540 | _GEN_1491 & _GEN_288 | _GEN_1474 | _GEN_1425 & _GEN_160) & (_GEN_1408 ? io_wb_resps_0_bits_predicated : ~_GEN_1375 & rob_predicated_2_15));
    rob_predicated_2_16 <= ~(_GEN_1689 & _GEN_674 | _GEN_1673 | _GEN_1623 & _GEN_546) & (_GEN_1607 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_418 | _GEN_1541 | _GEN_1491 & _GEN_290 | _GEN_1475 | _GEN_1425 & _GEN_162) & (_GEN_1409 ? io_wb_resps_0_bits_predicated : ~_GEN_1376 & rob_predicated_2_16));
    rob_predicated_2_17 <= ~(_GEN_1689 & _GEN_676 | _GEN_1674 | _GEN_1623 & _GEN_548) & (_GEN_1608 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_420 | _GEN_1542 | _GEN_1491 & _GEN_292 | _GEN_1476 | _GEN_1425 & _GEN_164) & (_GEN_1410 ? io_wb_resps_0_bits_predicated : ~_GEN_1377 & rob_predicated_2_17));
    rob_predicated_2_18 <= ~(_GEN_1689 & _GEN_678 | _GEN_1675 | _GEN_1623 & _GEN_550) & (_GEN_1609 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_422 | _GEN_1543 | _GEN_1491 & _GEN_294 | _GEN_1477 | _GEN_1425 & _GEN_166) & (_GEN_1411 ? io_wb_resps_0_bits_predicated : ~_GEN_1378 & rob_predicated_2_18));
    rob_predicated_2_19 <= ~(_GEN_1689 & _GEN_680 | _GEN_1676 | _GEN_1623 & _GEN_552) & (_GEN_1610 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_424 | _GEN_1544 | _GEN_1491 & _GEN_296 | _GEN_1478 | _GEN_1425 & _GEN_168) & (_GEN_1412 ? io_wb_resps_0_bits_predicated : ~_GEN_1379 & rob_predicated_2_19));
    rob_predicated_2_20 <= ~(_GEN_1689 & _GEN_682 | _GEN_1677 | _GEN_1623 & _GEN_554) & (_GEN_1611 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_426 | _GEN_1545 | _GEN_1491 & _GEN_298 | _GEN_1479 | _GEN_1425 & _GEN_170) & (_GEN_1413 ? io_wb_resps_0_bits_predicated : ~_GEN_1380 & rob_predicated_2_20));
    rob_predicated_2_21 <= ~(_GEN_1689 & _GEN_684 | _GEN_1678 | _GEN_1623 & _GEN_556) & (_GEN_1612 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_428 | _GEN_1546 | _GEN_1491 & _GEN_300 | _GEN_1480 | _GEN_1425 & _GEN_172) & (_GEN_1414 ? io_wb_resps_0_bits_predicated : ~_GEN_1381 & rob_predicated_2_21));
    rob_predicated_2_22 <= ~(_GEN_1689 & _GEN_686 | _GEN_1679 | _GEN_1623 & _GEN_558) & (_GEN_1613 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_430 | _GEN_1547 | _GEN_1491 & _GEN_302 | _GEN_1481 | _GEN_1425 & _GEN_174) & (_GEN_1415 ? io_wb_resps_0_bits_predicated : ~_GEN_1382 & rob_predicated_2_22));
    rob_predicated_2_23 <= ~(_GEN_1689 & _GEN_688 | _GEN_1680 | _GEN_1623 & _GEN_560) & (_GEN_1614 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_432 | _GEN_1548 | _GEN_1491 & _GEN_304 | _GEN_1482 | _GEN_1425 & _GEN_176) & (_GEN_1416 ? io_wb_resps_0_bits_predicated : ~_GEN_1383 & rob_predicated_2_23));
    rob_predicated_2_24 <= ~(_GEN_1689 & _GEN_690 | _GEN_1681 | _GEN_1623 & _GEN_562) & (_GEN_1615 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_434 | _GEN_1549 | _GEN_1491 & _GEN_306 | _GEN_1483 | _GEN_1425 & _GEN_178) & (_GEN_1417 ? io_wb_resps_0_bits_predicated : ~_GEN_1384 & rob_predicated_2_24));
    rob_predicated_2_25 <= ~(_GEN_1689 & _GEN_692 | _GEN_1682 | _GEN_1623 & _GEN_564) & (_GEN_1616 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_436 | _GEN_1550 | _GEN_1491 & _GEN_308 | _GEN_1484 | _GEN_1425 & _GEN_180) & (_GEN_1418 ? io_wb_resps_0_bits_predicated : ~_GEN_1385 & rob_predicated_2_25));
    rob_predicated_2_26 <= ~(_GEN_1689 & _GEN_694 | _GEN_1683 | _GEN_1623 & _GEN_566) & (_GEN_1617 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_438 | _GEN_1551 | _GEN_1491 & _GEN_310 | _GEN_1485 | _GEN_1425 & _GEN_182) & (_GEN_1419 ? io_wb_resps_0_bits_predicated : ~_GEN_1386 & rob_predicated_2_26));
    rob_predicated_2_27 <= ~(_GEN_1689 & _GEN_696 | _GEN_1684 | _GEN_1623 & _GEN_568) & (_GEN_1618 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_440 | _GEN_1552 | _GEN_1491 & _GEN_312 | _GEN_1486 | _GEN_1425 & _GEN_184) & (_GEN_1420 ? io_wb_resps_0_bits_predicated : ~_GEN_1387 & rob_predicated_2_27));
    rob_predicated_2_28 <= ~(_GEN_1689 & _GEN_698 | _GEN_1685 | _GEN_1623 & _GEN_570) & (_GEN_1619 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_442 | _GEN_1553 | _GEN_1491 & _GEN_314 | _GEN_1487 | _GEN_1425 & _GEN_186) & (_GEN_1421 ? io_wb_resps_0_bits_predicated : ~_GEN_1388 & rob_predicated_2_28));
    rob_predicated_2_29 <= ~(_GEN_1689 & _GEN_700 | _GEN_1686 | _GEN_1623 & _GEN_572) & (_GEN_1620 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_444 | _GEN_1554 | _GEN_1491 & _GEN_316 | _GEN_1488 | _GEN_1425 & _GEN_188) & (_GEN_1422 ? io_wb_resps_0_bits_predicated : ~_GEN_1389 & rob_predicated_2_29));
    rob_predicated_2_30 <= ~(_GEN_1689 & _GEN_702 | _GEN_1687 | _GEN_1623 & _GEN_574) & (_GEN_1621 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & _GEN_446 | _GEN_1555 | _GEN_1491 & _GEN_318 | _GEN_1489 | _GEN_1425 & _GEN_190) & (_GEN_1423 ? io_wb_resps_0_bits_predicated : ~_GEN_1390 & rob_predicated_2_30));
    rob_predicated_2_31 <= ~(_GEN_1689 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_1688 | _GEN_1623 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_1622 ? io_wb_resps_6_bits_predicated : ~(_GEN_1557 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_1556 | _GEN_1491 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1490 | _GEN_1425 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_1424 ? io_wb_resps_0_bits_predicated : ~_GEN_1391 & rob_predicated_2_31));
    if (_GEN_1822) begin
      rob_uop_3_0_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_0_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_0_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_0_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_0_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_0_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_0_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_0_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_0_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_0_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_0_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_0_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_0_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_0_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_0_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_0_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2711) | ~rob_val_3_0) begin
      if (_GEN_1822)
        rob_uop_3_0_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_0_br_mask <= rob_uop_3_0_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1823) begin
      rob_uop_3_1_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_1_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_1_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_1_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_1_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_1_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_1_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_1_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_1_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_1_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_1_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_1_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_1_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_1_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_1_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_1_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2712) | ~rob_val_3_1) begin
      if (_GEN_1823)
        rob_uop_3_1_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_1_br_mask <= rob_uop_3_1_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1824) begin
      rob_uop_3_2_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_2_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_2_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_2_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_2_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_2_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_2_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_2_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_2_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_2_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_2_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_2_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_2_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_2_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_2_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_2_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2713) | ~rob_val_3_2) begin
      if (_GEN_1824)
        rob_uop_3_2_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_2_br_mask <= rob_uop_3_2_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1825) begin
      rob_uop_3_3_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_3_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_3_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_3_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_3_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_3_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_3_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_3_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_3_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_3_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_3_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_3_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_3_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_3_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_3_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_3_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2714) | ~rob_val_3_3) begin
      if (_GEN_1825)
        rob_uop_3_3_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_3_br_mask <= rob_uop_3_3_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1826) begin
      rob_uop_3_4_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_4_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_4_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_4_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_4_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_4_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_4_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_4_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_4_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_4_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_4_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_4_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_4_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_4_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_4_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_4_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2715) | ~rob_val_3_4) begin
      if (_GEN_1826)
        rob_uop_3_4_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_4_br_mask <= rob_uop_3_4_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1827) begin
      rob_uop_3_5_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_5_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_5_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_5_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_5_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_5_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_5_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_5_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_5_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_5_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_5_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_5_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_5_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_5_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_5_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_5_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2716) | ~rob_val_3_5) begin
      if (_GEN_1827)
        rob_uop_3_5_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_5_br_mask <= rob_uop_3_5_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1828) begin
      rob_uop_3_6_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_6_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_6_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_6_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_6_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_6_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_6_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_6_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_6_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_6_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_6_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_6_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_6_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_6_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_6_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_6_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2717) | ~rob_val_3_6) begin
      if (_GEN_1828)
        rob_uop_3_6_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_6_br_mask <= rob_uop_3_6_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1829) begin
      rob_uop_3_7_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_7_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_7_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_7_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_7_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_7_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_7_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_7_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_7_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_7_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_7_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_7_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_7_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_7_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_7_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_7_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2718) | ~rob_val_3_7) begin
      if (_GEN_1829)
        rob_uop_3_7_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_7_br_mask <= rob_uop_3_7_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1830) begin
      rob_uop_3_8_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_8_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_8_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_8_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_8_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_8_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_8_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_8_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_8_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_8_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_8_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_8_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_8_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_8_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_8_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_8_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2719) | ~rob_val_3_8) begin
      if (_GEN_1830)
        rob_uop_3_8_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_8_br_mask <= rob_uop_3_8_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1831) begin
      rob_uop_3_9_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_9_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_9_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_9_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_9_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_9_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_9_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_9_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_9_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_9_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_9_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_9_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_9_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_9_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_9_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_9_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2720) | ~rob_val_3_9) begin
      if (_GEN_1831)
        rob_uop_3_9_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_9_br_mask <= rob_uop_3_9_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1832) begin
      rob_uop_3_10_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_10_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_10_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_10_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_10_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_10_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_10_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_10_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_10_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_10_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_10_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_10_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_10_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_10_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_10_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_10_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2721) | ~rob_val_3_10) begin
      if (_GEN_1832)
        rob_uop_3_10_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_10_br_mask <= rob_uop_3_10_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1833) begin
      rob_uop_3_11_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_11_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_11_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_11_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_11_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_11_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_11_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_11_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_11_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_11_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_11_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_11_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_11_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_11_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_11_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_11_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2722) | ~rob_val_3_11) begin
      if (_GEN_1833)
        rob_uop_3_11_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_11_br_mask <= rob_uop_3_11_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1834) begin
      rob_uop_3_12_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_12_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_12_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_12_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_12_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_12_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_12_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_12_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_12_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_12_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_12_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_12_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_12_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_12_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_12_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_12_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2723) | ~rob_val_3_12) begin
      if (_GEN_1834)
        rob_uop_3_12_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_12_br_mask <= rob_uop_3_12_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1835) begin
      rob_uop_3_13_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_13_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_13_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_13_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_13_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_13_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_13_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_13_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_13_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_13_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_13_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_13_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_13_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_13_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_13_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_13_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2724) | ~rob_val_3_13) begin
      if (_GEN_1835)
        rob_uop_3_13_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_13_br_mask <= rob_uop_3_13_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1836) begin
      rob_uop_3_14_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_14_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_14_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_14_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_14_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_14_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_14_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_14_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_14_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_14_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_14_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_14_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_14_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_14_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_14_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_14_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2725) | ~rob_val_3_14) begin
      if (_GEN_1836)
        rob_uop_3_14_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_14_br_mask <= rob_uop_3_14_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1837) begin
      rob_uop_3_15_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_15_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_15_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_15_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_15_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_15_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_15_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_15_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_15_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_15_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_15_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_15_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_15_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_15_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_15_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_15_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2726) | ~rob_val_3_15) begin
      if (_GEN_1837)
        rob_uop_3_15_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_15_br_mask <= rob_uop_3_15_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1838) begin
      rob_uop_3_16_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_16_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_16_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_16_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_16_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_16_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_16_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_16_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_16_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_16_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_16_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_16_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_16_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_16_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_16_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_16_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2727) | ~rob_val_3_16) begin
      if (_GEN_1838)
        rob_uop_3_16_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_16_br_mask <= rob_uop_3_16_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1839) begin
      rob_uop_3_17_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_17_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_17_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_17_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_17_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_17_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_17_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_17_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_17_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_17_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_17_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_17_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_17_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_17_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_17_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_17_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2728) | ~rob_val_3_17) begin
      if (_GEN_1839)
        rob_uop_3_17_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_17_br_mask <= rob_uop_3_17_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1840) begin
      rob_uop_3_18_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_18_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_18_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_18_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_18_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_18_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_18_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_18_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_18_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_18_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_18_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_18_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_18_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_18_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_18_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_18_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2729) | ~rob_val_3_18) begin
      if (_GEN_1840)
        rob_uop_3_18_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_18_br_mask <= rob_uop_3_18_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1841) begin
      rob_uop_3_19_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_19_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_19_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_19_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_19_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_19_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_19_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_19_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_19_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_19_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_19_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_19_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_19_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_19_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_19_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_19_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2730) | ~rob_val_3_19) begin
      if (_GEN_1841)
        rob_uop_3_19_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_19_br_mask <= rob_uop_3_19_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1842) begin
      rob_uop_3_20_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_20_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_20_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_20_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_20_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_20_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_20_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_20_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_20_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_20_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_20_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_20_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_20_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_20_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_20_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_20_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2731) | ~rob_val_3_20) begin
      if (_GEN_1842)
        rob_uop_3_20_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_20_br_mask <= rob_uop_3_20_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1843) begin
      rob_uop_3_21_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_21_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_21_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_21_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_21_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_21_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_21_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_21_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_21_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_21_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_21_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_21_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_21_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_21_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_21_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_21_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2732) | ~rob_val_3_21) begin
      if (_GEN_1843)
        rob_uop_3_21_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_21_br_mask <= rob_uop_3_21_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1844) begin
      rob_uop_3_22_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_22_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_22_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_22_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_22_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_22_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_22_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_22_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_22_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_22_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_22_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_22_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_22_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_22_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_22_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_22_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2733) | ~rob_val_3_22) begin
      if (_GEN_1844)
        rob_uop_3_22_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_22_br_mask <= rob_uop_3_22_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1845) begin
      rob_uop_3_23_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_23_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_23_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_23_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_23_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_23_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_23_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_23_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_23_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_23_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_23_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_23_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_23_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_23_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_23_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_23_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2734) | ~rob_val_3_23) begin
      if (_GEN_1845)
        rob_uop_3_23_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_23_br_mask <= rob_uop_3_23_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1846) begin
      rob_uop_3_24_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_24_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_24_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_24_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_24_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_24_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_24_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_24_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_24_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_24_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_24_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_24_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_24_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_24_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_24_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_24_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2735) | ~rob_val_3_24) begin
      if (_GEN_1846)
        rob_uop_3_24_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_24_br_mask <= rob_uop_3_24_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1847) begin
      rob_uop_3_25_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_25_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_25_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_25_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_25_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_25_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_25_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_25_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_25_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_25_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_25_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_25_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_25_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_25_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_25_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_25_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2736) | ~rob_val_3_25) begin
      if (_GEN_1847)
        rob_uop_3_25_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_25_br_mask <= rob_uop_3_25_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1848) begin
      rob_uop_3_26_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_26_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_26_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_26_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_26_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_26_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_26_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_26_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_26_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_26_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_26_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_26_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_26_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_26_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_26_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_26_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2737) | ~rob_val_3_26) begin
      if (_GEN_1848)
        rob_uop_3_26_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_26_br_mask <= rob_uop_3_26_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1849) begin
      rob_uop_3_27_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_27_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_27_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_27_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_27_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_27_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_27_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_27_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_27_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_27_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_27_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_27_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_27_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_27_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_27_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_27_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2738) | ~rob_val_3_27) begin
      if (_GEN_1849)
        rob_uop_3_27_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_27_br_mask <= rob_uop_3_27_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1850) begin
      rob_uop_3_28_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_28_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_28_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_28_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_28_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_28_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_28_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_28_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_28_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_28_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_28_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_28_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_28_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_28_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_28_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_28_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2739) | ~rob_val_3_28) begin
      if (_GEN_1850)
        rob_uop_3_28_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_28_br_mask <= rob_uop_3_28_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1851) begin
      rob_uop_3_29_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_29_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_29_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_29_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_29_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_29_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_29_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_29_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_29_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_29_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_29_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_29_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_29_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_29_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_29_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_29_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2740) | ~rob_val_3_29) begin
      if (_GEN_1851)
        rob_uop_3_29_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_29_br_mask <= rob_uop_3_29_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1852) begin
      rob_uop_3_30_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_30_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_30_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_30_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_30_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_30_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_30_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_30_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_30_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_30_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_30_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_30_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_30_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_30_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_30_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_30_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2741) | ~rob_val_3_30) begin
      if (_GEN_1852)
        rob_uop_3_30_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_30_br_mask <= rob_uop_3_30_br_mask & ~io_brupdate_b1_resolve_mask;
    if (_GEN_1853) begin
      rob_uop_3_31_uopc <= io_enq_uops_3_uopc;
      rob_uop_3_31_is_rvc <= io_enq_uops_3_is_rvc;
      rob_uop_3_31_ftq_idx <= io_enq_uops_3_ftq_idx;
      rob_uop_3_31_edge_inst <= io_enq_uops_3_edge_inst;
      rob_uop_3_31_pc_lob <= io_enq_uops_3_pc_lob;
      rob_uop_3_31_pdst <= io_enq_uops_3_pdst;
      rob_uop_3_31_stale_pdst <= io_enq_uops_3_stale_pdst;
      rob_uop_3_31_is_fencei <= io_enq_uops_3_is_fencei;
      rob_uop_3_31_uses_ldq <= io_enq_uops_3_uses_ldq;
      rob_uop_3_31_uses_stq <= io_enq_uops_3_uses_stq;
      rob_uop_3_31_is_sys_pc2epc <= io_enq_uops_3_is_sys_pc2epc;
      rob_uop_3_31_flush_on_commit <= io_enq_uops_3_flush_on_commit;
      rob_uop_3_31_ldst <= io_enq_uops_3_ldst;
      rob_uop_3_31_ldst_val <= io_enq_uops_3_ldst_val;
      rob_uop_3_31_dst_rtype <= io_enq_uops_3_dst_rtype;
      rob_uop_3_31_fp_val <= io_enq_uops_3_fp_val;
    end
    if ((|_GEN_2742) | ~rob_val_3_31) begin
      if (_GEN_1853)
        rob_uop_3_31_br_mask <= io_enq_uops_3_br_mask;
    end
    else
      rob_uop_3_31_br_mask <= rob_uop_3_31_br_mask & ~io_brupdate_b1_resolve_mask;
    rob_predicated_3_0 <= ~(_GEN_2151 & _GEN_642 | _GEN_2119 | _GEN_2085 & _GEN_514) & (_GEN_2053 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_386 | _GEN_1987 | _GEN_1953 & _GEN_258 | _GEN_1921 | _GEN_1887 & _GEN_130) & (_GEN_1855 ? io_wb_resps_0_bits_predicated : ~_GEN_1822 & rob_predicated_3_0));
    rob_predicated_3_1 <= ~(_GEN_2151 & _GEN_644 | _GEN_2120 | _GEN_2085 & _GEN_516) & (_GEN_2054 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_388 | _GEN_1988 | _GEN_1953 & _GEN_260 | _GEN_1922 | _GEN_1887 & _GEN_132) & (_GEN_1856 ? io_wb_resps_0_bits_predicated : ~_GEN_1823 & rob_predicated_3_1));
    rob_predicated_3_2 <= ~(_GEN_2151 & _GEN_646 | _GEN_2121 | _GEN_2085 & _GEN_518) & (_GEN_2055 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_390 | _GEN_1989 | _GEN_1953 & _GEN_262 | _GEN_1923 | _GEN_1887 & _GEN_134) & (_GEN_1857 ? io_wb_resps_0_bits_predicated : ~_GEN_1824 & rob_predicated_3_2));
    rob_predicated_3_3 <= ~(_GEN_2151 & _GEN_648 | _GEN_2122 | _GEN_2085 & _GEN_520) & (_GEN_2056 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_392 | _GEN_1990 | _GEN_1953 & _GEN_264 | _GEN_1924 | _GEN_1887 & _GEN_136) & (_GEN_1858 ? io_wb_resps_0_bits_predicated : ~_GEN_1825 & rob_predicated_3_3));
    rob_predicated_3_4 <= ~(_GEN_2151 & _GEN_650 | _GEN_2123 | _GEN_2085 & _GEN_522) & (_GEN_2057 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_394 | _GEN_1991 | _GEN_1953 & _GEN_266 | _GEN_1925 | _GEN_1887 & _GEN_138) & (_GEN_1859 ? io_wb_resps_0_bits_predicated : ~_GEN_1826 & rob_predicated_3_4));
    rob_predicated_3_5 <= ~(_GEN_2151 & _GEN_652 | _GEN_2124 | _GEN_2085 & _GEN_524) & (_GEN_2058 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_396 | _GEN_1992 | _GEN_1953 & _GEN_268 | _GEN_1926 | _GEN_1887 & _GEN_140) & (_GEN_1860 ? io_wb_resps_0_bits_predicated : ~_GEN_1827 & rob_predicated_3_5));
    rob_predicated_3_6 <= ~(_GEN_2151 & _GEN_654 | _GEN_2125 | _GEN_2085 & _GEN_526) & (_GEN_2059 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_398 | _GEN_1993 | _GEN_1953 & _GEN_270 | _GEN_1927 | _GEN_1887 & _GEN_142) & (_GEN_1861 ? io_wb_resps_0_bits_predicated : ~_GEN_1828 & rob_predicated_3_6));
    rob_predicated_3_7 <= ~(_GEN_2151 & _GEN_656 | _GEN_2126 | _GEN_2085 & _GEN_528) & (_GEN_2060 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_400 | _GEN_1994 | _GEN_1953 & _GEN_272 | _GEN_1928 | _GEN_1887 & _GEN_144) & (_GEN_1862 ? io_wb_resps_0_bits_predicated : ~_GEN_1829 & rob_predicated_3_7));
    rob_predicated_3_8 <= ~(_GEN_2151 & _GEN_658 | _GEN_2127 | _GEN_2085 & _GEN_530) & (_GEN_2061 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_402 | _GEN_1995 | _GEN_1953 & _GEN_274 | _GEN_1929 | _GEN_1887 & _GEN_146) & (_GEN_1863 ? io_wb_resps_0_bits_predicated : ~_GEN_1830 & rob_predicated_3_8));
    rob_predicated_3_9 <= ~(_GEN_2151 & _GEN_660 | _GEN_2128 | _GEN_2085 & _GEN_532) & (_GEN_2062 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_404 | _GEN_1996 | _GEN_1953 & _GEN_276 | _GEN_1930 | _GEN_1887 & _GEN_148) & (_GEN_1864 ? io_wb_resps_0_bits_predicated : ~_GEN_1831 & rob_predicated_3_9));
    rob_predicated_3_10 <= ~(_GEN_2151 & _GEN_662 | _GEN_2129 | _GEN_2085 & _GEN_534) & (_GEN_2063 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_406 | _GEN_1997 | _GEN_1953 & _GEN_278 | _GEN_1931 | _GEN_1887 & _GEN_150) & (_GEN_1865 ? io_wb_resps_0_bits_predicated : ~_GEN_1832 & rob_predicated_3_10));
    rob_predicated_3_11 <= ~(_GEN_2151 & _GEN_664 | _GEN_2130 | _GEN_2085 & _GEN_536) & (_GEN_2064 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_408 | _GEN_1998 | _GEN_1953 & _GEN_280 | _GEN_1932 | _GEN_1887 & _GEN_152) & (_GEN_1866 ? io_wb_resps_0_bits_predicated : ~_GEN_1833 & rob_predicated_3_11));
    rob_predicated_3_12 <= ~(_GEN_2151 & _GEN_666 | _GEN_2131 | _GEN_2085 & _GEN_538) & (_GEN_2065 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_410 | _GEN_1999 | _GEN_1953 & _GEN_282 | _GEN_1933 | _GEN_1887 & _GEN_154) & (_GEN_1867 ? io_wb_resps_0_bits_predicated : ~_GEN_1834 & rob_predicated_3_12));
    rob_predicated_3_13 <= ~(_GEN_2151 & _GEN_668 | _GEN_2132 | _GEN_2085 & _GEN_540) & (_GEN_2066 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_412 | _GEN_2000 | _GEN_1953 & _GEN_284 | _GEN_1934 | _GEN_1887 & _GEN_156) & (_GEN_1868 ? io_wb_resps_0_bits_predicated : ~_GEN_1835 & rob_predicated_3_13));
    rob_predicated_3_14 <= ~(_GEN_2151 & _GEN_670 | _GEN_2133 | _GEN_2085 & _GEN_542) & (_GEN_2067 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_414 | _GEN_2001 | _GEN_1953 & _GEN_286 | _GEN_1935 | _GEN_1887 & _GEN_158) & (_GEN_1869 ? io_wb_resps_0_bits_predicated : ~_GEN_1836 & rob_predicated_3_14));
    rob_predicated_3_15 <= ~(_GEN_2151 & _GEN_672 | _GEN_2134 | _GEN_2085 & _GEN_544) & (_GEN_2068 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_416 | _GEN_2002 | _GEN_1953 & _GEN_288 | _GEN_1936 | _GEN_1887 & _GEN_160) & (_GEN_1870 ? io_wb_resps_0_bits_predicated : ~_GEN_1837 & rob_predicated_3_15));
    rob_predicated_3_16 <= ~(_GEN_2151 & _GEN_674 | _GEN_2135 | _GEN_2085 & _GEN_546) & (_GEN_2069 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_418 | _GEN_2003 | _GEN_1953 & _GEN_290 | _GEN_1937 | _GEN_1887 & _GEN_162) & (_GEN_1871 ? io_wb_resps_0_bits_predicated : ~_GEN_1838 & rob_predicated_3_16));
    rob_predicated_3_17 <= ~(_GEN_2151 & _GEN_676 | _GEN_2136 | _GEN_2085 & _GEN_548) & (_GEN_2070 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_420 | _GEN_2004 | _GEN_1953 & _GEN_292 | _GEN_1938 | _GEN_1887 & _GEN_164) & (_GEN_1872 ? io_wb_resps_0_bits_predicated : ~_GEN_1839 & rob_predicated_3_17));
    rob_predicated_3_18 <= ~(_GEN_2151 & _GEN_678 | _GEN_2137 | _GEN_2085 & _GEN_550) & (_GEN_2071 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_422 | _GEN_2005 | _GEN_1953 & _GEN_294 | _GEN_1939 | _GEN_1887 & _GEN_166) & (_GEN_1873 ? io_wb_resps_0_bits_predicated : ~_GEN_1840 & rob_predicated_3_18));
    rob_predicated_3_19 <= ~(_GEN_2151 & _GEN_680 | _GEN_2138 | _GEN_2085 & _GEN_552) & (_GEN_2072 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_424 | _GEN_2006 | _GEN_1953 & _GEN_296 | _GEN_1940 | _GEN_1887 & _GEN_168) & (_GEN_1874 ? io_wb_resps_0_bits_predicated : ~_GEN_1841 & rob_predicated_3_19));
    rob_predicated_3_20 <= ~(_GEN_2151 & _GEN_682 | _GEN_2139 | _GEN_2085 & _GEN_554) & (_GEN_2073 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_426 | _GEN_2007 | _GEN_1953 & _GEN_298 | _GEN_1941 | _GEN_1887 & _GEN_170) & (_GEN_1875 ? io_wb_resps_0_bits_predicated : ~_GEN_1842 & rob_predicated_3_20));
    rob_predicated_3_21 <= ~(_GEN_2151 & _GEN_684 | _GEN_2140 | _GEN_2085 & _GEN_556) & (_GEN_2074 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_428 | _GEN_2008 | _GEN_1953 & _GEN_300 | _GEN_1942 | _GEN_1887 & _GEN_172) & (_GEN_1876 ? io_wb_resps_0_bits_predicated : ~_GEN_1843 & rob_predicated_3_21));
    rob_predicated_3_22 <= ~(_GEN_2151 & _GEN_686 | _GEN_2141 | _GEN_2085 & _GEN_558) & (_GEN_2075 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_430 | _GEN_2009 | _GEN_1953 & _GEN_302 | _GEN_1943 | _GEN_1887 & _GEN_174) & (_GEN_1877 ? io_wb_resps_0_bits_predicated : ~_GEN_1844 & rob_predicated_3_22));
    rob_predicated_3_23 <= ~(_GEN_2151 & _GEN_688 | _GEN_2142 | _GEN_2085 & _GEN_560) & (_GEN_2076 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_432 | _GEN_2010 | _GEN_1953 & _GEN_304 | _GEN_1944 | _GEN_1887 & _GEN_176) & (_GEN_1878 ? io_wb_resps_0_bits_predicated : ~_GEN_1845 & rob_predicated_3_23));
    rob_predicated_3_24 <= ~(_GEN_2151 & _GEN_690 | _GEN_2143 | _GEN_2085 & _GEN_562) & (_GEN_2077 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_434 | _GEN_2011 | _GEN_1953 & _GEN_306 | _GEN_1945 | _GEN_1887 & _GEN_178) & (_GEN_1879 ? io_wb_resps_0_bits_predicated : ~_GEN_1846 & rob_predicated_3_24));
    rob_predicated_3_25 <= ~(_GEN_2151 & _GEN_692 | _GEN_2144 | _GEN_2085 & _GEN_564) & (_GEN_2078 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_436 | _GEN_2012 | _GEN_1953 & _GEN_308 | _GEN_1946 | _GEN_1887 & _GEN_180) & (_GEN_1880 ? io_wb_resps_0_bits_predicated : ~_GEN_1847 & rob_predicated_3_25));
    rob_predicated_3_26 <= ~(_GEN_2151 & _GEN_694 | _GEN_2145 | _GEN_2085 & _GEN_566) & (_GEN_2079 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_438 | _GEN_2013 | _GEN_1953 & _GEN_310 | _GEN_1947 | _GEN_1887 & _GEN_182) & (_GEN_1881 ? io_wb_resps_0_bits_predicated : ~_GEN_1848 & rob_predicated_3_26));
    rob_predicated_3_27 <= ~(_GEN_2151 & _GEN_696 | _GEN_2146 | _GEN_2085 & _GEN_568) & (_GEN_2080 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_440 | _GEN_2014 | _GEN_1953 & _GEN_312 | _GEN_1948 | _GEN_1887 & _GEN_184) & (_GEN_1882 ? io_wb_resps_0_bits_predicated : ~_GEN_1849 & rob_predicated_3_27));
    rob_predicated_3_28 <= ~(_GEN_2151 & _GEN_698 | _GEN_2147 | _GEN_2085 & _GEN_570) & (_GEN_2081 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_442 | _GEN_2015 | _GEN_1953 & _GEN_314 | _GEN_1949 | _GEN_1887 & _GEN_186) & (_GEN_1883 ? io_wb_resps_0_bits_predicated : ~_GEN_1850 & rob_predicated_3_28));
    rob_predicated_3_29 <= ~(_GEN_2151 & _GEN_700 | _GEN_2148 | _GEN_2085 & _GEN_572) & (_GEN_2082 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_444 | _GEN_2016 | _GEN_1953 & _GEN_316 | _GEN_1950 | _GEN_1887 & _GEN_188) & (_GEN_1884 ? io_wb_resps_0_bits_predicated : ~_GEN_1851 & rob_predicated_3_29));
    rob_predicated_3_30 <= ~(_GEN_2151 & _GEN_702 | _GEN_2149 | _GEN_2085 & _GEN_574) & (_GEN_2083 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & _GEN_446 | _GEN_2017 | _GEN_1953 & _GEN_318 | _GEN_1951 | _GEN_1887 & _GEN_190) & (_GEN_1885 ? io_wb_resps_0_bits_predicated : ~_GEN_1852 & rob_predicated_3_30));
    rob_predicated_3_31 <= ~(_GEN_2151 & (&(io_wb_resps_9_bits_uop_rob_idx[6:2])) | _GEN_2150 | _GEN_2085 & (&(io_wb_resps_7_bits_uop_rob_idx[6:2]))) & (_GEN_2084 ? io_wb_resps_6_bits_predicated : ~(_GEN_2019 & (&(io_wb_resps_5_bits_uop_rob_idx[6:2])) | _GEN_2018 | _GEN_1953 & (&(io_wb_resps_3_bits_uop_rob_idx[6:2])) | _GEN_1952 | _GEN_1887 & (&(io_wb_resps_1_bits_uop_rob_idx[6:2]))) & (_GEN_1886 ? io_wb_resps_0_bits_predicated : ~_GEN_1853 & rob_predicated_3_31));
    block_commit_REG_1 <= exception_thrown;
    REG <= exception_thrown;
    REG_1 <= REG;
    REG_2 <= exception_thrown;
    io_com_load_is_at_rob_head_REG <= casez_tmp_96 & ~(_io_commit_valids_0_output | _io_commit_valids_1_output | _io_commit_valids_2_output | _io_commit_valids_3_output);
  end // always @(posedge)
  assign io_rob_tail_idx = rob_tail_idx;
  assign io_rob_head_idx = rob_head_idx;
  assign io_commit_valids_0 = _io_commit_valids_0_output;
  assign io_commit_valids_1 = _io_commit_valids_1_output;
  assign io_commit_valids_2 = _io_commit_valids_2_output;
  assign io_commit_valids_3 = _io_commit_valids_3_output;
  assign io_commit_arch_valids_0 = _io_commit_valids_0_output & ~casez_tmp_11;
  assign io_commit_arch_valids_1 = _io_commit_valids_1_output & ~casez_tmp_31;
  assign io_commit_arch_valids_2 = _io_commit_valids_2_output & ~casez_tmp_51;
  assign io_commit_arch_valids_3 = _io_commit_valids_3_output & ~casez_tmp_71;
  assign io_commit_uops_0_ftq_idx = casez_tmp_14;
  assign io_commit_uops_0_pdst = casez_tmp_17;
  assign io_commit_uops_0_stale_pdst = casez_tmp_18;
  assign io_commit_uops_0_is_fencei = casez_tmp_19;
  assign io_commit_uops_0_uses_ldq = casez_tmp_20;
  assign io_commit_uops_0_uses_stq = casez_tmp_21;
  assign io_commit_uops_0_ldst = casez_tmp_24;
  assign io_commit_uops_0_ldst_val = casez_tmp_25;
  assign io_commit_uops_0_dst_rtype = casez_tmp_26;
  assign io_commit_uops_1_ftq_idx = casez_tmp_34;
  assign io_commit_uops_1_pdst = casez_tmp_37;
  assign io_commit_uops_1_stale_pdst = casez_tmp_38;
  assign io_commit_uops_1_is_fencei = casez_tmp_39;
  assign io_commit_uops_1_uses_ldq = casez_tmp_40;
  assign io_commit_uops_1_uses_stq = casez_tmp_41;
  assign io_commit_uops_1_ldst = casez_tmp_44;
  assign io_commit_uops_1_ldst_val = casez_tmp_45;
  assign io_commit_uops_1_dst_rtype = casez_tmp_46;
  assign io_commit_uops_2_ftq_idx = casez_tmp_54;
  assign io_commit_uops_2_pdst = casez_tmp_57;
  assign io_commit_uops_2_stale_pdst = casez_tmp_58;
  assign io_commit_uops_2_is_fencei = casez_tmp_59;
  assign io_commit_uops_2_uses_ldq = casez_tmp_60;
  assign io_commit_uops_2_uses_stq = casez_tmp_61;
  assign io_commit_uops_2_ldst = casez_tmp_64;
  assign io_commit_uops_2_ldst_val = casez_tmp_65;
  assign io_commit_uops_2_dst_rtype = casez_tmp_66;
  assign io_commit_uops_3_ftq_idx = casez_tmp_74;
  assign io_commit_uops_3_pdst = casez_tmp_77;
  assign io_commit_uops_3_stale_pdst = casez_tmp_78;
  assign io_commit_uops_3_is_fencei = casez_tmp_79;
  assign io_commit_uops_3_uses_ldq = casez_tmp_80;
  assign io_commit_uops_3_uses_stq = casez_tmp_81;
  assign io_commit_uops_3_ldst = casez_tmp_84;
  assign io_commit_uops_3_ldst_val = casez_tmp_85;
  assign io_commit_uops_3_dst_rtype = casez_tmp_86;
  assign io_commit_fflags_valid = fflags_val_0 | fflags_val_1 | fflags_val_2 | fflags_val_3;
  assign io_commit_fflags_bits = (fflags_val_0 ? casez_tmp_29 : 5'h0) | (fflags_val_1 ? casez_tmp_49 : 5'h0) | (fflags_val_2 ? casez_tmp_69 : 5'h0) | (fflags_val_3 ? casez_tmp_89 : 5'h0);
  assign io_commit_rbk_valids_0 = _io_commit_rbk_valids_0_output;
  assign io_commit_rbk_valids_1 = _io_commit_rbk_valids_1_output;
  assign io_commit_rbk_valids_2 = _io_commit_rbk_valids_2_output;
  assign io_commit_rbk_valids_3 = _io_commit_rbk_valids_3_output;
  assign io_commit_rollback = _io_commit_rollback_T_3;
  assign io_com_load_is_at_rob_head = io_com_load_is_at_rob_head_REG;
  assign io_com_xcpt_valid = exception_thrown & ~is_mini_exception;
  assign io_com_xcpt_bits_ftq_idx = com_xcpt_uop_ftq_idx;
  assign io_com_xcpt_bits_edge_inst = com_xcpt_uop_edge_inst;
  assign io_com_xcpt_bits_pc_lob = com_xcpt_uop_pc_lob;
  assign io_com_xcpt_bits_cause = r_xcpt_uop_exc_cause;
  assign io_com_xcpt_bits_badvaddr = {{24{r_xcpt_badvaddr[39]}}, r_xcpt_badvaddr};
  assign io_flush_valid = _io_flush_valid_output;
  assign io_flush_bits_ftq_idx = exception_thrown ? com_xcpt_uop_ftq_idx : (flush_commit_mask_0 ? casez_tmp_14 : 6'h0) | (flush_commit_mask_1 ? casez_tmp_34 : 6'h0) | (flush_commit_mask_2 ? casez_tmp_54 : 6'h0) | (flush_commit_mask_3 ? casez_tmp_74 : 6'h0);
  assign io_flush_bits_edge_inst = exception_thrown ? com_xcpt_uop_edge_inst : flush_commit_mask_0 & casez_tmp_15 | flush_commit_mask_1 & casez_tmp_35 | flush_commit_mask_2 & casez_tmp_55 | flush_commit_mask_3 & casez_tmp_75;
  assign io_flush_bits_is_rvc = exception_thrown ? (casez_tmp ? casez_tmp_13 : casez_tmp_2 ? casez_tmp_33 : casez_tmp_5 ? casez_tmp_53 : casez_tmp_73) : flush_commit_mask_0 & casez_tmp_13 | flush_commit_mask_1 & casez_tmp_33 | flush_commit_mask_2 & casez_tmp_53 | flush_commit_mask_3 & casez_tmp_73;
  assign io_flush_bits_pc_lob = exception_thrown ? com_xcpt_uop_pc_lob : (flush_commit_mask_0 ? casez_tmp_16 : 6'h0) | (flush_commit_mask_1 ? casez_tmp_36 : 6'h0) | (flush_commit_mask_2 ? casez_tmp_56 : 6'h0) | (flush_commit_mask_3 ? casez_tmp_76 : 6'h0);
  assign io_flush_bits_flush_typ = _io_flush_valid_output ? (flush_commit & (exception_thrown ? (casez_tmp ? casez_tmp_12 : casez_tmp_2 ? casez_tmp_32 : casez_tmp_5 ? casez_tmp_52 : casez_tmp_72) : (flush_commit_mask_0 ? casez_tmp_12 : 7'h0) | (flush_commit_mask_1 ? casez_tmp_32 : 7'h0) | (flush_commit_mask_2 ? casez_tmp_52 : 7'h0) | (flush_commit_mask_3 ? casez_tmp_72 : 7'h0)) == 7'h6A ? 3'h3 : exception_thrown & ~is_mini_exception ? 3'h1 : exception_thrown | (casez_tmp | casez_tmp_2 | casez_tmp_5 | casez_tmp_8) & (casez_tmp ? casez_tmp_22 : casez_tmp_2 ? casez_tmp_42 : casez_tmp_5 ? casez_tmp_62 : casez_tmp_82) ? 3'h2 : 3'h4) : 3'h0;
  assign io_empty = empty;
  assign io_ready = _io_ready_T & ~full & ~r_xcpt_val;
  assign io_flush_frontend = r_xcpt_val;
endmodule

