// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

module LSU(
  input         clock,
                reset,
                io_ptw_req_ready,
                io_ptw_resp_valid,
                io_ptw_resp_bits_ae_final,
  input  [43:0] io_ptw_resp_bits_pte_ppn,
  input         io_ptw_resp_bits_pte_d,
                io_ptw_resp_bits_pte_a,
                io_ptw_resp_bits_pte_g,
                io_ptw_resp_bits_pte_u,
                io_ptw_resp_bits_pte_x,
                io_ptw_resp_bits_pte_w,
                io_ptw_resp_bits_pte_r,
                io_ptw_resp_bits_pte_v,
  input  [1:0]  io_ptw_resp_bits_level,
  input         io_ptw_resp_bits_homogeneous,
  input  [3:0]  io_ptw_ptbr_mode,
  input  [1:0]  io_ptw_status_dprv,
  input         io_ptw_status_mxr,
                io_ptw_status_sum,
                io_ptw_pmp_0_cfg_l,
  input  [1:0]  io_ptw_pmp_0_cfg_a,
  input         io_ptw_pmp_0_cfg_x,
                io_ptw_pmp_0_cfg_w,
                io_ptw_pmp_0_cfg_r,
  input  [29:0] io_ptw_pmp_0_addr,
  input  [31:0] io_ptw_pmp_0_mask,
  input         io_ptw_pmp_1_cfg_l,
  input  [1:0]  io_ptw_pmp_1_cfg_a,
  input         io_ptw_pmp_1_cfg_x,
                io_ptw_pmp_1_cfg_w,
                io_ptw_pmp_1_cfg_r,
  input  [29:0] io_ptw_pmp_1_addr,
  input  [31:0] io_ptw_pmp_1_mask,
  input         io_ptw_pmp_2_cfg_l,
  input  [1:0]  io_ptw_pmp_2_cfg_a,
  input         io_ptw_pmp_2_cfg_x,
                io_ptw_pmp_2_cfg_w,
                io_ptw_pmp_2_cfg_r,
  input  [29:0] io_ptw_pmp_2_addr,
  input  [31:0] io_ptw_pmp_2_mask,
  input         io_ptw_pmp_3_cfg_l,
  input  [1:0]  io_ptw_pmp_3_cfg_a,
  input         io_ptw_pmp_3_cfg_x,
                io_ptw_pmp_3_cfg_w,
                io_ptw_pmp_3_cfg_r,
  input  [29:0] io_ptw_pmp_3_addr,
  input  [31:0] io_ptw_pmp_3_mask,
  input         io_ptw_pmp_4_cfg_l,
  input  [1:0]  io_ptw_pmp_4_cfg_a,
  input         io_ptw_pmp_4_cfg_x,
                io_ptw_pmp_4_cfg_w,
                io_ptw_pmp_4_cfg_r,
  input  [29:0] io_ptw_pmp_4_addr,
  input  [31:0] io_ptw_pmp_4_mask,
  input         io_ptw_pmp_5_cfg_l,
  input  [1:0]  io_ptw_pmp_5_cfg_a,
  input         io_ptw_pmp_5_cfg_x,
                io_ptw_pmp_5_cfg_w,
                io_ptw_pmp_5_cfg_r,
  input  [29:0] io_ptw_pmp_5_addr,
  input  [31:0] io_ptw_pmp_5_mask,
  input         io_ptw_pmp_6_cfg_l,
  input  [1:0]  io_ptw_pmp_6_cfg_a,
  input         io_ptw_pmp_6_cfg_x,
                io_ptw_pmp_6_cfg_w,
                io_ptw_pmp_6_cfg_r,
  input  [29:0] io_ptw_pmp_6_addr,
  input  [31:0] io_ptw_pmp_6_mask,
  input         io_ptw_pmp_7_cfg_l,
  input  [1:0]  io_ptw_pmp_7_cfg_a,
  input         io_ptw_pmp_7_cfg_x,
                io_ptw_pmp_7_cfg_w,
                io_ptw_pmp_7_cfg_r,
  input  [29:0] io_ptw_pmp_7_addr,
  input  [31:0] io_ptw_pmp_7_mask,
  input         io_core_exe_0_req_valid,
                io_core_exe_0_req_bits_uop_ctrl_is_load,
                io_core_exe_0_req_bits_uop_ctrl_is_sta,
                io_core_exe_0_req_bits_uop_ctrl_is_std,
  input  [19:0] io_core_exe_0_req_bits_uop_br_mask,
  input  [6:0]  io_core_exe_0_req_bits_uop_rob_idx,
  input  [4:0]  io_core_exe_0_req_bits_uop_ldq_idx,
                io_core_exe_0_req_bits_uop_stq_idx,
  input  [6:0]  io_core_exe_0_req_bits_uop_pdst,
  input  [4:0]  io_core_exe_0_req_bits_uop_mem_cmd,
  input  [1:0]  io_core_exe_0_req_bits_uop_mem_size,
  input         io_core_exe_0_req_bits_uop_mem_signed,
                io_core_exe_0_req_bits_uop_is_fence,
                io_core_exe_0_req_bits_uop_is_amo,
                io_core_exe_0_req_bits_uop_uses_ldq,
                io_core_exe_0_req_bits_uop_uses_stq,
                io_core_exe_0_req_bits_uop_fp_val,
  input  [63:0] io_core_exe_0_req_bits_data,
  input  [39:0] io_core_exe_0_req_bits_addr,
  input         io_core_exe_0_req_bits_mxcpt_valid,
                io_core_exe_0_req_bits_sfence_valid,
                io_core_exe_0_req_bits_sfence_bits_rs1,
                io_core_exe_0_req_bits_sfence_bits_rs2,
  input  [38:0] io_core_exe_0_req_bits_sfence_bits_addr,
  input         io_core_exe_1_req_valid,
                io_core_exe_1_req_bits_uop_ctrl_is_load,
                io_core_exe_1_req_bits_uop_ctrl_is_sta,
                io_core_exe_1_req_bits_uop_ctrl_is_std,
  input  [19:0] io_core_exe_1_req_bits_uop_br_mask,
  input  [6:0]  io_core_exe_1_req_bits_uop_rob_idx,
  input  [4:0]  io_core_exe_1_req_bits_uop_ldq_idx,
                io_core_exe_1_req_bits_uop_stq_idx,
  input  [6:0]  io_core_exe_1_req_bits_uop_pdst,
  input  [4:0]  io_core_exe_1_req_bits_uop_mem_cmd,
  input  [1:0]  io_core_exe_1_req_bits_uop_mem_size,
  input         io_core_exe_1_req_bits_uop_mem_signed,
                io_core_exe_1_req_bits_uop_is_fence,
                io_core_exe_1_req_bits_uop_is_amo,
                io_core_exe_1_req_bits_uop_uses_ldq,
                io_core_exe_1_req_bits_uop_uses_stq,
                io_core_exe_1_req_bits_uop_fp_val,
  input  [63:0] io_core_exe_1_req_bits_data,
  input  [39:0] io_core_exe_1_req_bits_addr,
  input         io_core_exe_1_req_bits_mxcpt_valid,
                io_core_exe_1_req_bits_sfence_valid,
                io_core_exe_1_req_bits_sfence_bits_rs1,
                io_core_exe_1_req_bits_sfence_bits_rs2,
  input  [38:0] io_core_exe_1_req_bits_sfence_bits_addr,
  input         io_core_dis_uops_0_valid,
  input  [6:0]  io_core_dis_uops_0_bits_uopc,
  input         io_core_dis_uops_0_bits_ctrl_is_load,
                io_core_dis_uops_0_bits_ctrl_is_sta,
  input  [19:0] io_core_dis_uops_0_bits_br_mask,
  input  [6:0]  io_core_dis_uops_0_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_0_bits_ldq_idx,
                io_core_dis_uops_0_bits_stq_idx,
  input  [6:0]  io_core_dis_uops_0_bits_pdst,
  input         io_core_dis_uops_0_bits_exception,
  input  [4:0]  io_core_dis_uops_0_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_0_bits_mem_size,
  input         io_core_dis_uops_0_bits_mem_signed,
                io_core_dis_uops_0_bits_is_fence,
                io_core_dis_uops_0_bits_is_amo,
                io_core_dis_uops_0_bits_uses_ldq,
                io_core_dis_uops_0_bits_uses_stq,
  input  [1:0]  io_core_dis_uops_0_bits_dst_rtype,
  input         io_core_dis_uops_0_bits_fp_val,
                io_core_dis_uops_1_valid,
  input  [6:0]  io_core_dis_uops_1_bits_uopc,
  input         io_core_dis_uops_1_bits_ctrl_is_load,
                io_core_dis_uops_1_bits_ctrl_is_sta,
  input  [19:0] io_core_dis_uops_1_bits_br_mask,
  input  [6:0]  io_core_dis_uops_1_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_1_bits_ldq_idx,
                io_core_dis_uops_1_bits_stq_idx,
  input  [6:0]  io_core_dis_uops_1_bits_pdst,
  input         io_core_dis_uops_1_bits_exception,
  input  [4:0]  io_core_dis_uops_1_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_1_bits_mem_size,
  input         io_core_dis_uops_1_bits_mem_signed,
                io_core_dis_uops_1_bits_is_fence,
                io_core_dis_uops_1_bits_is_amo,
                io_core_dis_uops_1_bits_uses_ldq,
                io_core_dis_uops_1_bits_uses_stq,
  input  [1:0]  io_core_dis_uops_1_bits_dst_rtype,
  input         io_core_dis_uops_1_bits_fp_val,
                io_core_dis_uops_2_valid,
  input  [6:0]  io_core_dis_uops_2_bits_uopc,
  input         io_core_dis_uops_2_bits_ctrl_is_load,
                io_core_dis_uops_2_bits_ctrl_is_sta,
  input  [19:0] io_core_dis_uops_2_bits_br_mask,
  input  [6:0]  io_core_dis_uops_2_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_2_bits_ldq_idx,
                io_core_dis_uops_2_bits_stq_idx,
  input  [6:0]  io_core_dis_uops_2_bits_pdst,
  input         io_core_dis_uops_2_bits_exception,
  input  [4:0]  io_core_dis_uops_2_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_2_bits_mem_size,
  input         io_core_dis_uops_2_bits_mem_signed,
                io_core_dis_uops_2_bits_is_fence,
                io_core_dis_uops_2_bits_is_amo,
                io_core_dis_uops_2_bits_uses_ldq,
                io_core_dis_uops_2_bits_uses_stq,
  input  [1:0]  io_core_dis_uops_2_bits_dst_rtype,
  input         io_core_dis_uops_2_bits_fp_val,
                io_core_dis_uops_3_valid,
  input  [6:0]  io_core_dis_uops_3_bits_uopc,
  input         io_core_dis_uops_3_bits_ctrl_is_load,
                io_core_dis_uops_3_bits_ctrl_is_sta,
  input  [19:0] io_core_dis_uops_3_bits_br_mask,
  input  [6:0]  io_core_dis_uops_3_bits_rob_idx,
  input  [4:0]  io_core_dis_uops_3_bits_ldq_idx,
                io_core_dis_uops_3_bits_stq_idx,
  input  [6:0]  io_core_dis_uops_3_bits_pdst,
  input         io_core_dis_uops_3_bits_exception,
  input  [4:0]  io_core_dis_uops_3_bits_mem_cmd,
  input  [1:0]  io_core_dis_uops_3_bits_mem_size,
  input         io_core_dis_uops_3_bits_mem_signed,
                io_core_dis_uops_3_bits_is_fence,
                io_core_dis_uops_3_bits_is_amo,
                io_core_dis_uops_3_bits_uses_ldq,
                io_core_dis_uops_3_bits_uses_stq,
  input  [1:0]  io_core_dis_uops_3_bits_dst_rtype,
  input         io_core_dis_uops_3_bits_fp_val,
                io_core_fp_stdata_valid,
  input  [19:0] io_core_fp_stdata_bits_uop_br_mask,
  input  [6:0]  io_core_fp_stdata_bits_uop_rob_idx,
  input  [4:0]  io_core_fp_stdata_bits_uop_stq_idx,
  input  [63:0] io_core_fp_stdata_bits_data,
  input         io_core_commit_valids_0,
                io_core_commit_valids_1,
                io_core_commit_valids_2,
                io_core_commit_valids_3,
                io_core_commit_uops_0_uses_ldq,
                io_core_commit_uops_0_uses_stq,
                io_core_commit_uops_1_uses_ldq,
                io_core_commit_uops_1_uses_stq,
                io_core_commit_uops_2_uses_ldq,
                io_core_commit_uops_2_uses_stq,
                io_core_commit_uops_3_uses_ldq,
                io_core_commit_uops_3_uses_stq,
                io_core_commit_load_at_rob_head,
                io_core_fence_dmem,
  input  [19:0] io_core_brupdate_b1_resolve_mask,
                io_core_brupdate_b1_mispredict_mask,
  input  [4:0]  io_core_brupdate_b2_uop_ldq_idx,
                io_core_brupdate_b2_uop_stq_idx,
  input         io_core_brupdate_b2_mispredict,
  input  [6:0]  io_core_rob_head_idx,
  input         io_core_exception,
                io_dmem_req_ready,
                io_dmem_resp_0_valid,
  input  [4:0]  io_dmem_resp_0_bits_uop_ldq_idx,
                io_dmem_resp_0_bits_uop_stq_idx,
  input         io_dmem_resp_0_bits_uop_is_amo,
                io_dmem_resp_0_bits_uop_uses_ldq,
                io_dmem_resp_0_bits_uop_uses_stq,
  input  [63:0] io_dmem_resp_0_bits_data,
  input         io_dmem_resp_0_bits_is_hella,
                io_dmem_resp_1_valid,
  input  [4:0]  io_dmem_resp_1_bits_uop_ldq_idx,
                io_dmem_resp_1_bits_uop_stq_idx,
  input         io_dmem_resp_1_bits_uop_is_amo,
                io_dmem_resp_1_bits_uop_uses_ldq,
                io_dmem_resp_1_bits_uop_uses_stq,
  input  [63:0] io_dmem_resp_1_bits_data,
  input         io_dmem_resp_1_bits_is_hella,
                io_dmem_nack_0_valid,
  input  [4:0]  io_dmem_nack_0_bits_uop_ldq_idx,
                io_dmem_nack_0_bits_uop_stq_idx,
  input         io_dmem_nack_0_bits_uop_uses_ldq,
                io_dmem_nack_0_bits_uop_uses_stq,
                io_dmem_nack_0_bits_is_hella,
                io_dmem_nack_1_valid,
  input  [4:0]  io_dmem_nack_1_bits_uop_ldq_idx,
                io_dmem_nack_1_bits_uop_stq_idx,
  input         io_dmem_nack_1_bits_uop_uses_ldq,
                io_dmem_nack_1_bits_uop_uses_stq,
                io_dmem_nack_1_bits_is_hella,
                io_dmem_release_valid,
  input  [31:0] io_dmem_release_bits_address,
  input         io_dmem_ordered,
                io_hellacache_req_valid,
  input  [39:0] io_hellacache_req_bits_addr,
  input         io_hellacache_s1_kill,
  output        io_ptw_req_valid,
                io_ptw_req_bits_valid,
  output [26:0] io_ptw_req_bits_bits_addr,
  output        io_core_exe_0_iresp_valid,
  output [6:0]  io_core_exe_0_iresp_bits_uop_rob_idx,
                io_core_exe_0_iresp_bits_uop_pdst,
  output        io_core_exe_0_iresp_bits_uop_is_amo,
                io_core_exe_0_iresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_iresp_bits_uop_dst_rtype,
  output [63:0] io_core_exe_0_iresp_bits_data,
  output        io_core_exe_0_fresp_valid,
  output [6:0]  io_core_exe_0_fresp_bits_uop_uopc,
  output [19:0] io_core_exe_0_fresp_bits_uop_br_mask,
  output [6:0]  io_core_exe_0_fresp_bits_uop_rob_idx,
  output [4:0]  io_core_exe_0_fresp_bits_uop_stq_idx,
  output [6:0]  io_core_exe_0_fresp_bits_uop_pdst,
  output [1:0]  io_core_exe_0_fresp_bits_uop_mem_size,
  output        io_core_exe_0_fresp_bits_uop_is_amo,
                io_core_exe_0_fresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_0_fresp_bits_uop_dst_rtype,
  output        io_core_exe_0_fresp_bits_uop_fp_val,
  output [64:0] io_core_exe_0_fresp_bits_data,
  output        io_core_exe_1_iresp_valid,
  output [6:0]  io_core_exe_1_iresp_bits_uop_rob_idx,
                io_core_exe_1_iresp_bits_uop_pdst,
  output        io_core_exe_1_iresp_bits_uop_is_amo,
                io_core_exe_1_iresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_1_iresp_bits_uop_dst_rtype,
  output [63:0] io_core_exe_1_iresp_bits_data,
  output        io_core_exe_1_fresp_valid,
  output [6:0]  io_core_exe_1_fresp_bits_uop_uopc,
  output [19:0] io_core_exe_1_fresp_bits_uop_br_mask,
  output [6:0]  io_core_exe_1_fresp_bits_uop_rob_idx,
  output [4:0]  io_core_exe_1_fresp_bits_uop_stq_idx,
  output [6:0]  io_core_exe_1_fresp_bits_uop_pdst,
  output [1:0]  io_core_exe_1_fresp_bits_uop_mem_size,
  output        io_core_exe_1_fresp_bits_uop_is_amo,
                io_core_exe_1_fresp_bits_uop_uses_stq,
  output [1:0]  io_core_exe_1_fresp_bits_uop_dst_rtype,
  output        io_core_exe_1_fresp_bits_uop_fp_val,
  output [64:0] io_core_exe_1_fresp_bits_data,
  output [4:0]  io_core_dis_ldq_idx_0,
                io_core_dis_ldq_idx_1,
                io_core_dis_ldq_idx_2,
                io_core_dis_ldq_idx_3,
                io_core_dis_stq_idx_0,
                io_core_dis_stq_idx_1,
                io_core_dis_stq_idx_2,
                io_core_dis_stq_idx_3,
  output        io_core_ldq_full_0,
                io_core_ldq_full_1,
                io_core_ldq_full_2,
                io_core_ldq_full_3,
                io_core_stq_full_0,
                io_core_stq_full_1,
                io_core_stq_full_2,
                io_core_stq_full_3,
                io_core_fp_stdata_ready,
                io_core_clr_bsy_0_valid,
  output [6:0]  io_core_clr_bsy_0_bits,
  output        io_core_clr_bsy_1_valid,
  output [6:0]  io_core_clr_bsy_1_bits,
  output        io_core_clr_bsy_2_valid,
  output [6:0]  io_core_clr_bsy_2_bits,
  output        io_core_spec_ld_wakeup_0_valid,
  output [6:0]  io_core_spec_ld_wakeup_0_bits,
  output        io_core_spec_ld_wakeup_1_valid,
  output [6:0]  io_core_spec_ld_wakeup_1_bits,
  output        io_core_ld_miss,
                io_core_fencei_rdy,
                io_core_lxcpt_valid,
  output [19:0] io_core_lxcpt_bits_uop_br_mask,
  output [6:0]  io_core_lxcpt_bits_uop_rob_idx,
  output [4:0]  io_core_lxcpt_bits_cause,
  output [39:0] io_core_lxcpt_bits_badvaddr,
  output        io_dmem_req_valid,
                io_dmem_req_bits_0_valid,
  output [19:0] io_dmem_req_bits_0_bits_uop_br_mask,
  output [4:0]  io_dmem_req_bits_0_bits_uop_ldq_idx,
                io_dmem_req_bits_0_bits_uop_stq_idx,
                io_dmem_req_bits_0_bits_uop_mem_cmd,
  output [1:0]  io_dmem_req_bits_0_bits_uop_mem_size,
  output        io_dmem_req_bits_0_bits_uop_mem_signed,
                io_dmem_req_bits_0_bits_uop_is_amo,
                io_dmem_req_bits_0_bits_uop_uses_ldq,
                io_dmem_req_bits_0_bits_uop_uses_stq,
  output [39:0] io_dmem_req_bits_0_bits_addr,
  output [63:0] io_dmem_req_bits_0_bits_data,
  output        io_dmem_req_bits_1_valid,
  output [19:0] io_dmem_req_bits_1_bits_uop_br_mask,
  output [4:0]  io_dmem_req_bits_1_bits_uop_ldq_idx,
                io_dmem_req_bits_1_bits_uop_stq_idx,
                io_dmem_req_bits_1_bits_uop_mem_cmd,
  output [1:0]  io_dmem_req_bits_1_bits_uop_mem_size,
  output        io_dmem_req_bits_1_bits_uop_mem_signed,
                io_dmem_req_bits_1_bits_uop_is_amo,
                io_dmem_req_bits_1_bits_uop_uses_ldq,
                io_dmem_req_bits_1_bits_uop_uses_stq,
  output [39:0] io_dmem_req_bits_1_bits_addr,
  output [63:0] io_dmem_req_bits_1_bits_data,
  output        io_dmem_req_bits_1_bits_is_hella,
                io_dmem_s1_kill_0,
                io_dmem_s1_kill_1,
  output [19:0] io_dmem_brupdate_b1_resolve_mask,
                io_dmem_brupdate_b1_mispredict_mask,
  output        io_dmem_exception,
                io_dmem_release_ready,
                io_dmem_force_order,
                io_hellacache_req_ready,
                io_hellacache_s2_nack,
                io_hellacache_resp_valid,
  output [63:0] io_hellacache_resp_bits_data,
  output        io_hellacache_s2_xcpt_ae_ld
);

  wire        _will_fire_store_commit_0_T_2;
  wire        _will_fire_store_commit_1_T_2;
  wire [4:0]  _forwarding_age_logic_1_io_forwarding_idx;
  wire [4:0]  _forwarding_age_logic_0_io_forwarding_idx;
  wire        _dtlb_io_miss_rdy;
  wire        _dtlb_io_resp_0_miss;
  wire [31:0] _dtlb_io_resp_0_paddr;
  wire        _dtlb_io_resp_0_pf_ld;
  wire        _dtlb_io_resp_0_pf_st;
  wire        _dtlb_io_resp_0_ae_ld;
  wire        _dtlb_io_resp_0_ae_st;
  wire        _dtlb_io_resp_0_cacheable;
  wire        _dtlb_io_resp_1_miss;
  wire [31:0] _dtlb_io_resp_1_paddr;
  wire        _dtlb_io_resp_1_pf_ld;
  wire        _dtlb_io_resp_1_pf_st;
  wire        _dtlb_io_resp_1_ae_ld;
  wire        _dtlb_io_resp_1_ae_st;
  wire        _dtlb_io_resp_1_ma_ld;
  wire        _dtlb_io_resp_1_ma_st;
  wire        _dtlb_io_resp_1_cacheable;
  reg         casez_tmp;
  reg         casez_tmp_0;
  reg         casez_tmp_1;
  reg         casez_tmp_2;
  reg         casez_tmp_3;
  reg  [19:0] casez_tmp_4;
  reg  [4:0]  casez_tmp_5;
  reg  [1:0]  casez_tmp_6;
  reg  [31:0] casez_tmp_7;
  reg  [19:0] casez_tmp_8;
  reg  [4:0]  casez_tmp_9;
  reg  [1:0]  casez_tmp_10;
  reg  [31:0] casez_tmp_11;
  reg         casez_tmp_12;
  reg  [19:0] casez_tmp_13;
  reg  [6:0]  casez_tmp_14;
  reg  [4:0]  casez_tmp_15;
  reg  [1:0]  casez_tmp_16;
  reg         casez_tmp_17;
  reg         casez_tmp_18;
  reg         casez_tmp_19;
  reg         casez_tmp_20;
  reg         casez_tmp_21;
  reg  [19:0] casez_tmp_22;
  reg  [6:0]  casez_tmp_23;
  reg  [4:0]  casez_tmp_24;
  reg  [1:0]  casez_tmp_25;
  reg         casez_tmp_26;
  reg         casez_tmp_27;
  reg         casez_tmp_28;
  reg         casez_tmp_29;
  reg         casez_tmp_30;
  reg         casez_tmp_31;
  reg         casez_tmp_32;
  reg         casez_tmp_33;
  reg         casez_tmp_34;
  reg         casez_tmp_35;
  reg         casez_tmp_36;
  reg         casez_tmp_37;
  reg         casez_tmp_38;
  reg  [31:0] casez_tmp_39;
  reg         casez_tmp_40;
  reg         casez_tmp_41;
  reg         casez_tmp_42;
  reg         casez_tmp_43;
  reg         casez_tmp_44;
  reg         casez_tmp_45;
  reg         casez_tmp_46;
  reg         casez_tmp_47;
  reg         casez_tmp_48;
  reg         casez_tmp_49;
  reg         casez_tmp_50;
  reg         casez_tmp_51;
  reg         casez_tmp_52;
  reg         casez_tmp_53;
  reg         casez_tmp_54;
  reg         casez_tmp_55;
  reg  [19:0] casez_tmp_56;
  reg  [6:0]  casez_tmp_57;
  reg  [4:0]  casez_tmp_58;
  reg  [4:0]  casez_tmp_59;
  reg  [6:0]  casez_tmp_60;
  reg  [4:0]  casez_tmp_61;
  reg  [1:0]  casez_tmp_62;
  reg         casez_tmp_63;
  reg         casez_tmp_64;
  reg         casez_tmp_65;
  reg         casez_tmp_66;
  reg  [19:0] casez_tmp_67;
  reg  [6:0]  casez_tmp_68;
  reg  [4:0]  casez_tmp_69;
  reg  [4:0]  casez_tmp_70;
  reg  [6:0]  casez_tmp_71;
  reg  [4:0]  casez_tmp_72;
  reg  [1:0]  casez_tmp_73;
  reg         casez_tmp_74;
  reg         casez_tmp_75;
  reg         casez_tmp_76;
  reg         casez_tmp_77;
  reg  [39:0] casez_tmp_78;
  reg  [39:0] casez_tmp_79;
  reg  [39:0] casez_tmp_80;
  reg  [1:0]  casez_tmp_81;
  reg  [63:0] casez_tmp_82;
  reg  [63:0] casez_tmp_83;
  reg  [19:0] casez_tmp_84;
  reg  [4:0]  casez_tmp_85;
  reg  [4:0]  casez_tmp_86;
  reg  [4:0]  casez_tmp_87;
  reg         casez_tmp_88;
  reg         casez_tmp_89;
  reg         casez_tmp_90;
  reg  [39:0] casez_tmp_91;
  reg  [19:0] casez_tmp_92;
  reg  [4:0]  casez_tmp_93;
  reg  [4:0]  casez_tmp_94;
  reg  [4:0]  casez_tmp_95;
  reg  [1:0]  casez_tmp_96;
  reg         casez_tmp_97;
  reg         casez_tmp_98;
  reg         casez_tmp_99;
  reg         casez_tmp_100;
  reg  [63:0] casez_tmp_101;
  reg  [31:0] casez_tmp_102;
  reg         casez_tmp_103;
  reg         casez_tmp_104;
  reg         casez_tmp_105;
  reg         casez_tmp_106;
  reg         casez_tmp_107;
  reg  [7:0]  casez_tmp_108;
  reg  [7:0]  casez_tmp_109;
  reg         casez_tmp_110;
  reg         casez_tmp_111;
  reg  [7:0]  casez_tmp_112;
  reg  [7:0]  casez_tmp_113;
  reg  [7:0]  casez_tmp_114;
  reg  [7:0]  casez_tmp_115;
  reg  [7:0]  casez_tmp_116;
  reg  [7:0]  casez_tmp_117;
  reg  [7:0]  casez_tmp_118;
  reg  [7:0]  casez_tmp_119;
  reg  [7:0]  casez_tmp_120;
  reg  [7:0]  casez_tmp_121;
  reg  [7:0]  casez_tmp_122;
  reg  [7:0]  casez_tmp_123;
  reg  [7:0]  casez_tmp_124;
  reg  [7:0]  casez_tmp_125;
  reg  [7:0]  casez_tmp_126;
  reg  [7:0]  casez_tmp_127;
  reg  [7:0]  casez_tmp_128;
  reg  [7:0]  casez_tmp_129;
  reg  [7:0]  casez_tmp_130;
  reg  [7:0]  casez_tmp_131;
  reg  [7:0]  casez_tmp_132;
  reg  [7:0]  casez_tmp_133;
  reg  [7:0]  casez_tmp_134;
  reg  [7:0]  casez_tmp_135;
  reg  [7:0]  casez_tmp_136;
  reg  [7:0]  casez_tmp_137;
  reg  [7:0]  casez_tmp_138;
  reg  [7:0]  casez_tmp_139;
  reg  [7:0]  casez_tmp_140;
  reg  [7:0]  casez_tmp_141;
  reg  [7:0]  casez_tmp_142;
  reg  [7:0]  casez_tmp_143;
  reg  [7:0]  casez_tmp_144;
  reg  [7:0]  casez_tmp_145;
  reg  [7:0]  casez_tmp_146;
  reg  [7:0]  casez_tmp_147;
  reg  [7:0]  casez_tmp_148;
  reg  [7:0]  casez_tmp_149;
  reg  [7:0]  casez_tmp_150;
  reg  [7:0]  casez_tmp_151;
  reg  [7:0]  casez_tmp_152;
  reg  [7:0]  casez_tmp_153;
  reg  [7:0]  casez_tmp_154;
  reg  [7:0]  casez_tmp_155;
  reg  [7:0]  casez_tmp_156;
  reg  [7:0]  casez_tmp_157;
  reg  [7:0]  casez_tmp_158;
  reg  [7:0]  casez_tmp_159;
  reg  [7:0]  casez_tmp_160;
  reg  [7:0]  casez_tmp_161;
  reg  [7:0]  casez_tmp_162;
  reg  [7:0]  casez_tmp_163;
  reg  [7:0]  casez_tmp_164;
  reg  [7:0]  casez_tmp_165;
  reg  [7:0]  casez_tmp_166;
  reg  [7:0]  casez_tmp_167;
  reg  [7:0]  casez_tmp_168;
  reg  [7:0]  casez_tmp_169;
  reg  [7:0]  casez_tmp_170;
  reg  [7:0]  casez_tmp_171;
  reg  [7:0]  casez_tmp_172;
  reg  [7:0]  casez_tmp_173;
  reg  [7:0]  casez_tmp_174;
  reg  [7:0]  casez_tmp_175;
  reg         casez_tmp_176;
  reg         casez_tmp_177;
  reg  [6:0]  casez_tmp_178;
  reg  [19:0] casez_tmp_179;
  reg  [1:0]  casez_tmp_180;
  reg  [6:0]  casez_tmp_181;
  reg  [19:0] casez_tmp_182;
  reg  [6:0]  casez_tmp_183;
  reg  [4:0]  casez_tmp_184;
  reg  [4:0]  casez_tmp_185;
  reg  [6:0]  casez_tmp_186;
  reg  [1:0]  casez_tmp_187;
  reg         casez_tmp_188;
  reg         casez_tmp_189;
  reg         casez_tmp_190;
  reg  [6:0]  casez_tmp_191;
  reg  [4:0]  casez_tmp_192;
  reg  [6:0]  casez_tmp_193;
  reg         casez_tmp_194;
  reg         casez_tmp_195;
  reg  [1:0]  casez_tmp_196;
  reg  [19:0] casez_tmp_197;
  reg  [1:0]  casez_tmp_198;
  reg  [63:0] casez_tmp_199;
  reg  [63:0] casez_tmp_200;
  reg  [1:0]  casez_tmp_201;
  reg  [1:0]  casez_tmp_202;
  reg         casez_tmp_203;
  reg  [6:0]  casez_tmp_204;
  reg  [6:0]  casez_tmp_205;
  reg  [4:0]  casez_tmp_206;
  reg  [4:0]  casez_tmp_207;
  reg  [6:0]  casez_tmp_208;
  reg         casez_tmp_209;
  reg         casez_tmp_210;
  reg         casez_tmp_211;
  reg         casez_tmp_212;
  reg  [1:0]  casez_tmp_213;
  reg  [6:0]  casez_tmp_214;
  reg  [19:0] casez_tmp_215;
  reg  [6:0]  casez_tmp_216;
  reg  [4:0]  casez_tmp_217;
  reg  [4:0]  casez_tmp_218;
  reg  [6:0]  casez_tmp_219;
  reg  [1:0]  casez_tmp_220;
  reg         casez_tmp_221;
  reg         casez_tmp_222;
  reg         casez_tmp_223;
  reg  [6:0]  casez_tmp_224;
  reg  [4:0]  casez_tmp_225;
  reg  [6:0]  casez_tmp_226;
  reg         casez_tmp_227;
  reg         casez_tmp_228;
  reg  [1:0]  casez_tmp_229;
  reg  [19:0] casez_tmp_230;
  reg  [1:0]  casez_tmp_231;
  reg  [63:0] casez_tmp_232;
  reg  [63:0] casez_tmp_233;
  reg  [1:0]  casez_tmp_234;
  reg  [1:0]  casez_tmp_235;
  reg         casez_tmp_236;
  reg  [6:0]  casez_tmp_237;
  reg  [6:0]  casez_tmp_238;
  reg  [4:0]  casez_tmp_239;
  reg  [4:0]  casez_tmp_240;
  reg  [6:0]  casez_tmp_241;
  reg         casez_tmp_242;
  reg         casez_tmp_243;
  reg         casez_tmp_244;
  reg         casez_tmp_245;
  reg  [2:0]  casez_tmp_246;
  reg         ldq_0_valid;
  reg  [6:0]  ldq_0_bits_uop_uopc;
  reg  [19:0] ldq_0_bits_uop_br_mask;
  reg  [6:0]  ldq_0_bits_uop_rob_idx;
  reg  [4:0]  ldq_0_bits_uop_ldq_idx;
  reg  [4:0]  ldq_0_bits_uop_stq_idx;
  reg  [6:0]  ldq_0_bits_uop_pdst;
  reg  [4:0]  ldq_0_bits_uop_mem_cmd;
  reg  [1:0]  ldq_0_bits_uop_mem_size;
  reg         ldq_0_bits_uop_mem_signed;
  reg         ldq_0_bits_uop_is_amo;
  reg         ldq_0_bits_uop_uses_ldq;
  reg         ldq_0_bits_uop_uses_stq;
  reg  [1:0]  ldq_0_bits_uop_dst_rtype;
  reg         ldq_0_bits_uop_fp_val;
  reg         ldq_0_bits_addr_valid;
  reg  [39:0] ldq_0_bits_addr_bits;
  reg         ldq_0_bits_addr_is_virtual;
  reg         ldq_0_bits_addr_is_uncacheable;
  reg         ldq_0_bits_executed;
  reg         ldq_0_bits_succeeded;
  reg         ldq_0_bits_order_fail;
  reg         ldq_0_bits_observed;
  reg  [31:0] ldq_0_bits_st_dep_mask;
  reg  [4:0]  ldq_0_bits_youngest_stq_idx;
  reg         ldq_0_bits_forward_std_val;
  reg  [4:0]  ldq_0_bits_forward_stq_idx;
  reg         ldq_1_valid;
  reg  [6:0]  ldq_1_bits_uop_uopc;
  reg  [19:0] ldq_1_bits_uop_br_mask;
  reg  [6:0]  ldq_1_bits_uop_rob_idx;
  reg  [4:0]  ldq_1_bits_uop_ldq_idx;
  reg  [4:0]  ldq_1_bits_uop_stq_idx;
  reg  [6:0]  ldq_1_bits_uop_pdst;
  reg  [4:0]  ldq_1_bits_uop_mem_cmd;
  reg  [1:0]  ldq_1_bits_uop_mem_size;
  reg         ldq_1_bits_uop_mem_signed;
  reg         ldq_1_bits_uop_is_amo;
  reg         ldq_1_bits_uop_uses_ldq;
  reg         ldq_1_bits_uop_uses_stq;
  reg  [1:0]  ldq_1_bits_uop_dst_rtype;
  reg         ldq_1_bits_uop_fp_val;
  reg         ldq_1_bits_addr_valid;
  reg  [39:0] ldq_1_bits_addr_bits;
  reg         ldq_1_bits_addr_is_virtual;
  reg         ldq_1_bits_addr_is_uncacheable;
  reg         ldq_1_bits_executed;
  reg         ldq_1_bits_succeeded;
  reg         ldq_1_bits_order_fail;
  reg         ldq_1_bits_observed;
  reg  [31:0] ldq_1_bits_st_dep_mask;
  reg  [4:0]  ldq_1_bits_youngest_stq_idx;
  reg         ldq_1_bits_forward_std_val;
  reg  [4:0]  ldq_1_bits_forward_stq_idx;
  reg         ldq_2_valid;
  reg  [6:0]  ldq_2_bits_uop_uopc;
  reg  [19:0] ldq_2_bits_uop_br_mask;
  reg  [6:0]  ldq_2_bits_uop_rob_idx;
  reg  [4:0]  ldq_2_bits_uop_ldq_idx;
  reg  [4:0]  ldq_2_bits_uop_stq_idx;
  reg  [6:0]  ldq_2_bits_uop_pdst;
  reg  [4:0]  ldq_2_bits_uop_mem_cmd;
  reg  [1:0]  ldq_2_bits_uop_mem_size;
  reg         ldq_2_bits_uop_mem_signed;
  reg         ldq_2_bits_uop_is_amo;
  reg         ldq_2_bits_uop_uses_ldq;
  reg         ldq_2_bits_uop_uses_stq;
  reg  [1:0]  ldq_2_bits_uop_dst_rtype;
  reg         ldq_2_bits_uop_fp_val;
  reg         ldq_2_bits_addr_valid;
  reg  [39:0] ldq_2_bits_addr_bits;
  reg         ldq_2_bits_addr_is_virtual;
  reg         ldq_2_bits_addr_is_uncacheable;
  reg         ldq_2_bits_executed;
  reg         ldq_2_bits_succeeded;
  reg         ldq_2_bits_order_fail;
  reg         ldq_2_bits_observed;
  reg  [31:0] ldq_2_bits_st_dep_mask;
  reg  [4:0]  ldq_2_bits_youngest_stq_idx;
  reg         ldq_2_bits_forward_std_val;
  reg  [4:0]  ldq_2_bits_forward_stq_idx;
  reg         ldq_3_valid;
  reg  [6:0]  ldq_3_bits_uop_uopc;
  reg  [19:0] ldq_3_bits_uop_br_mask;
  reg  [6:0]  ldq_3_bits_uop_rob_idx;
  reg  [4:0]  ldq_3_bits_uop_ldq_idx;
  reg  [4:0]  ldq_3_bits_uop_stq_idx;
  reg  [6:0]  ldq_3_bits_uop_pdst;
  reg  [4:0]  ldq_3_bits_uop_mem_cmd;
  reg  [1:0]  ldq_3_bits_uop_mem_size;
  reg         ldq_3_bits_uop_mem_signed;
  reg         ldq_3_bits_uop_is_amo;
  reg         ldq_3_bits_uop_uses_ldq;
  reg         ldq_3_bits_uop_uses_stq;
  reg  [1:0]  ldq_3_bits_uop_dst_rtype;
  reg         ldq_3_bits_uop_fp_val;
  reg         ldq_3_bits_addr_valid;
  reg  [39:0] ldq_3_bits_addr_bits;
  reg         ldq_3_bits_addr_is_virtual;
  reg         ldq_3_bits_addr_is_uncacheable;
  reg         ldq_3_bits_executed;
  reg         ldq_3_bits_succeeded;
  reg         ldq_3_bits_order_fail;
  reg         ldq_3_bits_observed;
  reg  [31:0] ldq_3_bits_st_dep_mask;
  reg  [4:0]  ldq_3_bits_youngest_stq_idx;
  reg         ldq_3_bits_forward_std_val;
  reg  [4:0]  ldq_3_bits_forward_stq_idx;
  reg         ldq_4_valid;
  reg  [6:0]  ldq_4_bits_uop_uopc;
  reg  [19:0] ldq_4_bits_uop_br_mask;
  reg  [6:0]  ldq_4_bits_uop_rob_idx;
  reg  [4:0]  ldq_4_bits_uop_ldq_idx;
  reg  [4:0]  ldq_4_bits_uop_stq_idx;
  reg  [6:0]  ldq_4_bits_uop_pdst;
  reg  [4:0]  ldq_4_bits_uop_mem_cmd;
  reg  [1:0]  ldq_4_bits_uop_mem_size;
  reg         ldq_4_bits_uop_mem_signed;
  reg         ldq_4_bits_uop_is_amo;
  reg         ldq_4_bits_uop_uses_ldq;
  reg         ldq_4_bits_uop_uses_stq;
  reg  [1:0]  ldq_4_bits_uop_dst_rtype;
  reg         ldq_4_bits_uop_fp_val;
  reg         ldq_4_bits_addr_valid;
  reg  [39:0] ldq_4_bits_addr_bits;
  reg         ldq_4_bits_addr_is_virtual;
  reg         ldq_4_bits_addr_is_uncacheable;
  reg         ldq_4_bits_executed;
  reg         ldq_4_bits_succeeded;
  reg         ldq_4_bits_order_fail;
  reg         ldq_4_bits_observed;
  reg  [31:0] ldq_4_bits_st_dep_mask;
  reg  [4:0]  ldq_4_bits_youngest_stq_idx;
  reg         ldq_4_bits_forward_std_val;
  reg  [4:0]  ldq_4_bits_forward_stq_idx;
  reg         ldq_5_valid;
  reg  [6:0]  ldq_5_bits_uop_uopc;
  reg  [19:0] ldq_5_bits_uop_br_mask;
  reg  [6:0]  ldq_5_bits_uop_rob_idx;
  reg  [4:0]  ldq_5_bits_uop_ldq_idx;
  reg  [4:0]  ldq_5_bits_uop_stq_idx;
  reg  [6:0]  ldq_5_bits_uop_pdst;
  reg  [4:0]  ldq_5_bits_uop_mem_cmd;
  reg  [1:0]  ldq_5_bits_uop_mem_size;
  reg         ldq_5_bits_uop_mem_signed;
  reg         ldq_5_bits_uop_is_amo;
  reg         ldq_5_bits_uop_uses_ldq;
  reg         ldq_5_bits_uop_uses_stq;
  reg  [1:0]  ldq_5_bits_uop_dst_rtype;
  reg         ldq_5_bits_uop_fp_val;
  reg         ldq_5_bits_addr_valid;
  reg  [39:0] ldq_5_bits_addr_bits;
  reg         ldq_5_bits_addr_is_virtual;
  reg         ldq_5_bits_addr_is_uncacheable;
  reg         ldq_5_bits_executed;
  reg         ldq_5_bits_succeeded;
  reg         ldq_5_bits_order_fail;
  reg         ldq_5_bits_observed;
  reg  [31:0] ldq_5_bits_st_dep_mask;
  reg  [4:0]  ldq_5_bits_youngest_stq_idx;
  reg         ldq_5_bits_forward_std_val;
  reg  [4:0]  ldq_5_bits_forward_stq_idx;
  reg         ldq_6_valid;
  reg  [6:0]  ldq_6_bits_uop_uopc;
  reg  [19:0] ldq_6_bits_uop_br_mask;
  reg  [6:0]  ldq_6_bits_uop_rob_idx;
  reg  [4:0]  ldq_6_bits_uop_ldq_idx;
  reg  [4:0]  ldq_6_bits_uop_stq_idx;
  reg  [6:0]  ldq_6_bits_uop_pdst;
  reg  [4:0]  ldq_6_bits_uop_mem_cmd;
  reg  [1:0]  ldq_6_bits_uop_mem_size;
  reg         ldq_6_bits_uop_mem_signed;
  reg         ldq_6_bits_uop_is_amo;
  reg         ldq_6_bits_uop_uses_ldq;
  reg         ldq_6_bits_uop_uses_stq;
  reg  [1:0]  ldq_6_bits_uop_dst_rtype;
  reg         ldq_6_bits_uop_fp_val;
  reg         ldq_6_bits_addr_valid;
  reg  [39:0] ldq_6_bits_addr_bits;
  reg         ldq_6_bits_addr_is_virtual;
  reg         ldq_6_bits_addr_is_uncacheable;
  reg         ldq_6_bits_executed;
  reg         ldq_6_bits_succeeded;
  reg         ldq_6_bits_order_fail;
  reg         ldq_6_bits_observed;
  reg  [31:0] ldq_6_bits_st_dep_mask;
  reg  [4:0]  ldq_6_bits_youngest_stq_idx;
  reg         ldq_6_bits_forward_std_val;
  reg  [4:0]  ldq_6_bits_forward_stq_idx;
  reg         ldq_7_valid;
  reg  [6:0]  ldq_7_bits_uop_uopc;
  reg  [19:0] ldq_7_bits_uop_br_mask;
  reg  [6:0]  ldq_7_bits_uop_rob_idx;
  reg  [4:0]  ldq_7_bits_uop_ldq_idx;
  reg  [4:0]  ldq_7_bits_uop_stq_idx;
  reg  [6:0]  ldq_7_bits_uop_pdst;
  reg  [4:0]  ldq_7_bits_uop_mem_cmd;
  reg  [1:0]  ldq_7_bits_uop_mem_size;
  reg         ldq_7_bits_uop_mem_signed;
  reg         ldq_7_bits_uop_is_amo;
  reg         ldq_7_bits_uop_uses_ldq;
  reg         ldq_7_bits_uop_uses_stq;
  reg  [1:0]  ldq_7_bits_uop_dst_rtype;
  reg         ldq_7_bits_uop_fp_val;
  reg         ldq_7_bits_addr_valid;
  reg  [39:0] ldq_7_bits_addr_bits;
  reg         ldq_7_bits_addr_is_virtual;
  reg         ldq_7_bits_addr_is_uncacheable;
  reg         ldq_7_bits_executed;
  reg         ldq_7_bits_succeeded;
  reg         ldq_7_bits_order_fail;
  reg         ldq_7_bits_observed;
  reg  [31:0] ldq_7_bits_st_dep_mask;
  reg  [4:0]  ldq_7_bits_youngest_stq_idx;
  reg         ldq_7_bits_forward_std_val;
  reg  [4:0]  ldq_7_bits_forward_stq_idx;
  reg         ldq_8_valid;
  reg  [6:0]  ldq_8_bits_uop_uopc;
  reg  [19:0] ldq_8_bits_uop_br_mask;
  reg  [6:0]  ldq_8_bits_uop_rob_idx;
  reg  [4:0]  ldq_8_bits_uop_ldq_idx;
  reg  [4:0]  ldq_8_bits_uop_stq_idx;
  reg  [6:0]  ldq_8_bits_uop_pdst;
  reg  [4:0]  ldq_8_bits_uop_mem_cmd;
  reg  [1:0]  ldq_8_bits_uop_mem_size;
  reg         ldq_8_bits_uop_mem_signed;
  reg         ldq_8_bits_uop_is_amo;
  reg         ldq_8_bits_uop_uses_ldq;
  reg         ldq_8_bits_uop_uses_stq;
  reg  [1:0]  ldq_8_bits_uop_dst_rtype;
  reg         ldq_8_bits_uop_fp_val;
  reg         ldq_8_bits_addr_valid;
  reg  [39:0] ldq_8_bits_addr_bits;
  reg         ldq_8_bits_addr_is_virtual;
  reg         ldq_8_bits_addr_is_uncacheable;
  reg         ldq_8_bits_executed;
  reg         ldq_8_bits_succeeded;
  reg         ldq_8_bits_order_fail;
  reg         ldq_8_bits_observed;
  reg  [31:0] ldq_8_bits_st_dep_mask;
  reg  [4:0]  ldq_8_bits_youngest_stq_idx;
  reg         ldq_8_bits_forward_std_val;
  reg  [4:0]  ldq_8_bits_forward_stq_idx;
  reg         ldq_9_valid;
  reg  [6:0]  ldq_9_bits_uop_uopc;
  reg  [19:0] ldq_9_bits_uop_br_mask;
  reg  [6:0]  ldq_9_bits_uop_rob_idx;
  reg  [4:0]  ldq_9_bits_uop_ldq_idx;
  reg  [4:0]  ldq_9_bits_uop_stq_idx;
  reg  [6:0]  ldq_9_bits_uop_pdst;
  reg  [4:0]  ldq_9_bits_uop_mem_cmd;
  reg  [1:0]  ldq_9_bits_uop_mem_size;
  reg         ldq_9_bits_uop_mem_signed;
  reg         ldq_9_bits_uop_is_amo;
  reg         ldq_9_bits_uop_uses_ldq;
  reg         ldq_9_bits_uop_uses_stq;
  reg  [1:0]  ldq_9_bits_uop_dst_rtype;
  reg         ldq_9_bits_uop_fp_val;
  reg         ldq_9_bits_addr_valid;
  reg  [39:0] ldq_9_bits_addr_bits;
  reg         ldq_9_bits_addr_is_virtual;
  reg         ldq_9_bits_addr_is_uncacheable;
  reg         ldq_9_bits_executed;
  reg         ldq_9_bits_succeeded;
  reg         ldq_9_bits_order_fail;
  reg         ldq_9_bits_observed;
  reg  [31:0] ldq_9_bits_st_dep_mask;
  reg  [4:0]  ldq_9_bits_youngest_stq_idx;
  reg         ldq_9_bits_forward_std_val;
  reg  [4:0]  ldq_9_bits_forward_stq_idx;
  reg         ldq_10_valid;
  reg  [6:0]  ldq_10_bits_uop_uopc;
  reg  [19:0] ldq_10_bits_uop_br_mask;
  reg  [6:0]  ldq_10_bits_uop_rob_idx;
  reg  [4:0]  ldq_10_bits_uop_ldq_idx;
  reg  [4:0]  ldq_10_bits_uop_stq_idx;
  reg  [6:0]  ldq_10_bits_uop_pdst;
  reg  [4:0]  ldq_10_bits_uop_mem_cmd;
  reg  [1:0]  ldq_10_bits_uop_mem_size;
  reg         ldq_10_bits_uop_mem_signed;
  reg         ldq_10_bits_uop_is_amo;
  reg         ldq_10_bits_uop_uses_ldq;
  reg         ldq_10_bits_uop_uses_stq;
  reg  [1:0]  ldq_10_bits_uop_dst_rtype;
  reg         ldq_10_bits_uop_fp_val;
  reg         ldq_10_bits_addr_valid;
  reg  [39:0] ldq_10_bits_addr_bits;
  reg         ldq_10_bits_addr_is_virtual;
  reg         ldq_10_bits_addr_is_uncacheable;
  reg         ldq_10_bits_executed;
  reg         ldq_10_bits_succeeded;
  reg         ldq_10_bits_order_fail;
  reg         ldq_10_bits_observed;
  reg  [31:0] ldq_10_bits_st_dep_mask;
  reg  [4:0]  ldq_10_bits_youngest_stq_idx;
  reg         ldq_10_bits_forward_std_val;
  reg  [4:0]  ldq_10_bits_forward_stq_idx;
  reg         ldq_11_valid;
  reg  [6:0]  ldq_11_bits_uop_uopc;
  reg  [19:0] ldq_11_bits_uop_br_mask;
  reg  [6:0]  ldq_11_bits_uop_rob_idx;
  reg  [4:0]  ldq_11_bits_uop_ldq_idx;
  reg  [4:0]  ldq_11_bits_uop_stq_idx;
  reg  [6:0]  ldq_11_bits_uop_pdst;
  reg  [4:0]  ldq_11_bits_uop_mem_cmd;
  reg  [1:0]  ldq_11_bits_uop_mem_size;
  reg         ldq_11_bits_uop_mem_signed;
  reg         ldq_11_bits_uop_is_amo;
  reg         ldq_11_bits_uop_uses_ldq;
  reg         ldq_11_bits_uop_uses_stq;
  reg  [1:0]  ldq_11_bits_uop_dst_rtype;
  reg         ldq_11_bits_uop_fp_val;
  reg         ldq_11_bits_addr_valid;
  reg  [39:0] ldq_11_bits_addr_bits;
  reg         ldq_11_bits_addr_is_virtual;
  reg         ldq_11_bits_addr_is_uncacheable;
  reg         ldq_11_bits_executed;
  reg         ldq_11_bits_succeeded;
  reg         ldq_11_bits_order_fail;
  reg         ldq_11_bits_observed;
  reg  [31:0] ldq_11_bits_st_dep_mask;
  reg  [4:0]  ldq_11_bits_youngest_stq_idx;
  reg         ldq_11_bits_forward_std_val;
  reg  [4:0]  ldq_11_bits_forward_stq_idx;
  reg         ldq_12_valid;
  reg  [6:0]  ldq_12_bits_uop_uopc;
  reg  [19:0] ldq_12_bits_uop_br_mask;
  reg  [6:0]  ldq_12_bits_uop_rob_idx;
  reg  [4:0]  ldq_12_bits_uop_ldq_idx;
  reg  [4:0]  ldq_12_bits_uop_stq_idx;
  reg  [6:0]  ldq_12_bits_uop_pdst;
  reg  [4:0]  ldq_12_bits_uop_mem_cmd;
  reg  [1:0]  ldq_12_bits_uop_mem_size;
  reg         ldq_12_bits_uop_mem_signed;
  reg         ldq_12_bits_uop_is_amo;
  reg         ldq_12_bits_uop_uses_ldq;
  reg         ldq_12_bits_uop_uses_stq;
  reg  [1:0]  ldq_12_bits_uop_dst_rtype;
  reg         ldq_12_bits_uop_fp_val;
  reg         ldq_12_bits_addr_valid;
  reg  [39:0] ldq_12_bits_addr_bits;
  reg         ldq_12_bits_addr_is_virtual;
  reg         ldq_12_bits_addr_is_uncacheable;
  reg         ldq_12_bits_executed;
  reg         ldq_12_bits_succeeded;
  reg         ldq_12_bits_order_fail;
  reg         ldq_12_bits_observed;
  reg  [31:0] ldq_12_bits_st_dep_mask;
  reg  [4:0]  ldq_12_bits_youngest_stq_idx;
  reg         ldq_12_bits_forward_std_val;
  reg  [4:0]  ldq_12_bits_forward_stq_idx;
  reg         ldq_13_valid;
  reg  [6:0]  ldq_13_bits_uop_uopc;
  reg  [19:0] ldq_13_bits_uop_br_mask;
  reg  [6:0]  ldq_13_bits_uop_rob_idx;
  reg  [4:0]  ldq_13_bits_uop_ldq_idx;
  reg  [4:0]  ldq_13_bits_uop_stq_idx;
  reg  [6:0]  ldq_13_bits_uop_pdst;
  reg  [4:0]  ldq_13_bits_uop_mem_cmd;
  reg  [1:0]  ldq_13_bits_uop_mem_size;
  reg         ldq_13_bits_uop_mem_signed;
  reg         ldq_13_bits_uop_is_amo;
  reg         ldq_13_bits_uop_uses_ldq;
  reg         ldq_13_bits_uop_uses_stq;
  reg  [1:0]  ldq_13_bits_uop_dst_rtype;
  reg         ldq_13_bits_uop_fp_val;
  reg         ldq_13_bits_addr_valid;
  reg  [39:0] ldq_13_bits_addr_bits;
  reg         ldq_13_bits_addr_is_virtual;
  reg         ldq_13_bits_addr_is_uncacheable;
  reg         ldq_13_bits_executed;
  reg         ldq_13_bits_succeeded;
  reg         ldq_13_bits_order_fail;
  reg         ldq_13_bits_observed;
  reg  [31:0] ldq_13_bits_st_dep_mask;
  reg  [4:0]  ldq_13_bits_youngest_stq_idx;
  reg         ldq_13_bits_forward_std_val;
  reg  [4:0]  ldq_13_bits_forward_stq_idx;
  reg         ldq_14_valid;
  reg  [6:0]  ldq_14_bits_uop_uopc;
  reg  [19:0] ldq_14_bits_uop_br_mask;
  reg  [6:0]  ldq_14_bits_uop_rob_idx;
  reg  [4:0]  ldq_14_bits_uop_ldq_idx;
  reg  [4:0]  ldq_14_bits_uop_stq_idx;
  reg  [6:0]  ldq_14_bits_uop_pdst;
  reg  [4:0]  ldq_14_bits_uop_mem_cmd;
  reg  [1:0]  ldq_14_bits_uop_mem_size;
  reg         ldq_14_bits_uop_mem_signed;
  reg         ldq_14_bits_uop_is_amo;
  reg         ldq_14_bits_uop_uses_ldq;
  reg         ldq_14_bits_uop_uses_stq;
  reg  [1:0]  ldq_14_bits_uop_dst_rtype;
  reg         ldq_14_bits_uop_fp_val;
  reg         ldq_14_bits_addr_valid;
  reg  [39:0] ldq_14_bits_addr_bits;
  reg         ldq_14_bits_addr_is_virtual;
  reg         ldq_14_bits_addr_is_uncacheable;
  reg         ldq_14_bits_executed;
  reg         ldq_14_bits_succeeded;
  reg         ldq_14_bits_order_fail;
  reg         ldq_14_bits_observed;
  reg  [31:0] ldq_14_bits_st_dep_mask;
  reg  [4:0]  ldq_14_bits_youngest_stq_idx;
  reg         ldq_14_bits_forward_std_val;
  reg  [4:0]  ldq_14_bits_forward_stq_idx;
  reg         ldq_15_valid;
  reg  [6:0]  ldq_15_bits_uop_uopc;
  reg  [19:0] ldq_15_bits_uop_br_mask;
  reg  [6:0]  ldq_15_bits_uop_rob_idx;
  reg  [4:0]  ldq_15_bits_uop_ldq_idx;
  reg  [4:0]  ldq_15_bits_uop_stq_idx;
  reg  [6:0]  ldq_15_bits_uop_pdst;
  reg  [4:0]  ldq_15_bits_uop_mem_cmd;
  reg  [1:0]  ldq_15_bits_uop_mem_size;
  reg         ldq_15_bits_uop_mem_signed;
  reg         ldq_15_bits_uop_is_amo;
  reg         ldq_15_bits_uop_uses_ldq;
  reg         ldq_15_bits_uop_uses_stq;
  reg  [1:0]  ldq_15_bits_uop_dst_rtype;
  reg         ldq_15_bits_uop_fp_val;
  reg         ldq_15_bits_addr_valid;
  reg  [39:0] ldq_15_bits_addr_bits;
  reg         ldq_15_bits_addr_is_virtual;
  reg         ldq_15_bits_addr_is_uncacheable;
  reg         ldq_15_bits_executed;
  reg         ldq_15_bits_succeeded;
  reg         ldq_15_bits_order_fail;
  reg         ldq_15_bits_observed;
  reg  [31:0] ldq_15_bits_st_dep_mask;
  reg  [4:0]  ldq_15_bits_youngest_stq_idx;
  reg         ldq_15_bits_forward_std_val;
  reg  [4:0]  ldq_15_bits_forward_stq_idx;
  reg         ldq_16_valid;
  reg  [6:0]  ldq_16_bits_uop_uopc;
  reg  [19:0] ldq_16_bits_uop_br_mask;
  reg  [6:0]  ldq_16_bits_uop_rob_idx;
  reg  [4:0]  ldq_16_bits_uop_ldq_idx;
  reg  [4:0]  ldq_16_bits_uop_stq_idx;
  reg  [6:0]  ldq_16_bits_uop_pdst;
  reg  [4:0]  ldq_16_bits_uop_mem_cmd;
  reg  [1:0]  ldq_16_bits_uop_mem_size;
  reg         ldq_16_bits_uop_mem_signed;
  reg         ldq_16_bits_uop_is_amo;
  reg         ldq_16_bits_uop_uses_ldq;
  reg         ldq_16_bits_uop_uses_stq;
  reg  [1:0]  ldq_16_bits_uop_dst_rtype;
  reg         ldq_16_bits_uop_fp_val;
  reg         ldq_16_bits_addr_valid;
  reg  [39:0] ldq_16_bits_addr_bits;
  reg         ldq_16_bits_addr_is_virtual;
  reg         ldq_16_bits_addr_is_uncacheable;
  reg         ldq_16_bits_executed;
  reg         ldq_16_bits_succeeded;
  reg         ldq_16_bits_order_fail;
  reg         ldq_16_bits_observed;
  reg  [31:0] ldq_16_bits_st_dep_mask;
  reg  [4:0]  ldq_16_bits_youngest_stq_idx;
  reg         ldq_16_bits_forward_std_val;
  reg  [4:0]  ldq_16_bits_forward_stq_idx;
  reg         ldq_17_valid;
  reg  [6:0]  ldq_17_bits_uop_uopc;
  reg  [19:0] ldq_17_bits_uop_br_mask;
  reg  [6:0]  ldq_17_bits_uop_rob_idx;
  reg  [4:0]  ldq_17_bits_uop_ldq_idx;
  reg  [4:0]  ldq_17_bits_uop_stq_idx;
  reg  [6:0]  ldq_17_bits_uop_pdst;
  reg  [4:0]  ldq_17_bits_uop_mem_cmd;
  reg  [1:0]  ldq_17_bits_uop_mem_size;
  reg         ldq_17_bits_uop_mem_signed;
  reg         ldq_17_bits_uop_is_amo;
  reg         ldq_17_bits_uop_uses_ldq;
  reg         ldq_17_bits_uop_uses_stq;
  reg  [1:0]  ldq_17_bits_uop_dst_rtype;
  reg         ldq_17_bits_uop_fp_val;
  reg         ldq_17_bits_addr_valid;
  reg  [39:0] ldq_17_bits_addr_bits;
  reg         ldq_17_bits_addr_is_virtual;
  reg         ldq_17_bits_addr_is_uncacheable;
  reg         ldq_17_bits_executed;
  reg         ldq_17_bits_succeeded;
  reg         ldq_17_bits_order_fail;
  reg         ldq_17_bits_observed;
  reg  [31:0] ldq_17_bits_st_dep_mask;
  reg  [4:0]  ldq_17_bits_youngest_stq_idx;
  reg         ldq_17_bits_forward_std_val;
  reg  [4:0]  ldq_17_bits_forward_stq_idx;
  reg         ldq_18_valid;
  reg  [6:0]  ldq_18_bits_uop_uopc;
  reg  [19:0] ldq_18_bits_uop_br_mask;
  reg  [6:0]  ldq_18_bits_uop_rob_idx;
  reg  [4:0]  ldq_18_bits_uop_ldq_idx;
  reg  [4:0]  ldq_18_bits_uop_stq_idx;
  reg  [6:0]  ldq_18_bits_uop_pdst;
  reg  [4:0]  ldq_18_bits_uop_mem_cmd;
  reg  [1:0]  ldq_18_bits_uop_mem_size;
  reg         ldq_18_bits_uop_mem_signed;
  reg         ldq_18_bits_uop_is_amo;
  reg         ldq_18_bits_uop_uses_ldq;
  reg         ldq_18_bits_uop_uses_stq;
  reg  [1:0]  ldq_18_bits_uop_dst_rtype;
  reg         ldq_18_bits_uop_fp_val;
  reg         ldq_18_bits_addr_valid;
  reg  [39:0] ldq_18_bits_addr_bits;
  reg         ldq_18_bits_addr_is_virtual;
  reg         ldq_18_bits_addr_is_uncacheable;
  reg         ldq_18_bits_executed;
  reg         ldq_18_bits_succeeded;
  reg         ldq_18_bits_order_fail;
  reg         ldq_18_bits_observed;
  reg  [31:0] ldq_18_bits_st_dep_mask;
  reg  [4:0]  ldq_18_bits_youngest_stq_idx;
  reg         ldq_18_bits_forward_std_val;
  reg  [4:0]  ldq_18_bits_forward_stq_idx;
  reg         ldq_19_valid;
  reg  [6:0]  ldq_19_bits_uop_uopc;
  reg  [19:0] ldq_19_bits_uop_br_mask;
  reg  [6:0]  ldq_19_bits_uop_rob_idx;
  reg  [4:0]  ldq_19_bits_uop_ldq_idx;
  reg  [4:0]  ldq_19_bits_uop_stq_idx;
  reg  [6:0]  ldq_19_bits_uop_pdst;
  reg  [4:0]  ldq_19_bits_uop_mem_cmd;
  reg  [1:0]  ldq_19_bits_uop_mem_size;
  reg         ldq_19_bits_uop_mem_signed;
  reg         ldq_19_bits_uop_is_amo;
  reg         ldq_19_bits_uop_uses_ldq;
  reg         ldq_19_bits_uop_uses_stq;
  reg  [1:0]  ldq_19_bits_uop_dst_rtype;
  reg         ldq_19_bits_uop_fp_val;
  reg         ldq_19_bits_addr_valid;
  reg  [39:0] ldq_19_bits_addr_bits;
  reg         ldq_19_bits_addr_is_virtual;
  reg         ldq_19_bits_addr_is_uncacheable;
  reg         ldq_19_bits_executed;
  reg         ldq_19_bits_succeeded;
  reg         ldq_19_bits_order_fail;
  reg         ldq_19_bits_observed;
  reg  [31:0] ldq_19_bits_st_dep_mask;
  reg  [4:0]  ldq_19_bits_youngest_stq_idx;
  reg         ldq_19_bits_forward_std_val;
  reg  [4:0]  ldq_19_bits_forward_stq_idx;
  reg         ldq_20_valid;
  reg  [6:0]  ldq_20_bits_uop_uopc;
  reg  [19:0] ldq_20_bits_uop_br_mask;
  reg  [6:0]  ldq_20_bits_uop_rob_idx;
  reg  [4:0]  ldq_20_bits_uop_ldq_idx;
  reg  [4:0]  ldq_20_bits_uop_stq_idx;
  reg  [6:0]  ldq_20_bits_uop_pdst;
  reg  [4:0]  ldq_20_bits_uop_mem_cmd;
  reg  [1:0]  ldq_20_bits_uop_mem_size;
  reg         ldq_20_bits_uop_mem_signed;
  reg         ldq_20_bits_uop_is_amo;
  reg         ldq_20_bits_uop_uses_ldq;
  reg         ldq_20_bits_uop_uses_stq;
  reg  [1:0]  ldq_20_bits_uop_dst_rtype;
  reg         ldq_20_bits_uop_fp_val;
  reg         ldq_20_bits_addr_valid;
  reg  [39:0] ldq_20_bits_addr_bits;
  reg         ldq_20_bits_addr_is_virtual;
  reg         ldq_20_bits_addr_is_uncacheable;
  reg         ldq_20_bits_executed;
  reg         ldq_20_bits_succeeded;
  reg         ldq_20_bits_order_fail;
  reg         ldq_20_bits_observed;
  reg  [31:0] ldq_20_bits_st_dep_mask;
  reg  [4:0]  ldq_20_bits_youngest_stq_idx;
  reg         ldq_20_bits_forward_std_val;
  reg  [4:0]  ldq_20_bits_forward_stq_idx;
  reg         ldq_21_valid;
  reg  [6:0]  ldq_21_bits_uop_uopc;
  reg  [19:0] ldq_21_bits_uop_br_mask;
  reg  [6:0]  ldq_21_bits_uop_rob_idx;
  reg  [4:0]  ldq_21_bits_uop_ldq_idx;
  reg  [4:0]  ldq_21_bits_uop_stq_idx;
  reg  [6:0]  ldq_21_bits_uop_pdst;
  reg  [4:0]  ldq_21_bits_uop_mem_cmd;
  reg  [1:0]  ldq_21_bits_uop_mem_size;
  reg         ldq_21_bits_uop_mem_signed;
  reg         ldq_21_bits_uop_is_amo;
  reg         ldq_21_bits_uop_uses_ldq;
  reg         ldq_21_bits_uop_uses_stq;
  reg  [1:0]  ldq_21_bits_uop_dst_rtype;
  reg         ldq_21_bits_uop_fp_val;
  reg         ldq_21_bits_addr_valid;
  reg  [39:0] ldq_21_bits_addr_bits;
  reg         ldq_21_bits_addr_is_virtual;
  reg         ldq_21_bits_addr_is_uncacheable;
  reg         ldq_21_bits_executed;
  reg         ldq_21_bits_succeeded;
  reg         ldq_21_bits_order_fail;
  reg         ldq_21_bits_observed;
  reg  [31:0] ldq_21_bits_st_dep_mask;
  reg  [4:0]  ldq_21_bits_youngest_stq_idx;
  reg         ldq_21_bits_forward_std_val;
  reg  [4:0]  ldq_21_bits_forward_stq_idx;
  reg         ldq_22_valid;
  reg  [6:0]  ldq_22_bits_uop_uopc;
  reg  [19:0] ldq_22_bits_uop_br_mask;
  reg  [6:0]  ldq_22_bits_uop_rob_idx;
  reg  [4:0]  ldq_22_bits_uop_ldq_idx;
  reg  [4:0]  ldq_22_bits_uop_stq_idx;
  reg  [6:0]  ldq_22_bits_uop_pdst;
  reg  [4:0]  ldq_22_bits_uop_mem_cmd;
  reg  [1:0]  ldq_22_bits_uop_mem_size;
  reg         ldq_22_bits_uop_mem_signed;
  reg         ldq_22_bits_uop_is_amo;
  reg         ldq_22_bits_uop_uses_ldq;
  reg         ldq_22_bits_uop_uses_stq;
  reg  [1:0]  ldq_22_bits_uop_dst_rtype;
  reg         ldq_22_bits_uop_fp_val;
  reg         ldq_22_bits_addr_valid;
  reg  [39:0] ldq_22_bits_addr_bits;
  reg         ldq_22_bits_addr_is_virtual;
  reg         ldq_22_bits_addr_is_uncacheable;
  reg         ldq_22_bits_executed;
  reg         ldq_22_bits_succeeded;
  reg         ldq_22_bits_order_fail;
  reg         ldq_22_bits_observed;
  reg  [31:0] ldq_22_bits_st_dep_mask;
  reg  [4:0]  ldq_22_bits_youngest_stq_idx;
  reg         ldq_22_bits_forward_std_val;
  reg  [4:0]  ldq_22_bits_forward_stq_idx;
  reg         ldq_23_valid;
  reg  [6:0]  ldq_23_bits_uop_uopc;
  reg  [19:0] ldq_23_bits_uop_br_mask;
  reg  [6:0]  ldq_23_bits_uop_rob_idx;
  reg  [4:0]  ldq_23_bits_uop_ldq_idx;
  reg  [4:0]  ldq_23_bits_uop_stq_idx;
  reg  [6:0]  ldq_23_bits_uop_pdst;
  reg  [4:0]  ldq_23_bits_uop_mem_cmd;
  reg  [1:0]  ldq_23_bits_uop_mem_size;
  reg         ldq_23_bits_uop_mem_signed;
  reg         ldq_23_bits_uop_is_amo;
  reg         ldq_23_bits_uop_uses_ldq;
  reg         ldq_23_bits_uop_uses_stq;
  reg  [1:0]  ldq_23_bits_uop_dst_rtype;
  reg         ldq_23_bits_uop_fp_val;
  reg         ldq_23_bits_addr_valid;
  reg  [39:0] ldq_23_bits_addr_bits;
  reg         ldq_23_bits_addr_is_virtual;
  reg         ldq_23_bits_addr_is_uncacheable;
  reg         ldq_23_bits_executed;
  reg         ldq_23_bits_succeeded;
  reg         ldq_23_bits_order_fail;
  reg         ldq_23_bits_observed;
  reg  [31:0] ldq_23_bits_st_dep_mask;
  reg  [4:0]  ldq_23_bits_youngest_stq_idx;
  reg         ldq_23_bits_forward_std_val;
  reg  [4:0]  ldq_23_bits_forward_stq_idx;
  reg         ldq_24_valid;
  reg  [6:0]  ldq_24_bits_uop_uopc;
  reg  [19:0] ldq_24_bits_uop_br_mask;
  reg  [6:0]  ldq_24_bits_uop_rob_idx;
  reg  [4:0]  ldq_24_bits_uop_ldq_idx;
  reg  [4:0]  ldq_24_bits_uop_stq_idx;
  reg  [6:0]  ldq_24_bits_uop_pdst;
  reg  [4:0]  ldq_24_bits_uop_mem_cmd;
  reg  [1:0]  ldq_24_bits_uop_mem_size;
  reg         ldq_24_bits_uop_mem_signed;
  reg         ldq_24_bits_uop_is_amo;
  reg         ldq_24_bits_uop_uses_ldq;
  reg         ldq_24_bits_uop_uses_stq;
  reg  [1:0]  ldq_24_bits_uop_dst_rtype;
  reg         ldq_24_bits_uop_fp_val;
  reg         ldq_24_bits_addr_valid;
  reg  [39:0] ldq_24_bits_addr_bits;
  reg         ldq_24_bits_addr_is_virtual;
  reg         ldq_24_bits_addr_is_uncacheable;
  reg         ldq_24_bits_executed;
  reg         ldq_24_bits_succeeded;
  reg         ldq_24_bits_order_fail;
  reg         ldq_24_bits_observed;
  reg  [31:0] ldq_24_bits_st_dep_mask;
  reg  [4:0]  ldq_24_bits_youngest_stq_idx;
  reg         ldq_24_bits_forward_std_val;
  reg  [4:0]  ldq_24_bits_forward_stq_idx;
  reg         ldq_25_valid;
  reg  [6:0]  ldq_25_bits_uop_uopc;
  reg  [19:0] ldq_25_bits_uop_br_mask;
  reg  [6:0]  ldq_25_bits_uop_rob_idx;
  reg  [4:0]  ldq_25_bits_uop_ldq_idx;
  reg  [4:0]  ldq_25_bits_uop_stq_idx;
  reg  [6:0]  ldq_25_bits_uop_pdst;
  reg  [4:0]  ldq_25_bits_uop_mem_cmd;
  reg  [1:0]  ldq_25_bits_uop_mem_size;
  reg         ldq_25_bits_uop_mem_signed;
  reg         ldq_25_bits_uop_is_amo;
  reg         ldq_25_bits_uop_uses_ldq;
  reg         ldq_25_bits_uop_uses_stq;
  reg  [1:0]  ldq_25_bits_uop_dst_rtype;
  reg         ldq_25_bits_uop_fp_val;
  reg         ldq_25_bits_addr_valid;
  reg  [39:0] ldq_25_bits_addr_bits;
  reg         ldq_25_bits_addr_is_virtual;
  reg         ldq_25_bits_addr_is_uncacheable;
  reg         ldq_25_bits_executed;
  reg         ldq_25_bits_succeeded;
  reg         ldq_25_bits_order_fail;
  reg         ldq_25_bits_observed;
  reg  [31:0] ldq_25_bits_st_dep_mask;
  reg  [4:0]  ldq_25_bits_youngest_stq_idx;
  reg         ldq_25_bits_forward_std_val;
  reg  [4:0]  ldq_25_bits_forward_stq_idx;
  reg         ldq_26_valid;
  reg  [6:0]  ldq_26_bits_uop_uopc;
  reg  [19:0] ldq_26_bits_uop_br_mask;
  reg  [6:0]  ldq_26_bits_uop_rob_idx;
  reg  [4:0]  ldq_26_bits_uop_ldq_idx;
  reg  [4:0]  ldq_26_bits_uop_stq_idx;
  reg  [6:0]  ldq_26_bits_uop_pdst;
  reg  [4:0]  ldq_26_bits_uop_mem_cmd;
  reg  [1:0]  ldq_26_bits_uop_mem_size;
  reg         ldq_26_bits_uop_mem_signed;
  reg         ldq_26_bits_uop_is_amo;
  reg         ldq_26_bits_uop_uses_ldq;
  reg         ldq_26_bits_uop_uses_stq;
  reg  [1:0]  ldq_26_bits_uop_dst_rtype;
  reg         ldq_26_bits_uop_fp_val;
  reg         ldq_26_bits_addr_valid;
  reg  [39:0] ldq_26_bits_addr_bits;
  reg         ldq_26_bits_addr_is_virtual;
  reg         ldq_26_bits_addr_is_uncacheable;
  reg         ldq_26_bits_executed;
  reg         ldq_26_bits_succeeded;
  reg         ldq_26_bits_order_fail;
  reg         ldq_26_bits_observed;
  reg  [31:0] ldq_26_bits_st_dep_mask;
  reg  [4:0]  ldq_26_bits_youngest_stq_idx;
  reg         ldq_26_bits_forward_std_val;
  reg  [4:0]  ldq_26_bits_forward_stq_idx;
  reg         ldq_27_valid;
  reg  [6:0]  ldq_27_bits_uop_uopc;
  reg  [19:0] ldq_27_bits_uop_br_mask;
  reg  [6:0]  ldq_27_bits_uop_rob_idx;
  reg  [4:0]  ldq_27_bits_uop_ldq_idx;
  reg  [4:0]  ldq_27_bits_uop_stq_idx;
  reg  [6:0]  ldq_27_bits_uop_pdst;
  reg  [4:0]  ldq_27_bits_uop_mem_cmd;
  reg  [1:0]  ldq_27_bits_uop_mem_size;
  reg         ldq_27_bits_uop_mem_signed;
  reg         ldq_27_bits_uop_is_amo;
  reg         ldq_27_bits_uop_uses_ldq;
  reg         ldq_27_bits_uop_uses_stq;
  reg  [1:0]  ldq_27_bits_uop_dst_rtype;
  reg         ldq_27_bits_uop_fp_val;
  reg         ldq_27_bits_addr_valid;
  reg  [39:0] ldq_27_bits_addr_bits;
  reg         ldq_27_bits_addr_is_virtual;
  reg         ldq_27_bits_addr_is_uncacheable;
  reg         ldq_27_bits_executed;
  reg         ldq_27_bits_succeeded;
  reg         ldq_27_bits_order_fail;
  reg         ldq_27_bits_observed;
  reg  [31:0] ldq_27_bits_st_dep_mask;
  reg  [4:0]  ldq_27_bits_youngest_stq_idx;
  reg         ldq_27_bits_forward_std_val;
  reg  [4:0]  ldq_27_bits_forward_stq_idx;
  reg         ldq_28_valid;
  reg  [6:0]  ldq_28_bits_uop_uopc;
  reg  [19:0] ldq_28_bits_uop_br_mask;
  reg  [6:0]  ldq_28_bits_uop_rob_idx;
  reg  [4:0]  ldq_28_bits_uop_ldq_idx;
  reg  [4:0]  ldq_28_bits_uop_stq_idx;
  reg  [6:0]  ldq_28_bits_uop_pdst;
  reg  [4:0]  ldq_28_bits_uop_mem_cmd;
  reg  [1:0]  ldq_28_bits_uop_mem_size;
  reg         ldq_28_bits_uop_mem_signed;
  reg         ldq_28_bits_uop_is_amo;
  reg         ldq_28_bits_uop_uses_ldq;
  reg         ldq_28_bits_uop_uses_stq;
  reg  [1:0]  ldq_28_bits_uop_dst_rtype;
  reg         ldq_28_bits_uop_fp_val;
  reg         ldq_28_bits_addr_valid;
  reg  [39:0] ldq_28_bits_addr_bits;
  reg         ldq_28_bits_addr_is_virtual;
  reg         ldq_28_bits_addr_is_uncacheable;
  reg         ldq_28_bits_executed;
  reg         ldq_28_bits_succeeded;
  reg         ldq_28_bits_order_fail;
  reg         ldq_28_bits_observed;
  reg  [31:0] ldq_28_bits_st_dep_mask;
  reg  [4:0]  ldq_28_bits_youngest_stq_idx;
  reg         ldq_28_bits_forward_std_val;
  reg  [4:0]  ldq_28_bits_forward_stq_idx;
  reg         ldq_29_valid;
  reg  [6:0]  ldq_29_bits_uop_uopc;
  reg  [19:0] ldq_29_bits_uop_br_mask;
  reg  [6:0]  ldq_29_bits_uop_rob_idx;
  reg  [4:0]  ldq_29_bits_uop_ldq_idx;
  reg  [4:0]  ldq_29_bits_uop_stq_idx;
  reg  [6:0]  ldq_29_bits_uop_pdst;
  reg  [4:0]  ldq_29_bits_uop_mem_cmd;
  reg  [1:0]  ldq_29_bits_uop_mem_size;
  reg         ldq_29_bits_uop_mem_signed;
  reg         ldq_29_bits_uop_is_amo;
  reg         ldq_29_bits_uop_uses_ldq;
  reg         ldq_29_bits_uop_uses_stq;
  reg  [1:0]  ldq_29_bits_uop_dst_rtype;
  reg         ldq_29_bits_uop_fp_val;
  reg         ldq_29_bits_addr_valid;
  reg  [39:0] ldq_29_bits_addr_bits;
  reg         ldq_29_bits_addr_is_virtual;
  reg         ldq_29_bits_addr_is_uncacheable;
  reg         ldq_29_bits_executed;
  reg         ldq_29_bits_succeeded;
  reg         ldq_29_bits_order_fail;
  reg         ldq_29_bits_observed;
  reg  [31:0] ldq_29_bits_st_dep_mask;
  reg  [4:0]  ldq_29_bits_youngest_stq_idx;
  reg         ldq_29_bits_forward_std_val;
  reg  [4:0]  ldq_29_bits_forward_stq_idx;
  reg         ldq_30_valid;
  reg  [6:0]  ldq_30_bits_uop_uopc;
  reg  [19:0] ldq_30_bits_uop_br_mask;
  reg  [6:0]  ldq_30_bits_uop_rob_idx;
  reg  [4:0]  ldq_30_bits_uop_ldq_idx;
  reg  [4:0]  ldq_30_bits_uop_stq_idx;
  reg  [6:0]  ldq_30_bits_uop_pdst;
  reg  [4:0]  ldq_30_bits_uop_mem_cmd;
  reg  [1:0]  ldq_30_bits_uop_mem_size;
  reg         ldq_30_bits_uop_mem_signed;
  reg         ldq_30_bits_uop_is_amo;
  reg         ldq_30_bits_uop_uses_ldq;
  reg         ldq_30_bits_uop_uses_stq;
  reg  [1:0]  ldq_30_bits_uop_dst_rtype;
  reg         ldq_30_bits_uop_fp_val;
  reg         ldq_30_bits_addr_valid;
  reg  [39:0] ldq_30_bits_addr_bits;
  reg         ldq_30_bits_addr_is_virtual;
  reg         ldq_30_bits_addr_is_uncacheable;
  reg         ldq_30_bits_executed;
  reg         ldq_30_bits_succeeded;
  reg         ldq_30_bits_order_fail;
  reg         ldq_30_bits_observed;
  reg  [31:0] ldq_30_bits_st_dep_mask;
  reg  [4:0]  ldq_30_bits_youngest_stq_idx;
  reg         ldq_30_bits_forward_std_val;
  reg  [4:0]  ldq_30_bits_forward_stq_idx;
  reg         ldq_31_valid;
  reg  [6:0]  ldq_31_bits_uop_uopc;
  reg  [19:0] ldq_31_bits_uop_br_mask;
  reg  [6:0]  ldq_31_bits_uop_rob_idx;
  reg  [4:0]  ldq_31_bits_uop_ldq_idx;
  reg  [4:0]  ldq_31_bits_uop_stq_idx;
  reg  [6:0]  ldq_31_bits_uop_pdst;
  reg  [4:0]  ldq_31_bits_uop_mem_cmd;
  reg  [1:0]  ldq_31_bits_uop_mem_size;
  reg         ldq_31_bits_uop_mem_signed;
  reg         ldq_31_bits_uop_is_amo;
  reg         ldq_31_bits_uop_uses_ldq;
  reg         ldq_31_bits_uop_uses_stq;
  reg  [1:0]  ldq_31_bits_uop_dst_rtype;
  reg         ldq_31_bits_uop_fp_val;
  reg         ldq_31_bits_addr_valid;
  reg  [39:0] ldq_31_bits_addr_bits;
  reg         ldq_31_bits_addr_is_virtual;
  reg         ldq_31_bits_addr_is_uncacheable;
  reg         ldq_31_bits_executed;
  reg         ldq_31_bits_succeeded;
  reg         ldq_31_bits_order_fail;
  reg         ldq_31_bits_observed;
  reg  [31:0] ldq_31_bits_st_dep_mask;
  reg  [4:0]  ldq_31_bits_youngest_stq_idx;
  reg         ldq_31_bits_forward_std_val;
  reg  [4:0]  ldq_31_bits_forward_stq_idx;
  reg         stq_0_valid;
  reg  [19:0] stq_0_bits_uop_br_mask;
  reg  [6:0]  stq_0_bits_uop_rob_idx;
  reg  [4:0]  stq_0_bits_uop_ldq_idx;
  reg  [4:0]  stq_0_bits_uop_stq_idx;
  reg  [6:0]  stq_0_bits_uop_pdst;
  reg         stq_0_bits_uop_exception;
  reg  [4:0]  stq_0_bits_uop_mem_cmd;
  reg  [1:0]  stq_0_bits_uop_mem_size;
  reg         stq_0_bits_uop_mem_signed;
  reg         stq_0_bits_uop_is_fence;
  reg         stq_0_bits_uop_is_amo;
  reg         stq_0_bits_uop_uses_ldq;
  reg         stq_0_bits_uop_uses_stq;
  reg  [1:0]  stq_0_bits_uop_dst_rtype;
  reg         stq_0_bits_addr_valid;
  reg  [39:0] stq_0_bits_addr_bits;
  reg         stq_0_bits_addr_is_virtual;
  reg         stq_0_bits_data_valid;
  reg  [63:0] stq_0_bits_data_bits;
  reg         stq_0_bits_committed;
  reg         stq_0_bits_succeeded;
  reg         stq_1_valid;
  reg  [19:0] stq_1_bits_uop_br_mask;
  reg  [6:0]  stq_1_bits_uop_rob_idx;
  reg  [4:0]  stq_1_bits_uop_ldq_idx;
  reg  [4:0]  stq_1_bits_uop_stq_idx;
  reg  [6:0]  stq_1_bits_uop_pdst;
  reg         stq_1_bits_uop_exception;
  reg  [4:0]  stq_1_bits_uop_mem_cmd;
  reg  [1:0]  stq_1_bits_uop_mem_size;
  reg         stq_1_bits_uop_mem_signed;
  reg         stq_1_bits_uop_is_fence;
  reg         stq_1_bits_uop_is_amo;
  reg         stq_1_bits_uop_uses_ldq;
  reg         stq_1_bits_uop_uses_stq;
  reg  [1:0]  stq_1_bits_uop_dst_rtype;
  reg         stq_1_bits_addr_valid;
  reg  [39:0] stq_1_bits_addr_bits;
  reg         stq_1_bits_addr_is_virtual;
  reg         stq_1_bits_data_valid;
  reg  [63:0] stq_1_bits_data_bits;
  reg         stq_1_bits_committed;
  reg         stq_1_bits_succeeded;
  reg         stq_2_valid;
  reg  [19:0] stq_2_bits_uop_br_mask;
  reg  [6:0]  stq_2_bits_uop_rob_idx;
  reg  [4:0]  stq_2_bits_uop_ldq_idx;
  reg  [4:0]  stq_2_bits_uop_stq_idx;
  reg  [6:0]  stq_2_bits_uop_pdst;
  reg         stq_2_bits_uop_exception;
  reg  [4:0]  stq_2_bits_uop_mem_cmd;
  reg  [1:0]  stq_2_bits_uop_mem_size;
  reg         stq_2_bits_uop_mem_signed;
  reg         stq_2_bits_uop_is_fence;
  reg         stq_2_bits_uop_is_amo;
  reg         stq_2_bits_uop_uses_ldq;
  reg         stq_2_bits_uop_uses_stq;
  reg  [1:0]  stq_2_bits_uop_dst_rtype;
  reg         stq_2_bits_addr_valid;
  reg  [39:0] stq_2_bits_addr_bits;
  reg         stq_2_bits_addr_is_virtual;
  reg         stq_2_bits_data_valid;
  reg  [63:0] stq_2_bits_data_bits;
  reg         stq_2_bits_committed;
  reg         stq_2_bits_succeeded;
  reg         stq_3_valid;
  reg  [19:0] stq_3_bits_uop_br_mask;
  reg  [6:0]  stq_3_bits_uop_rob_idx;
  reg  [4:0]  stq_3_bits_uop_ldq_idx;
  reg  [4:0]  stq_3_bits_uop_stq_idx;
  reg  [6:0]  stq_3_bits_uop_pdst;
  reg         stq_3_bits_uop_exception;
  reg  [4:0]  stq_3_bits_uop_mem_cmd;
  reg  [1:0]  stq_3_bits_uop_mem_size;
  reg         stq_3_bits_uop_mem_signed;
  reg         stq_3_bits_uop_is_fence;
  reg         stq_3_bits_uop_is_amo;
  reg         stq_3_bits_uop_uses_ldq;
  reg         stq_3_bits_uop_uses_stq;
  reg  [1:0]  stq_3_bits_uop_dst_rtype;
  reg         stq_3_bits_addr_valid;
  reg  [39:0] stq_3_bits_addr_bits;
  reg         stq_3_bits_addr_is_virtual;
  reg         stq_3_bits_data_valid;
  reg  [63:0] stq_3_bits_data_bits;
  reg         stq_3_bits_committed;
  reg         stq_3_bits_succeeded;
  reg         stq_4_valid;
  reg  [19:0] stq_4_bits_uop_br_mask;
  reg  [6:0]  stq_4_bits_uop_rob_idx;
  reg  [4:0]  stq_4_bits_uop_ldq_idx;
  reg  [4:0]  stq_4_bits_uop_stq_idx;
  reg  [6:0]  stq_4_bits_uop_pdst;
  reg         stq_4_bits_uop_exception;
  reg  [4:0]  stq_4_bits_uop_mem_cmd;
  reg  [1:0]  stq_4_bits_uop_mem_size;
  reg         stq_4_bits_uop_mem_signed;
  reg         stq_4_bits_uop_is_fence;
  reg         stq_4_bits_uop_is_amo;
  reg         stq_4_bits_uop_uses_ldq;
  reg         stq_4_bits_uop_uses_stq;
  reg  [1:0]  stq_4_bits_uop_dst_rtype;
  reg         stq_4_bits_addr_valid;
  reg  [39:0] stq_4_bits_addr_bits;
  reg         stq_4_bits_addr_is_virtual;
  reg         stq_4_bits_data_valid;
  reg  [63:0] stq_4_bits_data_bits;
  reg         stq_4_bits_committed;
  reg         stq_4_bits_succeeded;
  reg         stq_5_valid;
  reg  [19:0] stq_5_bits_uop_br_mask;
  reg  [6:0]  stq_5_bits_uop_rob_idx;
  reg  [4:0]  stq_5_bits_uop_ldq_idx;
  reg  [4:0]  stq_5_bits_uop_stq_idx;
  reg  [6:0]  stq_5_bits_uop_pdst;
  reg         stq_5_bits_uop_exception;
  reg  [4:0]  stq_5_bits_uop_mem_cmd;
  reg  [1:0]  stq_5_bits_uop_mem_size;
  reg         stq_5_bits_uop_mem_signed;
  reg         stq_5_bits_uop_is_fence;
  reg         stq_5_bits_uop_is_amo;
  reg         stq_5_bits_uop_uses_ldq;
  reg         stq_5_bits_uop_uses_stq;
  reg  [1:0]  stq_5_bits_uop_dst_rtype;
  reg         stq_5_bits_addr_valid;
  reg  [39:0] stq_5_bits_addr_bits;
  reg         stq_5_bits_addr_is_virtual;
  reg         stq_5_bits_data_valid;
  reg  [63:0] stq_5_bits_data_bits;
  reg         stq_5_bits_committed;
  reg         stq_5_bits_succeeded;
  reg         stq_6_valid;
  reg  [19:0] stq_6_bits_uop_br_mask;
  reg  [6:0]  stq_6_bits_uop_rob_idx;
  reg  [4:0]  stq_6_bits_uop_ldq_idx;
  reg  [4:0]  stq_6_bits_uop_stq_idx;
  reg  [6:0]  stq_6_bits_uop_pdst;
  reg         stq_6_bits_uop_exception;
  reg  [4:0]  stq_6_bits_uop_mem_cmd;
  reg  [1:0]  stq_6_bits_uop_mem_size;
  reg         stq_6_bits_uop_mem_signed;
  reg         stq_6_bits_uop_is_fence;
  reg         stq_6_bits_uop_is_amo;
  reg         stq_6_bits_uop_uses_ldq;
  reg         stq_6_bits_uop_uses_stq;
  reg  [1:0]  stq_6_bits_uop_dst_rtype;
  reg         stq_6_bits_addr_valid;
  reg  [39:0] stq_6_bits_addr_bits;
  reg         stq_6_bits_addr_is_virtual;
  reg         stq_6_bits_data_valid;
  reg  [63:0] stq_6_bits_data_bits;
  reg         stq_6_bits_committed;
  reg         stq_6_bits_succeeded;
  reg         stq_7_valid;
  reg  [19:0] stq_7_bits_uop_br_mask;
  reg  [6:0]  stq_7_bits_uop_rob_idx;
  reg  [4:0]  stq_7_bits_uop_ldq_idx;
  reg  [4:0]  stq_7_bits_uop_stq_idx;
  reg  [6:0]  stq_7_bits_uop_pdst;
  reg         stq_7_bits_uop_exception;
  reg  [4:0]  stq_7_bits_uop_mem_cmd;
  reg  [1:0]  stq_7_bits_uop_mem_size;
  reg         stq_7_bits_uop_mem_signed;
  reg         stq_7_bits_uop_is_fence;
  reg         stq_7_bits_uop_is_amo;
  reg         stq_7_bits_uop_uses_ldq;
  reg         stq_7_bits_uop_uses_stq;
  reg  [1:0]  stq_7_bits_uop_dst_rtype;
  reg         stq_7_bits_addr_valid;
  reg  [39:0] stq_7_bits_addr_bits;
  reg         stq_7_bits_addr_is_virtual;
  reg         stq_7_bits_data_valid;
  reg  [63:0] stq_7_bits_data_bits;
  reg         stq_7_bits_committed;
  reg         stq_7_bits_succeeded;
  reg         stq_8_valid;
  reg  [19:0] stq_8_bits_uop_br_mask;
  reg  [6:0]  stq_8_bits_uop_rob_idx;
  reg  [4:0]  stq_8_bits_uop_ldq_idx;
  reg  [4:0]  stq_8_bits_uop_stq_idx;
  reg  [6:0]  stq_8_bits_uop_pdst;
  reg         stq_8_bits_uop_exception;
  reg  [4:0]  stq_8_bits_uop_mem_cmd;
  reg  [1:0]  stq_8_bits_uop_mem_size;
  reg         stq_8_bits_uop_mem_signed;
  reg         stq_8_bits_uop_is_fence;
  reg         stq_8_bits_uop_is_amo;
  reg         stq_8_bits_uop_uses_ldq;
  reg         stq_8_bits_uop_uses_stq;
  reg  [1:0]  stq_8_bits_uop_dst_rtype;
  reg         stq_8_bits_addr_valid;
  reg  [39:0] stq_8_bits_addr_bits;
  reg         stq_8_bits_addr_is_virtual;
  reg         stq_8_bits_data_valid;
  reg  [63:0] stq_8_bits_data_bits;
  reg         stq_8_bits_committed;
  reg         stq_8_bits_succeeded;
  reg         stq_9_valid;
  reg  [19:0] stq_9_bits_uop_br_mask;
  reg  [6:0]  stq_9_bits_uop_rob_idx;
  reg  [4:0]  stq_9_bits_uop_ldq_idx;
  reg  [4:0]  stq_9_bits_uop_stq_idx;
  reg  [6:0]  stq_9_bits_uop_pdst;
  reg         stq_9_bits_uop_exception;
  reg  [4:0]  stq_9_bits_uop_mem_cmd;
  reg  [1:0]  stq_9_bits_uop_mem_size;
  reg         stq_9_bits_uop_mem_signed;
  reg         stq_9_bits_uop_is_fence;
  reg         stq_9_bits_uop_is_amo;
  reg         stq_9_bits_uop_uses_ldq;
  reg         stq_9_bits_uop_uses_stq;
  reg  [1:0]  stq_9_bits_uop_dst_rtype;
  reg         stq_9_bits_addr_valid;
  reg  [39:0] stq_9_bits_addr_bits;
  reg         stq_9_bits_addr_is_virtual;
  reg         stq_9_bits_data_valid;
  reg  [63:0] stq_9_bits_data_bits;
  reg         stq_9_bits_committed;
  reg         stq_9_bits_succeeded;
  reg         stq_10_valid;
  reg  [19:0] stq_10_bits_uop_br_mask;
  reg  [6:0]  stq_10_bits_uop_rob_idx;
  reg  [4:0]  stq_10_bits_uop_ldq_idx;
  reg  [4:0]  stq_10_bits_uop_stq_idx;
  reg  [6:0]  stq_10_bits_uop_pdst;
  reg         stq_10_bits_uop_exception;
  reg  [4:0]  stq_10_bits_uop_mem_cmd;
  reg  [1:0]  stq_10_bits_uop_mem_size;
  reg         stq_10_bits_uop_mem_signed;
  reg         stq_10_bits_uop_is_fence;
  reg         stq_10_bits_uop_is_amo;
  reg         stq_10_bits_uop_uses_ldq;
  reg         stq_10_bits_uop_uses_stq;
  reg  [1:0]  stq_10_bits_uop_dst_rtype;
  reg         stq_10_bits_addr_valid;
  reg  [39:0] stq_10_bits_addr_bits;
  reg         stq_10_bits_addr_is_virtual;
  reg         stq_10_bits_data_valid;
  reg  [63:0] stq_10_bits_data_bits;
  reg         stq_10_bits_committed;
  reg         stq_10_bits_succeeded;
  reg         stq_11_valid;
  reg  [19:0] stq_11_bits_uop_br_mask;
  reg  [6:0]  stq_11_bits_uop_rob_idx;
  reg  [4:0]  stq_11_bits_uop_ldq_idx;
  reg  [4:0]  stq_11_bits_uop_stq_idx;
  reg  [6:0]  stq_11_bits_uop_pdst;
  reg         stq_11_bits_uop_exception;
  reg  [4:0]  stq_11_bits_uop_mem_cmd;
  reg  [1:0]  stq_11_bits_uop_mem_size;
  reg         stq_11_bits_uop_mem_signed;
  reg         stq_11_bits_uop_is_fence;
  reg         stq_11_bits_uop_is_amo;
  reg         stq_11_bits_uop_uses_ldq;
  reg         stq_11_bits_uop_uses_stq;
  reg  [1:0]  stq_11_bits_uop_dst_rtype;
  reg         stq_11_bits_addr_valid;
  reg  [39:0] stq_11_bits_addr_bits;
  reg         stq_11_bits_addr_is_virtual;
  reg         stq_11_bits_data_valid;
  reg  [63:0] stq_11_bits_data_bits;
  reg         stq_11_bits_committed;
  reg         stq_11_bits_succeeded;
  reg         stq_12_valid;
  reg  [19:0] stq_12_bits_uop_br_mask;
  reg  [6:0]  stq_12_bits_uop_rob_idx;
  reg  [4:0]  stq_12_bits_uop_ldq_idx;
  reg  [4:0]  stq_12_bits_uop_stq_idx;
  reg  [6:0]  stq_12_bits_uop_pdst;
  reg         stq_12_bits_uop_exception;
  reg  [4:0]  stq_12_bits_uop_mem_cmd;
  reg  [1:0]  stq_12_bits_uop_mem_size;
  reg         stq_12_bits_uop_mem_signed;
  reg         stq_12_bits_uop_is_fence;
  reg         stq_12_bits_uop_is_amo;
  reg         stq_12_bits_uop_uses_ldq;
  reg         stq_12_bits_uop_uses_stq;
  reg  [1:0]  stq_12_bits_uop_dst_rtype;
  reg         stq_12_bits_addr_valid;
  reg  [39:0] stq_12_bits_addr_bits;
  reg         stq_12_bits_addr_is_virtual;
  reg         stq_12_bits_data_valid;
  reg  [63:0] stq_12_bits_data_bits;
  reg         stq_12_bits_committed;
  reg         stq_12_bits_succeeded;
  reg         stq_13_valid;
  reg  [19:0] stq_13_bits_uop_br_mask;
  reg  [6:0]  stq_13_bits_uop_rob_idx;
  reg  [4:0]  stq_13_bits_uop_ldq_idx;
  reg  [4:0]  stq_13_bits_uop_stq_idx;
  reg  [6:0]  stq_13_bits_uop_pdst;
  reg         stq_13_bits_uop_exception;
  reg  [4:0]  stq_13_bits_uop_mem_cmd;
  reg  [1:0]  stq_13_bits_uop_mem_size;
  reg         stq_13_bits_uop_mem_signed;
  reg         stq_13_bits_uop_is_fence;
  reg         stq_13_bits_uop_is_amo;
  reg         stq_13_bits_uop_uses_ldq;
  reg         stq_13_bits_uop_uses_stq;
  reg  [1:0]  stq_13_bits_uop_dst_rtype;
  reg         stq_13_bits_addr_valid;
  reg  [39:0] stq_13_bits_addr_bits;
  reg         stq_13_bits_addr_is_virtual;
  reg         stq_13_bits_data_valid;
  reg  [63:0] stq_13_bits_data_bits;
  reg         stq_13_bits_committed;
  reg         stq_13_bits_succeeded;
  reg         stq_14_valid;
  reg  [19:0] stq_14_bits_uop_br_mask;
  reg  [6:0]  stq_14_bits_uop_rob_idx;
  reg  [4:0]  stq_14_bits_uop_ldq_idx;
  reg  [4:0]  stq_14_bits_uop_stq_idx;
  reg  [6:0]  stq_14_bits_uop_pdst;
  reg         stq_14_bits_uop_exception;
  reg  [4:0]  stq_14_bits_uop_mem_cmd;
  reg  [1:0]  stq_14_bits_uop_mem_size;
  reg         stq_14_bits_uop_mem_signed;
  reg         stq_14_bits_uop_is_fence;
  reg         stq_14_bits_uop_is_amo;
  reg         stq_14_bits_uop_uses_ldq;
  reg         stq_14_bits_uop_uses_stq;
  reg  [1:0]  stq_14_bits_uop_dst_rtype;
  reg         stq_14_bits_addr_valid;
  reg  [39:0] stq_14_bits_addr_bits;
  reg         stq_14_bits_addr_is_virtual;
  reg         stq_14_bits_data_valid;
  reg  [63:0] stq_14_bits_data_bits;
  reg         stq_14_bits_committed;
  reg         stq_14_bits_succeeded;
  reg         stq_15_valid;
  reg  [19:0] stq_15_bits_uop_br_mask;
  reg  [6:0]  stq_15_bits_uop_rob_idx;
  reg  [4:0]  stq_15_bits_uop_ldq_idx;
  reg  [4:0]  stq_15_bits_uop_stq_idx;
  reg  [6:0]  stq_15_bits_uop_pdst;
  reg         stq_15_bits_uop_exception;
  reg  [4:0]  stq_15_bits_uop_mem_cmd;
  reg  [1:0]  stq_15_bits_uop_mem_size;
  reg         stq_15_bits_uop_mem_signed;
  reg         stq_15_bits_uop_is_fence;
  reg         stq_15_bits_uop_is_amo;
  reg         stq_15_bits_uop_uses_ldq;
  reg         stq_15_bits_uop_uses_stq;
  reg  [1:0]  stq_15_bits_uop_dst_rtype;
  reg         stq_15_bits_addr_valid;
  reg  [39:0] stq_15_bits_addr_bits;
  reg         stq_15_bits_addr_is_virtual;
  reg         stq_15_bits_data_valid;
  reg  [63:0] stq_15_bits_data_bits;
  reg         stq_15_bits_committed;
  reg         stq_15_bits_succeeded;
  reg         stq_16_valid;
  reg  [19:0] stq_16_bits_uop_br_mask;
  reg  [6:0]  stq_16_bits_uop_rob_idx;
  reg  [4:0]  stq_16_bits_uop_ldq_idx;
  reg  [4:0]  stq_16_bits_uop_stq_idx;
  reg  [6:0]  stq_16_bits_uop_pdst;
  reg         stq_16_bits_uop_exception;
  reg  [4:0]  stq_16_bits_uop_mem_cmd;
  reg  [1:0]  stq_16_bits_uop_mem_size;
  reg         stq_16_bits_uop_mem_signed;
  reg         stq_16_bits_uop_is_fence;
  reg         stq_16_bits_uop_is_amo;
  reg         stq_16_bits_uop_uses_ldq;
  reg         stq_16_bits_uop_uses_stq;
  reg  [1:0]  stq_16_bits_uop_dst_rtype;
  reg         stq_16_bits_addr_valid;
  reg  [39:0] stq_16_bits_addr_bits;
  reg         stq_16_bits_addr_is_virtual;
  reg         stq_16_bits_data_valid;
  reg  [63:0] stq_16_bits_data_bits;
  reg         stq_16_bits_committed;
  reg         stq_16_bits_succeeded;
  reg         stq_17_valid;
  reg  [19:0] stq_17_bits_uop_br_mask;
  reg  [6:0]  stq_17_bits_uop_rob_idx;
  reg  [4:0]  stq_17_bits_uop_ldq_idx;
  reg  [4:0]  stq_17_bits_uop_stq_idx;
  reg  [6:0]  stq_17_bits_uop_pdst;
  reg         stq_17_bits_uop_exception;
  reg  [4:0]  stq_17_bits_uop_mem_cmd;
  reg  [1:0]  stq_17_bits_uop_mem_size;
  reg         stq_17_bits_uop_mem_signed;
  reg         stq_17_bits_uop_is_fence;
  reg         stq_17_bits_uop_is_amo;
  reg         stq_17_bits_uop_uses_ldq;
  reg         stq_17_bits_uop_uses_stq;
  reg  [1:0]  stq_17_bits_uop_dst_rtype;
  reg         stq_17_bits_addr_valid;
  reg  [39:0] stq_17_bits_addr_bits;
  reg         stq_17_bits_addr_is_virtual;
  reg         stq_17_bits_data_valid;
  reg  [63:0] stq_17_bits_data_bits;
  reg         stq_17_bits_committed;
  reg         stq_17_bits_succeeded;
  reg         stq_18_valid;
  reg  [19:0] stq_18_bits_uop_br_mask;
  reg  [6:0]  stq_18_bits_uop_rob_idx;
  reg  [4:0]  stq_18_bits_uop_ldq_idx;
  reg  [4:0]  stq_18_bits_uop_stq_idx;
  reg  [6:0]  stq_18_bits_uop_pdst;
  reg         stq_18_bits_uop_exception;
  reg  [4:0]  stq_18_bits_uop_mem_cmd;
  reg  [1:0]  stq_18_bits_uop_mem_size;
  reg         stq_18_bits_uop_mem_signed;
  reg         stq_18_bits_uop_is_fence;
  reg         stq_18_bits_uop_is_amo;
  reg         stq_18_bits_uop_uses_ldq;
  reg         stq_18_bits_uop_uses_stq;
  reg  [1:0]  stq_18_bits_uop_dst_rtype;
  reg         stq_18_bits_addr_valid;
  reg  [39:0] stq_18_bits_addr_bits;
  reg         stq_18_bits_addr_is_virtual;
  reg         stq_18_bits_data_valid;
  reg  [63:0] stq_18_bits_data_bits;
  reg         stq_18_bits_committed;
  reg         stq_18_bits_succeeded;
  reg         stq_19_valid;
  reg  [19:0] stq_19_bits_uop_br_mask;
  reg  [6:0]  stq_19_bits_uop_rob_idx;
  reg  [4:0]  stq_19_bits_uop_ldq_idx;
  reg  [4:0]  stq_19_bits_uop_stq_idx;
  reg  [6:0]  stq_19_bits_uop_pdst;
  reg         stq_19_bits_uop_exception;
  reg  [4:0]  stq_19_bits_uop_mem_cmd;
  reg  [1:0]  stq_19_bits_uop_mem_size;
  reg         stq_19_bits_uop_mem_signed;
  reg         stq_19_bits_uop_is_fence;
  reg         stq_19_bits_uop_is_amo;
  reg         stq_19_bits_uop_uses_ldq;
  reg         stq_19_bits_uop_uses_stq;
  reg  [1:0]  stq_19_bits_uop_dst_rtype;
  reg         stq_19_bits_addr_valid;
  reg  [39:0] stq_19_bits_addr_bits;
  reg         stq_19_bits_addr_is_virtual;
  reg         stq_19_bits_data_valid;
  reg  [63:0] stq_19_bits_data_bits;
  reg         stq_19_bits_committed;
  reg         stq_19_bits_succeeded;
  reg         stq_20_valid;
  reg  [19:0] stq_20_bits_uop_br_mask;
  reg  [6:0]  stq_20_bits_uop_rob_idx;
  reg  [4:0]  stq_20_bits_uop_ldq_idx;
  reg  [4:0]  stq_20_bits_uop_stq_idx;
  reg  [6:0]  stq_20_bits_uop_pdst;
  reg         stq_20_bits_uop_exception;
  reg  [4:0]  stq_20_bits_uop_mem_cmd;
  reg  [1:0]  stq_20_bits_uop_mem_size;
  reg         stq_20_bits_uop_mem_signed;
  reg         stq_20_bits_uop_is_fence;
  reg         stq_20_bits_uop_is_amo;
  reg         stq_20_bits_uop_uses_ldq;
  reg         stq_20_bits_uop_uses_stq;
  reg  [1:0]  stq_20_bits_uop_dst_rtype;
  reg         stq_20_bits_addr_valid;
  reg  [39:0] stq_20_bits_addr_bits;
  reg         stq_20_bits_addr_is_virtual;
  reg         stq_20_bits_data_valid;
  reg  [63:0] stq_20_bits_data_bits;
  reg         stq_20_bits_committed;
  reg         stq_20_bits_succeeded;
  reg         stq_21_valid;
  reg  [19:0] stq_21_bits_uop_br_mask;
  reg  [6:0]  stq_21_bits_uop_rob_idx;
  reg  [4:0]  stq_21_bits_uop_ldq_idx;
  reg  [4:0]  stq_21_bits_uop_stq_idx;
  reg  [6:0]  stq_21_bits_uop_pdst;
  reg         stq_21_bits_uop_exception;
  reg  [4:0]  stq_21_bits_uop_mem_cmd;
  reg  [1:0]  stq_21_bits_uop_mem_size;
  reg         stq_21_bits_uop_mem_signed;
  reg         stq_21_bits_uop_is_fence;
  reg         stq_21_bits_uop_is_amo;
  reg         stq_21_bits_uop_uses_ldq;
  reg         stq_21_bits_uop_uses_stq;
  reg  [1:0]  stq_21_bits_uop_dst_rtype;
  reg         stq_21_bits_addr_valid;
  reg  [39:0] stq_21_bits_addr_bits;
  reg         stq_21_bits_addr_is_virtual;
  reg         stq_21_bits_data_valid;
  reg  [63:0] stq_21_bits_data_bits;
  reg         stq_21_bits_committed;
  reg         stq_21_bits_succeeded;
  reg         stq_22_valid;
  reg  [19:0] stq_22_bits_uop_br_mask;
  reg  [6:0]  stq_22_bits_uop_rob_idx;
  reg  [4:0]  stq_22_bits_uop_ldq_idx;
  reg  [4:0]  stq_22_bits_uop_stq_idx;
  reg  [6:0]  stq_22_bits_uop_pdst;
  reg         stq_22_bits_uop_exception;
  reg  [4:0]  stq_22_bits_uop_mem_cmd;
  reg  [1:0]  stq_22_bits_uop_mem_size;
  reg         stq_22_bits_uop_mem_signed;
  reg         stq_22_bits_uop_is_fence;
  reg         stq_22_bits_uop_is_amo;
  reg         stq_22_bits_uop_uses_ldq;
  reg         stq_22_bits_uop_uses_stq;
  reg  [1:0]  stq_22_bits_uop_dst_rtype;
  reg         stq_22_bits_addr_valid;
  reg  [39:0] stq_22_bits_addr_bits;
  reg         stq_22_bits_addr_is_virtual;
  reg         stq_22_bits_data_valid;
  reg  [63:0] stq_22_bits_data_bits;
  reg         stq_22_bits_committed;
  reg         stq_22_bits_succeeded;
  reg         stq_23_valid;
  reg  [19:0] stq_23_bits_uop_br_mask;
  reg  [6:0]  stq_23_bits_uop_rob_idx;
  reg  [4:0]  stq_23_bits_uop_ldq_idx;
  reg  [4:0]  stq_23_bits_uop_stq_idx;
  reg  [6:0]  stq_23_bits_uop_pdst;
  reg         stq_23_bits_uop_exception;
  reg  [4:0]  stq_23_bits_uop_mem_cmd;
  reg  [1:0]  stq_23_bits_uop_mem_size;
  reg         stq_23_bits_uop_mem_signed;
  reg         stq_23_bits_uop_is_fence;
  reg         stq_23_bits_uop_is_amo;
  reg         stq_23_bits_uop_uses_ldq;
  reg         stq_23_bits_uop_uses_stq;
  reg  [1:0]  stq_23_bits_uop_dst_rtype;
  reg         stq_23_bits_addr_valid;
  reg  [39:0] stq_23_bits_addr_bits;
  reg         stq_23_bits_addr_is_virtual;
  reg         stq_23_bits_data_valid;
  reg  [63:0] stq_23_bits_data_bits;
  reg         stq_23_bits_committed;
  reg         stq_23_bits_succeeded;
  reg         stq_24_valid;
  reg  [19:0] stq_24_bits_uop_br_mask;
  reg  [6:0]  stq_24_bits_uop_rob_idx;
  reg  [4:0]  stq_24_bits_uop_ldq_idx;
  reg  [4:0]  stq_24_bits_uop_stq_idx;
  reg  [6:0]  stq_24_bits_uop_pdst;
  reg         stq_24_bits_uop_exception;
  reg  [4:0]  stq_24_bits_uop_mem_cmd;
  reg  [1:0]  stq_24_bits_uop_mem_size;
  reg         stq_24_bits_uop_mem_signed;
  reg         stq_24_bits_uop_is_fence;
  reg         stq_24_bits_uop_is_amo;
  reg         stq_24_bits_uop_uses_ldq;
  reg         stq_24_bits_uop_uses_stq;
  reg  [1:0]  stq_24_bits_uop_dst_rtype;
  reg         stq_24_bits_addr_valid;
  reg  [39:0] stq_24_bits_addr_bits;
  reg         stq_24_bits_addr_is_virtual;
  reg         stq_24_bits_data_valid;
  reg  [63:0] stq_24_bits_data_bits;
  reg         stq_24_bits_committed;
  reg         stq_24_bits_succeeded;
  reg         stq_25_valid;
  reg  [19:0] stq_25_bits_uop_br_mask;
  reg  [6:0]  stq_25_bits_uop_rob_idx;
  reg  [4:0]  stq_25_bits_uop_ldq_idx;
  reg  [4:0]  stq_25_bits_uop_stq_idx;
  reg  [6:0]  stq_25_bits_uop_pdst;
  reg         stq_25_bits_uop_exception;
  reg  [4:0]  stq_25_bits_uop_mem_cmd;
  reg  [1:0]  stq_25_bits_uop_mem_size;
  reg         stq_25_bits_uop_mem_signed;
  reg         stq_25_bits_uop_is_fence;
  reg         stq_25_bits_uop_is_amo;
  reg         stq_25_bits_uop_uses_ldq;
  reg         stq_25_bits_uop_uses_stq;
  reg  [1:0]  stq_25_bits_uop_dst_rtype;
  reg         stq_25_bits_addr_valid;
  reg  [39:0] stq_25_bits_addr_bits;
  reg         stq_25_bits_addr_is_virtual;
  reg         stq_25_bits_data_valid;
  reg  [63:0] stq_25_bits_data_bits;
  reg         stq_25_bits_committed;
  reg         stq_25_bits_succeeded;
  reg         stq_26_valid;
  reg  [19:0] stq_26_bits_uop_br_mask;
  reg  [6:0]  stq_26_bits_uop_rob_idx;
  reg  [4:0]  stq_26_bits_uop_ldq_idx;
  reg  [4:0]  stq_26_bits_uop_stq_idx;
  reg  [6:0]  stq_26_bits_uop_pdst;
  reg         stq_26_bits_uop_exception;
  reg  [4:0]  stq_26_bits_uop_mem_cmd;
  reg  [1:0]  stq_26_bits_uop_mem_size;
  reg         stq_26_bits_uop_mem_signed;
  reg         stq_26_bits_uop_is_fence;
  reg         stq_26_bits_uop_is_amo;
  reg         stq_26_bits_uop_uses_ldq;
  reg         stq_26_bits_uop_uses_stq;
  reg  [1:0]  stq_26_bits_uop_dst_rtype;
  reg         stq_26_bits_addr_valid;
  reg  [39:0] stq_26_bits_addr_bits;
  reg         stq_26_bits_addr_is_virtual;
  reg         stq_26_bits_data_valid;
  reg  [63:0] stq_26_bits_data_bits;
  reg         stq_26_bits_committed;
  reg         stq_26_bits_succeeded;
  reg         stq_27_valid;
  reg  [19:0] stq_27_bits_uop_br_mask;
  reg  [6:0]  stq_27_bits_uop_rob_idx;
  reg  [4:0]  stq_27_bits_uop_ldq_idx;
  reg  [4:0]  stq_27_bits_uop_stq_idx;
  reg  [6:0]  stq_27_bits_uop_pdst;
  reg         stq_27_bits_uop_exception;
  reg  [4:0]  stq_27_bits_uop_mem_cmd;
  reg  [1:0]  stq_27_bits_uop_mem_size;
  reg         stq_27_bits_uop_mem_signed;
  reg         stq_27_bits_uop_is_fence;
  reg         stq_27_bits_uop_is_amo;
  reg         stq_27_bits_uop_uses_ldq;
  reg         stq_27_bits_uop_uses_stq;
  reg  [1:0]  stq_27_bits_uop_dst_rtype;
  reg         stq_27_bits_addr_valid;
  reg  [39:0] stq_27_bits_addr_bits;
  reg         stq_27_bits_addr_is_virtual;
  reg         stq_27_bits_data_valid;
  reg  [63:0] stq_27_bits_data_bits;
  reg         stq_27_bits_committed;
  reg         stq_27_bits_succeeded;
  reg         stq_28_valid;
  reg  [19:0] stq_28_bits_uop_br_mask;
  reg  [6:0]  stq_28_bits_uop_rob_idx;
  reg  [4:0]  stq_28_bits_uop_ldq_idx;
  reg  [4:0]  stq_28_bits_uop_stq_idx;
  reg  [6:0]  stq_28_bits_uop_pdst;
  reg         stq_28_bits_uop_exception;
  reg  [4:0]  stq_28_bits_uop_mem_cmd;
  reg  [1:0]  stq_28_bits_uop_mem_size;
  reg         stq_28_bits_uop_mem_signed;
  reg         stq_28_bits_uop_is_fence;
  reg         stq_28_bits_uop_is_amo;
  reg         stq_28_bits_uop_uses_ldq;
  reg         stq_28_bits_uop_uses_stq;
  reg  [1:0]  stq_28_bits_uop_dst_rtype;
  reg         stq_28_bits_addr_valid;
  reg  [39:0] stq_28_bits_addr_bits;
  reg         stq_28_bits_addr_is_virtual;
  reg         stq_28_bits_data_valid;
  reg  [63:0] stq_28_bits_data_bits;
  reg         stq_28_bits_committed;
  reg         stq_28_bits_succeeded;
  reg         stq_29_valid;
  reg  [19:0] stq_29_bits_uop_br_mask;
  reg  [6:0]  stq_29_bits_uop_rob_idx;
  reg  [4:0]  stq_29_bits_uop_ldq_idx;
  reg  [4:0]  stq_29_bits_uop_stq_idx;
  reg  [6:0]  stq_29_bits_uop_pdst;
  reg         stq_29_bits_uop_exception;
  reg  [4:0]  stq_29_bits_uop_mem_cmd;
  reg  [1:0]  stq_29_bits_uop_mem_size;
  reg         stq_29_bits_uop_mem_signed;
  reg         stq_29_bits_uop_is_fence;
  reg         stq_29_bits_uop_is_amo;
  reg         stq_29_bits_uop_uses_ldq;
  reg         stq_29_bits_uop_uses_stq;
  reg  [1:0]  stq_29_bits_uop_dst_rtype;
  reg         stq_29_bits_addr_valid;
  reg  [39:0] stq_29_bits_addr_bits;
  reg         stq_29_bits_addr_is_virtual;
  reg         stq_29_bits_data_valid;
  reg  [63:0] stq_29_bits_data_bits;
  reg         stq_29_bits_committed;
  reg         stq_29_bits_succeeded;
  reg         stq_30_valid;
  reg  [19:0] stq_30_bits_uop_br_mask;
  reg  [6:0]  stq_30_bits_uop_rob_idx;
  reg  [4:0]  stq_30_bits_uop_ldq_idx;
  reg  [4:0]  stq_30_bits_uop_stq_idx;
  reg  [6:0]  stq_30_bits_uop_pdst;
  reg         stq_30_bits_uop_exception;
  reg  [4:0]  stq_30_bits_uop_mem_cmd;
  reg  [1:0]  stq_30_bits_uop_mem_size;
  reg         stq_30_bits_uop_mem_signed;
  reg         stq_30_bits_uop_is_fence;
  reg         stq_30_bits_uop_is_amo;
  reg         stq_30_bits_uop_uses_ldq;
  reg         stq_30_bits_uop_uses_stq;
  reg  [1:0]  stq_30_bits_uop_dst_rtype;
  reg         stq_30_bits_addr_valid;
  reg  [39:0] stq_30_bits_addr_bits;
  reg         stq_30_bits_addr_is_virtual;
  reg         stq_30_bits_data_valid;
  reg  [63:0] stq_30_bits_data_bits;
  reg         stq_30_bits_committed;
  reg         stq_30_bits_succeeded;
  reg         stq_31_valid;
  reg  [19:0] stq_31_bits_uop_br_mask;
  reg  [6:0]  stq_31_bits_uop_rob_idx;
  reg  [4:0]  stq_31_bits_uop_ldq_idx;
  reg  [4:0]  stq_31_bits_uop_stq_idx;
  reg  [6:0]  stq_31_bits_uop_pdst;
  reg         stq_31_bits_uop_exception;
  reg  [4:0]  stq_31_bits_uop_mem_cmd;
  reg  [1:0]  stq_31_bits_uop_mem_size;
  reg         stq_31_bits_uop_mem_signed;
  reg         stq_31_bits_uop_is_fence;
  reg         stq_31_bits_uop_is_amo;
  reg         stq_31_bits_uop_uses_ldq;
  reg         stq_31_bits_uop_uses_stq;
  reg  [1:0]  stq_31_bits_uop_dst_rtype;
  reg         stq_31_bits_addr_valid;
  reg  [39:0] stq_31_bits_addr_bits;
  reg         stq_31_bits_addr_is_virtual;
  reg         stq_31_bits_data_valid;
  reg  [63:0] stq_31_bits_data_bits;
  reg         stq_31_bits_committed;
  reg         stq_31_bits_succeeded;
  reg  [4:0]  ldq_head;
  reg  [4:0]  ldq_tail;
  reg  [4:0]  stq_head;
  reg  [4:0]  stq_tail;
  reg  [4:0]  stq_commit_head;
  reg  [4:0]  stq_execute_head;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp = stq_0_valid;
      5'b00001:
        casez_tmp = stq_1_valid;
      5'b00010:
        casez_tmp = stq_2_valid;
      5'b00011:
        casez_tmp = stq_3_valid;
      5'b00100:
        casez_tmp = stq_4_valid;
      5'b00101:
        casez_tmp = stq_5_valid;
      5'b00110:
        casez_tmp = stq_6_valid;
      5'b00111:
        casez_tmp = stq_7_valid;
      5'b01000:
        casez_tmp = stq_8_valid;
      5'b01001:
        casez_tmp = stq_9_valid;
      5'b01010:
        casez_tmp = stq_10_valid;
      5'b01011:
        casez_tmp = stq_11_valid;
      5'b01100:
        casez_tmp = stq_12_valid;
      5'b01101:
        casez_tmp = stq_13_valid;
      5'b01110:
        casez_tmp = stq_14_valid;
      5'b01111:
        casez_tmp = stq_15_valid;
      5'b10000:
        casez_tmp = stq_16_valid;
      5'b10001:
        casez_tmp = stq_17_valid;
      5'b10010:
        casez_tmp = stq_18_valid;
      5'b10011:
        casez_tmp = stq_19_valid;
      5'b10100:
        casez_tmp = stq_20_valid;
      5'b10101:
        casez_tmp = stq_21_valid;
      5'b10110:
        casez_tmp = stq_22_valid;
      5'b10111:
        casez_tmp = stq_23_valid;
      5'b11000:
        casez_tmp = stq_24_valid;
      5'b11001:
        casez_tmp = stq_25_valid;
      5'b11010:
        casez_tmp = stq_26_valid;
      5'b11011:
        casez_tmp = stq_27_valid;
      5'b11100:
        casez_tmp = stq_28_valid;
      5'b11101:
        casez_tmp = stq_29_valid;
      5'b11110:
        casez_tmp = stq_30_valid;
      default:
        casez_tmp = stq_31_valid;
    endcase
  end // always @(*)
  reg  [2:0]  hella_state;
  reg  [39:0] hella_req_addr;
  reg  [4:0]  hella_req_cmd;
  reg  [1:0]  hella_req_size;
  reg         hella_req_signed;
  reg         hella_req_phys;
  reg  [63:0] hella_data_data;
  reg  [31:0] hella_paddr;
  reg         hella_xcpt_ma_ld;
  reg         hella_xcpt_ma_st;
  reg         hella_xcpt_pf_ld;
  reg         hella_xcpt_pf_st;
  reg         hella_xcpt_gf_ld;
  reg         hella_xcpt_gf_st;
  reg         hella_xcpt_ae_ld;
  reg         hella_xcpt_ae_st;
  reg  [31:0] live_store_mask;
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_0 = stq_0_valid;
      5'b00001:
        casez_tmp_0 = stq_1_valid;
      5'b00010:
        casez_tmp_0 = stq_2_valid;
      5'b00011:
        casez_tmp_0 = stq_3_valid;
      5'b00100:
        casez_tmp_0 = stq_4_valid;
      5'b00101:
        casez_tmp_0 = stq_5_valid;
      5'b00110:
        casez_tmp_0 = stq_6_valid;
      5'b00111:
        casez_tmp_0 = stq_7_valid;
      5'b01000:
        casez_tmp_0 = stq_8_valid;
      5'b01001:
        casez_tmp_0 = stq_9_valid;
      5'b01010:
        casez_tmp_0 = stq_10_valid;
      5'b01011:
        casez_tmp_0 = stq_11_valid;
      5'b01100:
        casez_tmp_0 = stq_12_valid;
      5'b01101:
        casez_tmp_0 = stq_13_valid;
      5'b01110:
        casez_tmp_0 = stq_14_valid;
      5'b01111:
        casez_tmp_0 = stq_15_valid;
      5'b10000:
        casez_tmp_0 = stq_16_valid;
      5'b10001:
        casez_tmp_0 = stq_17_valid;
      5'b10010:
        casez_tmp_0 = stq_18_valid;
      5'b10011:
        casez_tmp_0 = stq_19_valid;
      5'b10100:
        casez_tmp_0 = stq_20_valid;
      5'b10101:
        casez_tmp_0 = stq_21_valid;
      5'b10110:
        casez_tmp_0 = stq_22_valid;
      5'b10111:
        casez_tmp_0 = stq_23_valid;
      5'b11000:
        casez_tmp_0 = stq_24_valid;
      5'b11001:
        casez_tmp_0 = stq_25_valid;
      5'b11010:
        casez_tmp_0 = stq_26_valid;
      5'b11011:
        casez_tmp_0 = stq_27_valid;
      5'b11100:
        casez_tmp_0 = stq_28_valid;
      5'b11101:
        casez_tmp_0 = stq_29_valid;
      5'b11110:
        casez_tmp_0 = stq_30_valid;
      default:
        casez_tmp_0 = stq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_1 = stq_0_bits_committed;
      5'b00001:
        casez_tmp_1 = stq_1_bits_committed;
      5'b00010:
        casez_tmp_1 = stq_2_bits_committed;
      5'b00011:
        casez_tmp_1 = stq_3_bits_committed;
      5'b00100:
        casez_tmp_1 = stq_4_bits_committed;
      5'b00101:
        casez_tmp_1 = stq_5_bits_committed;
      5'b00110:
        casez_tmp_1 = stq_6_bits_committed;
      5'b00111:
        casez_tmp_1 = stq_7_bits_committed;
      5'b01000:
        casez_tmp_1 = stq_8_bits_committed;
      5'b01001:
        casez_tmp_1 = stq_9_bits_committed;
      5'b01010:
        casez_tmp_1 = stq_10_bits_committed;
      5'b01011:
        casez_tmp_1 = stq_11_bits_committed;
      5'b01100:
        casez_tmp_1 = stq_12_bits_committed;
      5'b01101:
        casez_tmp_1 = stq_13_bits_committed;
      5'b01110:
        casez_tmp_1 = stq_14_bits_committed;
      5'b01111:
        casez_tmp_1 = stq_15_bits_committed;
      5'b10000:
        casez_tmp_1 = stq_16_bits_committed;
      5'b10001:
        casez_tmp_1 = stq_17_bits_committed;
      5'b10010:
        casez_tmp_1 = stq_18_bits_committed;
      5'b10011:
        casez_tmp_1 = stq_19_bits_committed;
      5'b10100:
        casez_tmp_1 = stq_20_bits_committed;
      5'b10101:
        casez_tmp_1 = stq_21_bits_committed;
      5'b10110:
        casez_tmp_1 = stq_22_bits_committed;
      5'b10111:
        casez_tmp_1 = stq_23_bits_committed;
      5'b11000:
        casez_tmp_1 = stq_24_bits_committed;
      5'b11001:
        casez_tmp_1 = stq_25_bits_committed;
      5'b11010:
        casez_tmp_1 = stq_26_bits_committed;
      5'b11011:
        casez_tmp_1 = stq_27_bits_committed;
      5'b11100:
        casez_tmp_1 = stq_28_bits_committed;
      5'b11101:
        casez_tmp_1 = stq_29_bits_committed;
      5'b11110:
        casez_tmp_1 = stq_30_bits_committed;
      default:
        casez_tmp_1 = stq_31_bits_committed;
    endcase
  end // always @(*)
  wire        _GEN = casez_tmp_0 & casez_tmp_1;
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_2 = stq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_2 = stq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_2 = stq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_2 = stq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_2 = stq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_2 = stq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_2 = stq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_2 = stq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_2 = stq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_2 = stq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_2 = stq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_2 = stq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_2 = stq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_2 = stq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_2 = stq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_2 = stq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_2 = stq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_2 = stq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_2 = stq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_2 = stq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_2 = stq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_2 = stq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_2 = stq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_2 = stq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_2 = stq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_2 = stq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_2 = stq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_2 = stq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_2 = stq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_2 = stq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_2 = stq_30_bits_uop_is_fence;
      default:
        casez_tmp_2 = stq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_head)
      5'b00000:
        casez_tmp_3 = stq_0_bits_succeeded;
      5'b00001:
        casez_tmp_3 = stq_1_bits_succeeded;
      5'b00010:
        casez_tmp_3 = stq_2_bits_succeeded;
      5'b00011:
        casez_tmp_3 = stq_3_bits_succeeded;
      5'b00100:
        casez_tmp_3 = stq_4_bits_succeeded;
      5'b00101:
        casez_tmp_3 = stq_5_bits_succeeded;
      5'b00110:
        casez_tmp_3 = stq_6_bits_succeeded;
      5'b00111:
        casez_tmp_3 = stq_7_bits_succeeded;
      5'b01000:
        casez_tmp_3 = stq_8_bits_succeeded;
      5'b01001:
        casez_tmp_3 = stq_9_bits_succeeded;
      5'b01010:
        casez_tmp_3 = stq_10_bits_succeeded;
      5'b01011:
        casez_tmp_3 = stq_11_bits_succeeded;
      5'b01100:
        casez_tmp_3 = stq_12_bits_succeeded;
      5'b01101:
        casez_tmp_3 = stq_13_bits_succeeded;
      5'b01110:
        casez_tmp_3 = stq_14_bits_succeeded;
      5'b01111:
        casez_tmp_3 = stq_15_bits_succeeded;
      5'b10000:
        casez_tmp_3 = stq_16_bits_succeeded;
      5'b10001:
        casez_tmp_3 = stq_17_bits_succeeded;
      5'b10010:
        casez_tmp_3 = stq_18_bits_succeeded;
      5'b10011:
        casez_tmp_3 = stq_19_bits_succeeded;
      5'b10100:
        casez_tmp_3 = stq_20_bits_succeeded;
      5'b10101:
        casez_tmp_3 = stq_21_bits_succeeded;
      5'b10110:
        casez_tmp_3 = stq_22_bits_succeeded;
      5'b10111:
        casez_tmp_3 = stq_23_bits_succeeded;
      5'b11000:
        casez_tmp_3 = stq_24_bits_succeeded;
      5'b11001:
        casez_tmp_3 = stq_25_bits_succeeded;
      5'b11010:
        casez_tmp_3 = stq_26_bits_succeeded;
      5'b11011:
        casez_tmp_3 = stq_27_bits_succeeded;
      5'b11100:
        casez_tmp_3 = stq_28_bits_succeeded;
      5'b11101:
        casez_tmp_3 = stq_29_bits_succeeded;
      5'b11110:
        casez_tmp_3 = stq_30_bits_succeeded;
      default:
        casez_tmp_3 = stq_31_bits_succeeded;
    endcase
  end // always @(*)
  wire [4:0]  _GEN_0 = ldq_tail + 5'h1;
  wire [4:0]  _GEN_1 = stq_tail + 5'h1;
  wire        dis_ld_val = io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_ldq & ~io_core_dis_uops_0_bits_exception;
  wire        dis_st_val = io_core_dis_uops_0_valid & io_core_dis_uops_0_bits_uses_stq & ~io_core_dis_uops_0_bits_exception;
  wire        _GEN_2 = dis_st_val & stq_tail == 5'h0;
  wire        _GEN_3 = dis_st_val & stq_tail == 5'h1;
  wire        _GEN_4 = dis_st_val & stq_tail == 5'h2;
  wire        _GEN_5 = dis_st_val & stq_tail == 5'h3;
  wire        _GEN_6 = dis_st_val & stq_tail == 5'h4;
  wire        _GEN_7 = dis_st_val & stq_tail == 5'h5;
  wire        _GEN_8 = dis_st_val & stq_tail == 5'h6;
  wire        _GEN_9 = dis_st_val & stq_tail == 5'h7;
  wire        _GEN_10 = dis_st_val & stq_tail == 5'h8;
  wire        _GEN_11 = dis_st_val & stq_tail == 5'h9;
  wire        _GEN_12 = dis_st_val & stq_tail == 5'hA;
  wire        _GEN_13 = dis_st_val & stq_tail == 5'hB;
  wire        _GEN_14 = dis_st_val & stq_tail == 5'hC;
  wire        _GEN_15 = dis_st_val & stq_tail == 5'hD;
  wire        _GEN_16 = dis_st_val & stq_tail == 5'hE;
  wire        _GEN_17 = dis_st_val & stq_tail == 5'hF;
  wire        _GEN_18 = dis_st_val & stq_tail == 5'h10;
  wire        _GEN_19 = dis_st_val & stq_tail == 5'h11;
  wire        _GEN_20 = dis_st_val & stq_tail == 5'h12;
  wire        _GEN_21 = dis_st_val & stq_tail == 5'h13;
  wire        _GEN_22 = dis_st_val & stq_tail == 5'h14;
  wire        _GEN_23 = dis_st_val & stq_tail == 5'h15;
  wire        _GEN_24 = dis_st_val & stq_tail == 5'h16;
  wire        _GEN_25 = dis_st_val & stq_tail == 5'h17;
  wire        _GEN_26 = dis_st_val & stq_tail == 5'h18;
  wire        _GEN_27 = dis_st_val & stq_tail == 5'h19;
  wire        _GEN_28 = dis_st_val & stq_tail == 5'h1A;
  wire        _GEN_29 = dis_st_val & stq_tail == 5'h1B;
  wire        _GEN_30 = dis_st_val & stq_tail == 5'h1C;
  wire        _GEN_31 = dis_st_val & stq_tail == 5'h1D;
  wire        _GEN_32 = dis_st_val & stq_tail == 5'h1E;
  wire        _GEN_33 = dis_st_val & (&stq_tail);
  wire        _GEN_34 = dis_ld_val & ldq_tail == 5'h0;
  wire        _GEN_35 = dis_ld_val & ldq_tail == 5'h1;
  wire        _GEN_36 = dis_ld_val & ldq_tail == 5'h2;
  wire        _GEN_37 = dis_ld_val & ldq_tail == 5'h3;
  wire        _GEN_38 = dis_ld_val & ldq_tail == 5'h4;
  wire        _GEN_39 = dis_ld_val & ldq_tail == 5'h5;
  wire        _GEN_40 = dis_ld_val & ldq_tail == 5'h6;
  wire        _GEN_41 = dis_ld_val & ldq_tail == 5'h7;
  wire        _GEN_42 = dis_ld_val & ldq_tail == 5'h8;
  wire        _GEN_43 = dis_ld_val & ldq_tail == 5'h9;
  wire        _GEN_44 = dis_ld_val & ldq_tail == 5'hA;
  wire        _GEN_45 = dis_ld_val & ldq_tail == 5'hB;
  wire        _GEN_46 = dis_ld_val & ldq_tail == 5'hC;
  wire        _GEN_47 = dis_ld_val & ldq_tail == 5'hD;
  wire        _GEN_48 = dis_ld_val & ldq_tail == 5'hE;
  wire        _GEN_49 = dis_ld_val & ldq_tail == 5'hF;
  wire        _GEN_50 = dis_ld_val & ldq_tail == 5'h10;
  wire        _GEN_51 = dis_ld_val & ldq_tail == 5'h11;
  wire        _GEN_52 = dis_ld_val & ldq_tail == 5'h12;
  wire        _GEN_53 = dis_ld_val & ldq_tail == 5'h13;
  wire        _GEN_54 = dis_ld_val & ldq_tail == 5'h14;
  wire        _GEN_55 = dis_ld_val & ldq_tail == 5'h15;
  wire        _GEN_56 = dis_ld_val & ldq_tail == 5'h16;
  wire        _GEN_57 = dis_ld_val & ldq_tail == 5'h17;
  wire        _GEN_58 = dis_ld_val & ldq_tail == 5'h18;
  wire        _GEN_59 = dis_ld_val & ldq_tail == 5'h19;
  wire        _GEN_60 = dis_ld_val & ldq_tail == 5'h1A;
  wire        _GEN_61 = dis_ld_val & ldq_tail == 5'h1B;
  wire        _GEN_62 = dis_ld_val & ldq_tail == 5'h1C;
  wire        _GEN_63 = dis_ld_val & ldq_tail == 5'h1D;
  wire        _GEN_64 = dis_ld_val & ldq_tail == 5'h1E;
  wire        _GEN_65 = dis_ld_val & (&ldq_tail);
  wire [4:0]  _GEN_66 = dis_ld_val ? _GEN_0 : ldq_tail;
  wire [4:0]  _ldq_T_35_bits_youngest_stq_idx = dis_st_val ? _GEN_1 : stq_tail;
  wire [4:0]  _GEN_67 = _GEN_66 + 5'h1;
  wire [4:0]  _GEN_68 = _ldq_T_35_bits_youngest_stq_idx + 5'h1;
  wire        dis_ld_val_1 = io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_ldq & ~io_core_dis_uops_1_bits_exception;
  wire        dis_st_val_1 = io_core_dis_uops_1_valid & io_core_dis_uops_1_bits_uses_stq & ~io_core_dis_uops_1_bits_exception;
  wire        _GEN_69 = _GEN_66 == 5'h0;
  wire        _GEN_70 = _GEN_66 == 5'h1;
  wire        _GEN_71 = _GEN_66 == 5'h2;
  wire        _GEN_72 = _GEN_66 == 5'h3;
  wire        _GEN_73 = _GEN_66 == 5'h4;
  wire        _GEN_74 = _GEN_66 == 5'h5;
  wire        _GEN_75 = _GEN_66 == 5'h6;
  wire        _GEN_76 = _GEN_66 == 5'h7;
  wire        _GEN_77 = _GEN_66 == 5'h8;
  wire        _GEN_78 = _GEN_66 == 5'h9;
  wire        _GEN_79 = _GEN_66 == 5'hA;
  wire        _GEN_80 = _GEN_66 == 5'hB;
  wire        _GEN_81 = _GEN_66 == 5'hC;
  wire        _GEN_82 = _GEN_66 == 5'hD;
  wire        _GEN_83 = _GEN_66 == 5'hE;
  wire        _GEN_84 = _GEN_66 == 5'hF;
  wire        _GEN_85 = _GEN_66 == 5'h10;
  wire        _GEN_86 = _GEN_66 == 5'h11;
  wire        _GEN_87 = _GEN_66 == 5'h12;
  wire        _GEN_88 = _GEN_66 == 5'h13;
  wire        _GEN_89 = _GEN_66 == 5'h14;
  wire        _GEN_90 = _GEN_66 == 5'h15;
  wire        _GEN_91 = _GEN_66 == 5'h16;
  wire        _GEN_92 = _GEN_66 == 5'h17;
  wire        _GEN_93 = _GEN_66 == 5'h18;
  wire        _GEN_94 = _GEN_66 == 5'h19;
  wire        _GEN_95 = _GEN_66 == 5'h1A;
  wire        _GEN_96 = _GEN_66 == 5'h1B;
  wire        _GEN_97 = _GEN_66 == 5'h1C;
  wire        _GEN_98 = _GEN_66 == 5'h1D;
  wire        _GEN_99 = _GEN_66 == 5'h1E;
  wire        _GEN_100 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h0;
  wire        _GEN_101 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h1;
  wire        _GEN_102 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h2;
  wire        _GEN_103 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h3;
  wire        _GEN_104 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h4;
  wire        _GEN_105 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h5;
  wire        _GEN_106 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h6;
  wire        _GEN_107 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h7;
  wire        _GEN_108 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h8;
  wire        _GEN_109 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h9;
  wire        _GEN_110 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'hA;
  wire        _GEN_111 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'hB;
  wire        _GEN_112 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'hC;
  wire        _GEN_113 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'hD;
  wire        _GEN_114 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'hE;
  wire        _GEN_115 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'hF;
  wire        _GEN_116 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h10;
  wire        _GEN_117 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h11;
  wire        _GEN_118 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h12;
  wire        _GEN_119 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h13;
  wire        _GEN_120 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h14;
  wire        _GEN_121 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h15;
  wire        _GEN_122 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h16;
  wire        _GEN_123 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h17;
  wire        _GEN_124 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h18;
  wire        _GEN_125 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h19;
  wire        _GEN_126 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h1A;
  wire        _GEN_127 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h1B;
  wire        _GEN_128 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h1C;
  wire        _GEN_129 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h1D;
  wire        _GEN_130 = dis_st_val_1 & _ldq_T_35_bits_youngest_stq_idx == 5'h1E;
  wire        _GEN_131 = dis_st_val_1 & (&_ldq_T_35_bits_youngest_stq_idx);
  wire        _GEN_132 = dis_ld_val_1 & _GEN_69;
  wire        _GEN_133 = dis_ld_val_1 & _GEN_70;
  wire        _GEN_134 = dis_ld_val_1 & _GEN_71;
  wire        _GEN_135 = dis_ld_val_1 & _GEN_72;
  wire        _GEN_136 = dis_ld_val_1 & _GEN_73;
  wire        _GEN_137 = dis_ld_val_1 & _GEN_74;
  wire        _GEN_138 = dis_ld_val_1 & _GEN_75;
  wire        _GEN_139 = dis_ld_val_1 & _GEN_76;
  wire        _GEN_140 = dis_ld_val_1 & _GEN_77;
  wire        _GEN_141 = dis_ld_val_1 & _GEN_78;
  wire        _GEN_142 = dis_ld_val_1 & _GEN_79;
  wire        _GEN_143 = dis_ld_val_1 & _GEN_80;
  wire        _GEN_144 = dis_ld_val_1 & _GEN_81;
  wire        _GEN_145 = dis_ld_val_1 & _GEN_82;
  wire        _GEN_146 = dis_ld_val_1 & _GEN_83;
  wire        _GEN_147 = dis_ld_val_1 & _GEN_84;
  wire        _GEN_148 = dis_ld_val_1 & _GEN_85;
  wire        _GEN_149 = dis_ld_val_1 & _GEN_86;
  wire        _GEN_150 = dis_ld_val_1 & _GEN_87;
  wire        _GEN_151 = dis_ld_val_1 & _GEN_88;
  wire        _GEN_152 = dis_ld_val_1 & _GEN_89;
  wire        _GEN_153 = dis_ld_val_1 & _GEN_90;
  wire        _GEN_154 = dis_ld_val_1 & _GEN_91;
  wire        _GEN_155 = dis_ld_val_1 & _GEN_92;
  wire        _GEN_156 = dis_ld_val_1 & _GEN_93;
  wire        _GEN_157 = dis_ld_val_1 & _GEN_94;
  wire        _GEN_158 = dis_ld_val_1 & _GEN_95;
  wire        _GEN_159 = dis_ld_val_1 & _GEN_96;
  wire        _GEN_160 = dis_ld_val_1 & _GEN_97;
  wire        _GEN_161 = dis_ld_val_1 & _GEN_98;
  wire        _GEN_162 = dis_ld_val_1 & _GEN_99;
  wire        _GEN_163 = dis_ld_val_1 & (&_GEN_66);
  wire [4:0]  _GEN_164 = dis_ld_val_1 ? _GEN_67 : _GEN_66;
  wire [4:0]  _ldq_T_75_bits_youngest_stq_idx = dis_st_val_1 ? _GEN_68 : _ldq_T_35_bits_youngest_stq_idx;
  wire [4:0]  _GEN_165 = _GEN_164 + 5'h1;
  wire [4:0]  _GEN_166 = _ldq_T_75_bits_youngest_stq_idx + 5'h1;
  wire        dis_ld_val_2 = io_core_dis_uops_2_valid & io_core_dis_uops_2_bits_uses_ldq & ~io_core_dis_uops_2_bits_exception;
  wire        dis_st_val_2 = io_core_dis_uops_2_valid & io_core_dis_uops_2_bits_uses_stq & ~io_core_dis_uops_2_bits_exception;
  wire        _GEN_167 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h0;
  wire        _GEN_168 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h1;
  wire        _GEN_169 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h2;
  wire        _GEN_170 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h3;
  wire        _GEN_171 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h4;
  wire        _GEN_172 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h5;
  wire        _GEN_173 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h6;
  wire        _GEN_174 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h7;
  wire        _GEN_175 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h8;
  wire        _GEN_176 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h9;
  wire        _GEN_177 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'hA;
  wire        _GEN_178 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'hB;
  wire        _GEN_179 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'hC;
  wire        _GEN_180 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'hD;
  wire        _GEN_181 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'hE;
  wire        _GEN_182 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'hF;
  wire        _GEN_183 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h10;
  wire        _GEN_184 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h11;
  wire        _GEN_185 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h12;
  wire        _GEN_186 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h13;
  wire        _GEN_187 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h14;
  wire        _GEN_188 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h15;
  wire        _GEN_189 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h16;
  wire        _GEN_190 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h17;
  wire        _GEN_191 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h18;
  wire        _GEN_192 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h19;
  wire        _GEN_193 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h1A;
  wire        _GEN_194 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h1B;
  wire        _GEN_195 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h1C;
  wire        _GEN_196 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h1D;
  wire        _GEN_197 = dis_st_val_2 & _ldq_T_75_bits_youngest_stq_idx == 5'h1E;
  wire        _GEN_198 = dis_st_val_2 & (&_ldq_T_75_bits_youngest_stq_idx);
  wire        _GEN_199 = dis_ld_val_2 & _GEN_164 == 5'h0;
  wire        _GEN_200 = dis_ld_val_2 & _GEN_164 == 5'h1;
  wire        _GEN_201 = dis_ld_val_2 & _GEN_164 == 5'h2;
  wire        _GEN_202 = dis_ld_val_2 & _GEN_164 == 5'h3;
  wire        _GEN_203 = dis_ld_val_2 & _GEN_164 == 5'h4;
  wire        _GEN_204 = dis_ld_val_2 & _GEN_164 == 5'h5;
  wire        _GEN_205 = dis_ld_val_2 & _GEN_164 == 5'h6;
  wire        _GEN_206 = dis_ld_val_2 & _GEN_164 == 5'h7;
  wire        _GEN_207 = dis_ld_val_2 & _GEN_164 == 5'h8;
  wire        _GEN_208 = dis_ld_val_2 & _GEN_164 == 5'h9;
  wire        _GEN_209 = dis_ld_val_2 & _GEN_164 == 5'hA;
  wire        _GEN_210 = dis_ld_val_2 & _GEN_164 == 5'hB;
  wire        _GEN_211 = dis_ld_val_2 & _GEN_164 == 5'hC;
  wire        _GEN_212 = dis_ld_val_2 & _GEN_164 == 5'hD;
  wire        _GEN_213 = dis_ld_val_2 & _GEN_164 == 5'hE;
  wire        _GEN_214 = dis_ld_val_2 & _GEN_164 == 5'hF;
  wire        _GEN_215 = dis_ld_val_2 & _GEN_164 == 5'h10;
  wire        _GEN_216 = dis_ld_val_2 & _GEN_164 == 5'h11;
  wire        _GEN_217 = dis_ld_val_2 & _GEN_164 == 5'h12;
  wire        _GEN_218 = dis_ld_val_2 & _GEN_164 == 5'h13;
  wire        _GEN_219 = dis_ld_val_2 & _GEN_164 == 5'h14;
  wire        _GEN_220 = dis_ld_val_2 & _GEN_164 == 5'h15;
  wire        _GEN_221 = dis_ld_val_2 & _GEN_164 == 5'h16;
  wire        _GEN_222 = dis_ld_val_2 & _GEN_164 == 5'h17;
  wire        _GEN_223 = dis_ld_val_2 & _GEN_164 == 5'h18;
  wire        _GEN_224 = dis_ld_val_2 & _GEN_164 == 5'h19;
  wire        _GEN_225 = dis_ld_val_2 & _GEN_164 == 5'h1A;
  wire        _GEN_226 = dis_ld_val_2 & _GEN_164 == 5'h1B;
  wire        _GEN_227 = dis_ld_val_2 & _GEN_164 == 5'h1C;
  wire        _GEN_228 = dis_ld_val_2 & _GEN_164 == 5'h1D;
  wire        _GEN_229 = dis_ld_val_2 & _GEN_164 == 5'h1E;
  wire        _GEN_230 = dis_ld_val_2 & (&_GEN_164);
  wire [4:0]  _GEN_231 = dis_ld_val_2 ? _GEN_165 : _GEN_164;
  wire [4:0]  _ldq_T_115_bits_youngest_stq_idx = dis_st_val_2 ? _GEN_166 : _ldq_T_75_bits_youngest_stq_idx;
  wire [4:0]  _GEN_232 = _GEN_231 + 5'h1;
  wire [4:0]  _GEN_233 = _ldq_T_115_bits_youngest_stq_idx + 5'h1;
  wire        dis_ld_val_3 = io_core_dis_uops_3_valid & io_core_dis_uops_3_bits_uses_ldq & ~io_core_dis_uops_3_bits_exception;
  wire        dis_st_val_3 = io_core_dis_uops_3_valid & io_core_dis_uops_3_bits_uses_stq & ~io_core_dis_uops_3_bits_exception;
  wire        _GEN_234 = _GEN_231 == 5'h0;
  wire        _GEN_235 = _GEN_231 == 5'h1;
  wire        _GEN_236 = _GEN_231 == 5'h2;
  wire        _GEN_237 = _GEN_231 == 5'h3;
  wire        _GEN_238 = _GEN_231 == 5'h4;
  wire        _GEN_239 = _GEN_231 == 5'h5;
  wire        _GEN_240 = _GEN_231 == 5'h6;
  wire        _GEN_241 = _GEN_231 == 5'h7;
  wire        _GEN_242 = _GEN_231 == 5'h8;
  wire        _GEN_243 = _GEN_231 == 5'h9;
  wire        _GEN_244 = _GEN_231 == 5'hA;
  wire        _GEN_245 = _GEN_231 == 5'hB;
  wire        _GEN_246 = _GEN_231 == 5'hC;
  wire        _GEN_247 = _GEN_231 == 5'hD;
  wire        _GEN_248 = _GEN_231 == 5'hE;
  wire        _GEN_249 = _GEN_231 == 5'hF;
  wire        _GEN_250 = _GEN_231 == 5'h10;
  wire        _GEN_251 = _GEN_231 == 5'h11;
  wire        _GEN_252 = _GEN_231 == 5'h12;
  wire        _GEN_253 = _GEN_231 == 5'h13;
  wire        _GEN_254 = _GEN_231 == 5'h14;
  wire        _GEN_255 = _GEN_231 == 5'h15;
  wire        _GEN_256 = _GEN_231 == 5'h16;
  wire        _GEN_257 = _GEN_231 == 5'h17;
  wire        _GEN_258 = _GEN_231 == 5'h18;
  wire        _GEN_259 = _GEN_231 == 5'h19;
  wire        _GEN_260 = _GEN_231 == 5'h1A;
  wire        _GEN_261 = _GEN_231 == 5'h1B;
  wire        _GEN_262 = _GEN_231 == 5'h1C;
  wire        _GEN_263 = _GEN_231 == 5'h1D;
  wire        _GEN_264 = _GEN_231 == 5'h1E;
  wire        _GEN_265 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h0;
  wire        _GEN_266 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h1;
  wire        _GEN_267 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h2;
  wire        _GEN_268 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h3;
  wire        _GEN_269 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h4;
  wire        _GEN_270 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h5;
  wire        _GEN_271 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h6;
  wire        _GEN_272 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h7;
  wire        _GEN_273 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h8;
  wire        _GEN_274 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h9;
  wire        _GEN_275 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'hA;
  wire        _GEN_276 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'hB;
  wire        _GEN_277 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'hC;
  wire        _GEN_278 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'hD;
  wire        _GEN_279 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'hE;
  wire        _GEN_280 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'hF;
  wire        _GEN_281 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h10;
  wire        _GEN_282 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h11;
  wire        _GEN_283 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h12;
  wire        _GEN_284 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h13;
  wire        _GEN_285 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h14;
  wire        _GEN_286 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h15;
  wire        _GEN_287 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h16;
  wire        _GEN_288 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h17;
  wire        _GEN_289 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h18;
  wire        _GEN_290 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h19;
  wire        _GEN_291 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h1A;
  wire        _GEN_292 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h1B;
  wire        _GEN_293 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h1C;
  wire        _GEN_294 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h1D;
  wire        _GEN_295 = dis_st_val_3 & _ldq_T_115_bits_youngest_stq_idx == 5'h1E;
  wire        _GEN_296 = dis_st_val_3 & (&_ldq_T_115_bits_youngest_stq_idx);
  wire        _GEN_297 = dis_ld_val_3 & _GEN_234;
  wire        _GEN_298 = dis_ld_val_3 & _GEN_235;
  wire        _GEN_299 = dis_ld_val_3 & _GEN_236;
  wire        _GEN_300 = dis_ld_val_3 & _GEN_237;
  wire        _GEN_301 = dis_ld_val_3 & _GEN_238;
  wire        _GEN_302 = dis_ld_val_3 & _GEN_239;
  wire        _GEN_303 = dis_ld_val_3 & _GEN_240;
  wire        _GEN_304 = dis_ld_val_3 & _GEN_241;
  wire        _GEN_305 = dis_ld_val_3 & _GEN_242;
  wire        _GEN_306 = dis_ld_val_3 & _GEN_243;
  wire        _GEN_307 = dis_ld_val_3 & _GEN_244;
  wire        _GEN_308 = dis_ld_val_3 & _GEN_245;
  wire        _GEN_309 = dis_ld_val_3 & _GEN_246;
  wire        _GEN_310 = dis_ld_val_3 & _GEN_247;
  wire        _GEN_311 = dis_ld_val_3 & _GEN_248;
  wire        _GEN_312 = dis_ld_val_3 & _GEN_249;
  wire        _GEN_313 = dis_ld_val_3 & _GEN_250;
  wire        _GEN_314 = dis_ld_val_3 & _GEN_251;
  wire        _GEN_315 = dis_ld_val_3 & _GEN_252;
  wire        _GEN_316 = dis_ld_val_3 & _GEN_253;
  wire        _GEN_317 = dis_ld_val_3 & _GEN_254;
  wire        _GEN_318 = dis_ld_val_3 & _GEN_255;
  wire        _GEN_319 = dis_ld_val_3 & _GEN_256;
  wire        _GEN_320 = dis_ld_val_3 & _GEN_257;
  wire        _GEN_321 = dis_ld_val_3 & _GEN_258;
  wire        _GEN_322 = dis_ld_val_3 & _GEN_259;
  wire        _GEN_323 = dis_ld_val_3 & _GEN_260;
  wire        _GEN_324 = dis_ld_val_3 & _GEN_261;
  wire        _GEN_325 = dis_ld_val_3 & _GEN_262;
  wire        _GEN_326 = dis_ld_val_3 & _GEN_263;
  wire        _GEN_327 = dis_ld_val_3 & _GEN_264;
  wire        _GEN_328 = dis_ld_val_3 & (&_GEN_231);
  wire [38:0] exe_req_0_bits_sfence_bits_addr = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_bits_addr : io_core_exe_0_req_bits_sfence_bits_addr;
  wire        exe_req_0_bits_sfence_valid = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_valid : io_core_exe_0_req_bits_sfence_valid;
  wire        exe_req_0_bits_mxcpt_valid = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_mxcpt_valid : io_core_exe_0_req_bits_mxcpt_valid;
  wire [1:0]  mem_incoming_uop_out_mem_size = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_mem_size : io_core_exe_0_req_bits_uop_mem_size;
  wire [4:0]  mem_incoming_uop_out_mem_cmd = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_mem_cmd : io_core_exe_0_req_bits_uop_mem_cmd;
  wire [4:0]  stq_incoming_idx_0 = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_stq_idx : io_core_exe_0_req_bits_uop_stq_idx;
  wire [4:0]  ldq_incoming_idx_0 = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ldq_idx : io_core_exe_0_req_bits_uop_ldq_idx;
  wire [19:0] exe_req_0_bits_uop_br_mask = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_br_mask : io_core_exe_0_req_bits_uop_br_mask;
  wire        mem_incoming_uop_out_ctrl_is_std = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_is_std : io_core_exe_0_req_bits_uop_ctrl_is_std;
  wire        mem_incoming_uop_out_ctrl_is_sta = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_is_sta : io_core_exe_0_req_bits_uop_ctrl_is_sta;
  wire        mem_incoming_uop_out_ctrl_is_load = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_ctrl_is_load : io_core_exe_0_req_bits_uop_ctrl_is_load;
  wire        exe_req_0_valid = io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_valid : io_core_exe_0_req_valid;
  wire        _GEN_329 = io_core_exe_1_req_bits_sfence_valid | ~io_core_exe_0_req_bits_sfence_valid;
  wire [38:0] exe_req_1_bits_sfence_bits_addr = _GEN_329 ? io_core_exe_1_req_bits_sfence_bits_addr : io_core_exe_0_req_bits_sfence_bits_addr;
  wire        exe_req_1_bits_sfence_valid = _GEN_329 ? io_core_exe_1_req_bits_sfence_valid : io_core_exe_0_req_bits_sfence_valid;
  wire        exe_req_1_bits_mxcpt_valid = _GEN_329 ? io_core_exe_1_req_bits_mxcpt_valid : io_core_exe_0_req_bits_mxcpt_valid;
  wire        exe_req_1_bits_uop_uses_stq = _GEN_329 ? io_core_exe_1_req_bits_uop_uses_stq : io_core_exe_0_req_bits_uop_uses_stq;
  wire        exe_req_1_bits_uop_uses_ldq = _GEN_329 ? io_core_exe_1_req_bits_uop_uses_ldq : io_core_exe_0_req_bits_uop_uses_ldq;
  wire        exe_req_1_bits_uop_is_amo = _GEN_329 ? io_core_exe_1_req_bits_uop_is_amo : io_core_exe_0_req_bits_uop_is_amo;
  wire        exe_req_1_bits_uop_mem_signed = _GEN_329 ? io_core_exe_1_req_bits_uop_mem_signed : io_core_exe_0_req_bits_uop_mem_signed;
  wire [1:0]  exe_req_1_bits_uop_mem_size = _GEN_329 ? io_core_exe_1_req_bits_uop_mem_size : io_core_exe_0_req_bits_uop_mem_size;
  wire [4:0]  exe_req_1_bits_uop_mem_cmd = _GEN_329 ? io_core_exe_1_req_bits_uop_mem_cmd : io_core_exe_0_req_bits_uop_mem_cmd;
  wire [4:0]  stq_incoming_idx_1 = _GEN_329 ? io_core_exe_1_req_bits_uop_stq_idx : io_core_exe_0_req_bits_uop_stq_idx;
  wire [4:0]  ldq_incoming_idx_1 = _GEN_329 ? io_core_exe_1_req_bits_uop_ldq_idx : io_core_exe_0_req_bits_uop_ldq_idx;
  wire [19:0] exe_req_1_bits_uop_br_mask = _GEN_329 ? io_core_exe_1_req_bits_uop_br_mask : io_core_exe_0_req_bits_uop_br_mask;
  wire        exe_req_1_bits_uop_ctrl_is_std = _GEN_329 ? io_core_exe_1_req_bits_uop_ctrl_is_std : io_core_exe_0_req_bits_uop_ctrl_is_std;
  wire        exe_req_1_bits_uop_ctrl_is_sta = _GEN_329 ? io_core_exe_1_req_bits_uop_ctrl_is_sta : io_core_exe_0_req_bits_uop_ctrl_is_sta;
  wire        exe_req_1_bits_uop_ctrl_is_load = _GEN_329 ? io_core_exe_1_req_bits_uop_ctrl_is_load : io_core_exe_0_req_bits_uop_ctrl_is_load;
  wire        exe_req_1_valid = _GEN_329 ? io_core_exe_1_req_valid : io_core_exe_0_req_valid;
  reg         p1_block_load_mask_0;
  reg         p1_block_load_mask_1;
  reg         p1_block_load_mask_2;
  reg         p1_block_load_mask_3;
  reg         p1_block_load_mask_4;
  reg         p1_block_load_mask_5;
  reg         p1_block_load_mask_6;
  reg         p1_block_load_mask_7;
  reg         p1_block_load_mask_8;
  reg         p1_block_load_mask_9;
  reg         p1_block_load_mask_10;
  reg         p1_block_load_mask_11;
  reg         p1_block_load_mask_12;
  reg         p1_block_load_mask_13;
  reg         p1_block_load_mask_14;
  reg         p1_block_load_mask_15;
  reg         p1_block_load_mask_16;
  reg         p1_block_load_mask_17;
  reg         p1_block_load_mask_18;
  reg         p1_block_load_mask_19;
  reg         p1_block_load_mask_20;
  reg         p1_block_load_mask_21;
  reg         p1_block_load_mask_22;
  reg         p1_block_load_mask_23;
  reg         p1_block_load_mask_24;
  reg         p1_block_load_mask_25;
  reg         p1_block_load_mask_26;
  reg         p1_block_load_mask_27;
  reg         p1_block_load_mask_28;
  reg         p1_block_load_mask_29;
  reg         p1_block_load_mask_30;
  reg         p1_block_load_mask_31;
  reg         p2_block_load_mask_0;
  reg         p2_block_load_mask_1;
  reg         p2_block_load_mask_2;
  reg         p2_block_load_mask_3;
  reg         p2_block_load_mask_4;
  reg         p2_block_load_mask_5;
  reg         p2_block_load_mask_6;
  reg         p2_block_load_mask_7;
  reg         p2_block_load_mask_8;
  reg         p2_block_load_mask_9;
  reg         p2_block_load_mask_10;
  reg         p2_block_load_mask_11;
  reg         p2_block_load_mask_12;
  reg         p2_block_load_mask_13;
  reg         p2_block_load_mask_14;
  reg         p2_block_load_mask_15;
  reg         p2_block_load_mask_16;
  reg         p2_block_load_mask_17;
  reg         p2_block_load_mask_18;
  reg         p2_block_load_mask_19;
  reg         p2_block_load_mask_20;
  reg         p2_block_load_mask_21;
  reg         p2_block_load_mask_22;
  reg         p2_block_load_mask_23;
  reg         p2_block_load_mask_24;
  reg         p2_block_load_mask_25;
  reg         p2_block_load_mask_26;
  reg         p2_block_load_mask_27;
  reg         p2_block_load_mask_28;
  reg         p2_block_load_mask_29;
  reg         p2_block_load_mask_30;
  reg         p2_block_load_mask_31;
  always @(*) begin
    casez (ldq_incoming_idx_0)
      5'b00000:
        casez_tmp_4 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_4 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_4 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_4 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_4 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_4 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_4 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_4 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_4 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_4 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_4 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_4 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_4 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_4 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_4 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_4 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_4 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_4 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_4 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_4 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_4 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_4 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_4 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_4 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_4 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_4 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_4 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_4 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_4 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_4 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_4 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_4 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_0)
      5'b00000:
        casez_tmp_5 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_5 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_5 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_5 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_5 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_5 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_5 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_5 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_5 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_5 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_5 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_5 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_5 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_5 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_5 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_5 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_5 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_5 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_5 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_5 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_5 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_5 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_5 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_5 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_5 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_5 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_5 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_5 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_5 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_5 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_5 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_5 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_0)
      5'b00000:
        casez_tmp_6 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_6 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_6 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_6 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_6 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_6 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_6 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_6 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_6 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_6 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_6 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_6 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_6 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_6 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_6 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_6 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_6 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_6 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_6 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_6 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_6 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_6 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_6 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_6 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_6 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_6 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_6 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_6 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_6 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_6 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_6 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_6 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_0)
      5'b00000:
        casez_tmp_7 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_7 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_7 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_7 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_7 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_7 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_7 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_7 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_7 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_7 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_7 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_7 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_7 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_7 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_7 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_7 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_7 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_7 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_7 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_7 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_7 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_7 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_7 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_7 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_7 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_7 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_7 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_7 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_7 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_7 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_7 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_7 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_1)
      5'b00000:
        casez_tmp_8 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_8 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_8 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_8 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_8 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_8 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_8 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_8 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_8 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_8 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_8 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_8 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_8 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_8 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_8 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_8 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_8 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_8 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_8 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_8 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_8 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_8 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_8 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_8 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_8 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_8 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_8 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_8 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_8 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_8 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_8 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_8 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_1)
      5'b00000:
        casez_tmp_9 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_9 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_9 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_9 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_9 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_9 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_9 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_9 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_9 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_9 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_9 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_9 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_9 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_9 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_9 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_9 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_9 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_9 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_9 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_9 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_9 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_9 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_9 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_9 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_9 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_9 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_9 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_9 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_9 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_9 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_9 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_9 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_1)
      5'b00000:
        casez_tmp_10 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_10 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_10 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_10 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_10 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_10 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_10 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_10 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_10 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_10 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_10 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_10 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_10 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_10 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_10 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_10 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_10 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_10 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_10 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_10 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_10 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_10 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_10 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_10 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_10 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_10 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_10 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_10 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_10 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_10 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_10 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_10 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_incoming_idx_1)
      5'b00000:
        casez_tmp_11 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_11 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_11 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_11 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_11 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_11 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_11 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_11 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_11 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_11 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_11 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_11 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_11 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_11 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_11 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_11 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_11 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_11 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_11 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_11 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_11 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_11 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_11 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_11 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_11 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_11 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_11 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_11 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_11 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_11 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_11 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_11 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_12 = stq_0_valid;
      5'b00001:
        casez_tmp_12 = stq_1_valid;
      5'b00010:
        casez_tmp_12 = stq_2_valid;
      5'b00011:
        casez_tmp_12 = stq_3_valid;
      5'b00100:
        casez_tmp_12 = stq_4_valid;
      5'b00101:
        casez_tmp_12 = stq_5_valid;
      5'b00110:
        casez_tmp_12 = stq_6_valid;
      5'b00111:
        casez_tmp_12 = stq_7_valid;
      5'b01000:
        casez_tmp_12 = stq_8_valid;
      5'b01001:
        casez_tmp_12 = stq_9_valid;
      5'b01010:
        casez_tmp_12 = stq_10_valid;
      5'b01011:
        casez_tmp_12 = stq_11_valid;
      5'b01100:
        casez_tmp_12 = stq_12_valid;
      5'b01101:
        casez_tmp_12 = stq_13_valid;
      5'b01110:
        casez_tmp_12 = stq_14_valid;
      5'b01111:
        casez_tmp_12 = stq_15_valid;
      5'b10000:
        casez_tmp_12 = stq_16_valid;
      5'b10001:
        casez_tmp_12 = stq_17_valid;
      5'b10010:
        casez_tmp_12 = stq_18_valid;
      5'b10011:
        casez_tmp_12 = stq_19_valid;
      5'b10100:
        casez_tmp_12 = stq_20_valid;
      5'b10101:
        casez_tmp_12 = stq_21_valid;
      5'b10110:
        casez_tmp_12 = stq_22_valid;
      5'b10111:
        casez_tmp_12 = stq_23_valid;
      5'b11000:
        casez_tmp_12 = stq_24_valid;
      5'b11001:
        casez_tmp_12 = stq_25_valid;
      5'b11010:
        casez_tmp_12 = stq_26_valid;
      5'b11011:
        casez_tmp_12 = stq_27_valid;
      5'b11100:
        casez_tmp_12 = stq_28_valid;
      5'b11101:
        casez_tmp_12 = stq_29_valid;
      5'b11110:
        casez_tmp_12 = stq_30_valid;
      default:
        casez_tmp_12 = stq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_13 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_13 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_13 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_13 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_13 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_13 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_13 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_13 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_13 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_13 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_13 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_13 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_13 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_13 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_13 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_13 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_13 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_13 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_13 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_13 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_13 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_13 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_13 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_13 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_13 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_13 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_13 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_13 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_13 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_13 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_13 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_13 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_14 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_14 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_14 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_14 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_14 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_14 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_14 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_14 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_14 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_14 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_14 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_14 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_14 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_14 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_14 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_14 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_14 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_14 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_14 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_14 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_14 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_14 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_14 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_14 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_14 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_14 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_14 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_14 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_14 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_14 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_14 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_14 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_15 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_15 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_15 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_15 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_15 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_15 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_15 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_15 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_15 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_15 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_15 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_15 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_15 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_15 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_15 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_15 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_15 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_15 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_15 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_15 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_15 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_15 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_15 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_15 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_15 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_15 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_15 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_15 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_15 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_15 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_15 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_15 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_16 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_16 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_16 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_16 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_16 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_16 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_16 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_16 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_16 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_16 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_16 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_16 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_16 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_16 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_16 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_16 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_16 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_16 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_16 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_16 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_16 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_16 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_16 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_16 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_16 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_16 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_16 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_16 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_16 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_16 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_16 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_16 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_17 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_17 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_17 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_17 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_17 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_17 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_17 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_17 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_17 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_17 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_17 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_17 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_17 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_17 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_17 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_17 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_17 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_17 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_17 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_17 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_17 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_17 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_17 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_17 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_17 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_17 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_17 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_17 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_17 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_17 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_17 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_17 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_18 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_18 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_18 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_18 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_18 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_18 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_18 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_18 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_18 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_18 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_18 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_18 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_18 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_18 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_18 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_18 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_18 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_18 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_18 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_18 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_18 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_18 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_18 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_18 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_18 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_18 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_18 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_18 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_18 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_18 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_18 = stq_30_bits_addr_valid;
      default:
        casez_tmp_18 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_19 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_19 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_19 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_19 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_19 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_19 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_19 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_19 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_19 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_19 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_19 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_19 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_19 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_19 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_19 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_19 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_19 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_19 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_19 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_19 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_19 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_19 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_19 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_19 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_19 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_19 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_19 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_19 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_19 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_19 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_19 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_19 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_0)
      5'b00000:
        casez_tmp_20 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_20 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_20 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_20 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_20 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_20 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_20 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_20 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_20 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_20 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_20 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_20 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_20 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_20 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_20 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_20 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_20 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_20 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_20 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_20 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_20 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_20 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_20 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_20 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_20 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_20 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_20 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_20 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_20 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_20 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_20 = stq_30_bits_data_valid;
      default:
        casez_tmp_20 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_21 = stq_0_valid;
      5'b00001:
        casez_tmp_21 = stq_1_valid;
      5'b00010:
        casez_tmp_21 = stq_2_valid;
      5'b00011:
        casez_tmp_21 = stq_3_valid;
      5'b00100:
        casez_tmp_21 = stq_4_valid;
      5'b00101:
        casez_tmp_21 = stq_5_valid;
      5'b00110:
        casez_tmp_21 = stq_6_valid;
      5'b00111:
        casez_tmp_21 = stq_7_valid;
      5'b01000:
        casez_tmp_21 = stq_8_valid;
      5'b01001:
        casez_tmp_21 = stq_9_valid;
      5'b01010:
        casez_tmp_21 = stq_10_valid;
      5'b01011:
        casez_tmp_21 = stq_11_valid;
      5'b01100:
        casez_tmp_21 = stq_12_valid;
      5'b01101:
        casez_tmp_21 = stq_13_valid;
      5'b01110:
        casez_tmp_21 = stq_14_valid;
      5'b01111:
        casez_tmp_21 = stq_15_valid;
      5'b10000:
        casez_tmp_21 = stq_16_valid;
      5'b10001:
        casez_tmp_21 = stq_17_valid;
      5'b10010:
        casez_tmp_21 = stq_18_valid;
      5'b10011:
        casez_tmp_21 = stq_19_valid;
      5'b10100:
        casez_tmp_21 = stq_20_valid;
      5'b10101:
        casez_tmp_21 = stq_21_valid;
      5'b10110:
        casez_tmp_21 = stq_22_valid;
      5'b10111:
        casez_tmp_21 = stq_23_valid;
      5'b11000:
        casez_tmp_21 = stq_24_valid;
      5'b11001:
        casez_tmp_21 = stq_25_valid;
      5'b11010:
        casez_tmp_21 = stq_26_valid;
      5'b11011:
        casez_tmp_21 = stq_27_valid;
      5'b11100:
        casez_tmp_21 = stq_28_valid;
      5'b11101:
        casez_tmp_21 = stq_29_valid;
      5'b11110:
        casez_tmp_21 = stq_30_valid;
      default:
        casez_tmp_21 = stq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_22 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_22 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_22 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_22 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_22 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_22 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_22 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_22 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_22 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_22 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_22 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_22 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_22 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_22 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_22 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_22 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_22 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_22 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_22 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_22 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_22 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_22 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_22 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_22 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_22 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_22 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_22 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_22 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_22 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_22 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_22 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_22 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_23 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_23 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_23 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_23 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_23 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_23 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_23 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_23 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_23 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_23 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_23 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_23 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_23 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_23 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_23 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_23 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_23 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_23 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_23 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_23 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_23 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_23 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_23 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_23 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_23 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_23 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_23 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_23 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_23 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_23 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_23 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_23 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_24 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_24 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_24 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_24 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_24 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_24 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_24 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_24 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_24 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_24 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_24 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_24 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_24 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_24 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_24 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_24 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_24 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_24 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_24 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_24 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_24 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_24 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_24 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_24 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_24 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_24 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_24 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_24 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_24 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_24 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_24 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_24 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_25 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_25 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_25 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_25 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_25 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_25 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_25 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_25 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_25 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_25 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_25 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_25 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_25 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_25 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_25 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_25 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_25 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_25 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_25 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_25 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_25 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_25 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_25 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_25 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_25 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_25 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_25 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_25 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_25 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_25 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_25 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_25 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_26 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_26 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_26 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_26 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_26 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_26 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_26 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_26 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_26 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_26 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_26 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_26 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_26 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_26 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_26 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_26 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_26 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_26 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_26 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_26 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_26 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_26 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_26 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_26 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_26 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_26 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_26 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_26 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_26 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_26 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_26 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_26 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_27 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_27 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_27 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_27 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_27 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_27 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_27 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_27 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_27 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_27 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_27 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_27 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_27 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_27 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_27 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_27 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_27 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_27 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_27 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_27 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_27 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_27 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_27 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_27 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_27 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_27 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_27 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_27 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_27 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_27 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_27 = stq_30_bits_addr_valid;
      default:
        casez_tmp_27 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_28 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_28 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_28 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_28 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_28 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_28 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_28 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_28 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_28 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_28 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_28 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_28 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_28 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_28 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_28 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_28 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_28 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_28 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_28 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_28 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_28 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_28 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_28 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_28 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_28 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_28 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_28 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_28 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_28 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_28 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_28 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_28 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_incoming_idx_1)
      5'b00000:
        casez_tmp_29 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_29 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_29 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_29 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_29 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_29 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_29 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_29 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_29 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_29 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_29 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_29 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_29 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_29 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_29 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_29 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_29 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_29 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_29 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_29 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_29 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_29 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_29 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_29 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_29 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_29 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_29 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_29 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_29 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_29 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_29 = stq_30_bits_data_valid;
      default:
        casez_tmp_29 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg  [4:0]  ldq_wakeup_idx;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_30 = ldq_0_valid;
      5'b00001:
        casez_tmp_30 = ldq_1_valid;
      5'b00010:
        casez_tmp_30 = ldq_2_valid;
      5'b00011:
        casez_tmp_30 = ldq_3_valid;
      5'b00100:
        casez_tmp_30 = ldq_4_valid;
      5'b00101:
        casez_tmp_30 = ldq_5_valid;
      5'b00110:
        casez_tmp_30 = ldq_6_valid;
      5'b00111:
        casez_tmp_30 = ldq_7_valid;
      5'b01000:
        casez_tmp_30 = ldq_8_valid;
      5'b01001:
        casez_tmp_30 = ldq_9_valid;
      5'b01010:
        casez_tmp_30 = ldq_10_valid;
      5'b01011:
        casez_tmp_30 = ldq_11_valid;
      5'b01100:
        casez_tmp_30 = ldq_12_valid;
      5'b01101:
        casez_tmp_30 = ldq_13_valid;
      5'b01110:
        casez_tmp_30 = ldq_14_valid;
      5'b01111:
        casez_tmp_30 = ldq_15_valid;
      5'b10000:
        casez_tmp_30 = ldq_16_valid;
      5'b10001:
        casez_tmp_30 = ldq_17_valid;
      5'b10010:
        casez_tmp_30 = ldq_18_valid;
      5'b10011:
        casez_tmp_30 = ldq_19_valid;
      5'b10100:
        casez_tmp_30 = ldq_20_valid;
      5'b10101:
        casez_tmp_30 = ldq_21_valid;
      5'b10110:
        casez_tmp_30 = ldq_22_valid;
      5'b10111:
        casez_tmp_30 = ldq_23_valid;
      5'b11000:
        casez_tmp_30 = ldq_24_valid;
      5'b11001:
        casez_tmp_30 = ldq_25_valid;
      5'b11010:
        casez_tmp_30 = ldq_26_valid;
      5'b11011:
        casez_tmp_30 = ldq_27_valid;
      5'b11100:
        casez_tmp_30 = ldq_28_valid;
      5'b11101:
        casez_tmp_30 = ldq_29_valid;
      5'b11110:
        casez_tmp_30 = ldq_30_valid;
      default:
        casez_tmp_30 = ldq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_31 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_31 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_31 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_31 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_31 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_31 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_31 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_31 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_31 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_31 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_31 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_31 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_31 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_31 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_31 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_31 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_31 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_31 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_31 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_31 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_31 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_31 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_31 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_31 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_31 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_31 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_31 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_31 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_31 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_31 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_31 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_31 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_32 = ldq_0_bits_succeeded;
      5'b00001:
        casez_tmp_32 = ldq_1_bits_succeeded;
      5'b00010:
        casez_tmp_32 = ldq_2_bits_succeeded;
      5'b00011:
        casez_tmp_32 = ldq_3_bits_succeeded;
      5'b00100:
        casez_tmp_32 = ldq_4_bits_succeeded;
      5'b00101:
        casez_tmp_32 = ldq_5_bits_succeeded;
      5'b00110:
        casez_tmp_32 = ldq_6_bits_succeeded;
      5'b00111:
        casez_tmp_32 = ldq_7_bits_succeeded;
      5'b01000:
        casez_tmp_32 = ldq_8_bits_succeeded;
      5'b01001:
        casez_tmp_32 = ldq_9_bits_succeeded;
      5'b01010:
        casez_tmp_32 = ldq_10_bits_succeeded;
      5'b01011:
        casez_tmp_32 = ldq_11_bits_succeeded;
      5'b01100:
        casez_tmp_32 = ldq_12_bits_succeeded;
      5'b01101:
        casez_tmp_32 = ldq_13_bits_succeeded;
      5'b01110:
        casez_tmp_32 = ldq_14_bits_succeeded;
      5'b01111:
        casez_tmp_32 = ldq_15_bits_succeeded;
      5'b10000:
        casez_tmp_32 = ldq_16_bits_succeeded;
      5'b10001:
        casez_tmp_32 = ldq_17_bits_succeeded;
      5'b10010:
        casez_tmp_32 = ldq_18_bits_succeeded;
      5'b10011:
        casez_tmp_32 = ldq_19_bits_succeeded;
      5'b10100:
        casez_tmp_32 = ldq_20_bits_succeeded;
      5'b10101:
        casez_tmp_32 = ldq_21_bits_succeeded;
      5'b10110:
        casez_tmp_32 = ldq_22_bits_succeeded;
      5'b10111:
        casez_tmp_32 = ldq_23_bits_succeeded;
      5'b11000:
        casez_tmp_32 = ldq_24_bits_succeeded;
      5'b11001:
        casez_tmp_32 = ldq_25_bits_succeeded;
      5'b11010:
        casez_tmp_32 = ldq_26_bits_succeeded;
      5'b11011:
        casez_tmp_32 = ldq_27_bits_succeeded;
      5'b11100:
        casez_tmp_32 = ldq_28_bits_succeeded;
      5'b11101:
        casez_tmp_32 = ldq_29_bits_succeeded;
      5'b11110:
        casez_tmp_32 = ldq_30_bits_succeeded;
      default:
        casez_tmp_32 = ldq_31_bits_succeeded;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_33 = ldq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_33 = ldq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_33 = ldq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_33 = ldq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_33 = ldq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_33 = ldq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_33 = ldq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_33 = ldq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_33 = ldq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_33 = ldq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_33 = ldq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_33 = ldq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_33 = ldq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_33 = ldq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_33 = ldq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_33 = ldq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_33 = ldq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_33 = ldq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_33 = ldq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_33 = ldq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_33 = ldq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_33 = ldq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_33 = ldq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_33 = ldq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_33 = ldq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_33 = ldq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_33 = ldq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_33 = ldq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_33 = ldq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_33 = ldq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_33 = ldq_30_bits_addr_is_virtual;
      default:
        casez_tmp_33 = ldq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_34 = ldq_0_bits_executed;
      5'b00001:
        casez_tmp_34 = ldq_1_bits_executed;
      5'b00010:
        casez_tmp_34 = ldq_2_bits_executed;
      5'b00011:
        casez_tmp_34 = ldq_3_bits_executed;
      5'b00100:
        casez_tmp_34 = ldq_4_bits_executed;
      5'b00101:
        casez_tmp_34 = ldq_5_bits_executed;
      5'b00110:
        casez_tmp_34 = ldq_6_bits_executed;
      5'b00111:
        casez_tmp_34 = ldq_7_bits_executed;
      5'b01000:
        casez_tmp_34 = ldq_8_bits_executed;
      5'b01001:
        casez_tmp_34 = ldq_9_bits_executed;
      5'b01010:
        casez_tmp_34 = ldq_10_bits_executed;
      5'b01011:
        casez_tmp_34 = ldq_11_bits_executed;
      5'b01100:
        casez_tmp_34 = ldq_12_bits_executed;
      5'b01101:
        casez_tmp_34 = ldq_13_bits_executed;
      5'b01110:
        casez_tmp_34 = ldq_14_bits_executed;
      5'b01111:
        casez_tmp_34 = ldq_15_bits_executed;
      5'b10000:
        casez_tmp_34 = ldq_16_bits_executed;
      5'b10001:
        casez_tmp_34 = ldq_17_bits_executed;
      5'b10010:
        casez_tmp_34 = ldq_18_bits_executed;
      5'b10011:
        casez_tmp_34 = ldq_19_bits_executed;
      5'b10100:
        casez_tmp_34 = ldq_20_bits_executed;
      5'b10101:
        casez_tmp_34 = ldq_21_bits_executed;
      5'b10110:
        casez_tmp_34 = ldq_22_bits_executed;
      5'b10111:
        casez_tmp_34 = ldq_23_bits_executed;
      5'b11000:
        casez_tmp_34 = ldq_24_bits_executed;
      5'b11001:
        casez_tmp_34 = ldq_25_bits_executed;
      5'b11010:
        casez_tmp_34 = ldq_26_bits_executed;
      5'b11011:
        casez_tmp_34 = ldq_27_bits_executed;
      5'b11100:
        casez_tmp_34 = ldq_28_bits_executed;
      5'b11101:
        casez_tmp_34 = ldq_29_bits_executed;
      5'b11110:
        casez_tmp_34 = ldq_30_bits_executed;
      default:
        casez_tmp_34 = ldq_31_bits_executed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_35 = ldq_0_bits_order_fail;
      5'b00001:
        casez_tmp_35 = ldq_1_bits_order_fail;
      5'b00010:
        casez_tmp_35 = ldq_2_bits_order_fail;
      5'b00011:
        casez_tmp_35 = ldq_3_bits_order_fail;
      5'b00100:
        casez_tmp_35 = ldq_4_bits_order_fail;
      5'b00101:
        casez_tmp_35 = ldq_5_bits_order_fail;
      5'b00110:
        casez_tmp_35 = ldq_6_bits_order_fail;
      5'b00111:
        casez_tmp_35 = ldq_7_bits_order_fail;
      5'b01000:
        casez_tmp_35 = ldq_8_bits_order_fail;
      5'b01001:
        casez_tmp_35 = ldq_9_bits_order_fail;
      5'b01010:
        casez_tmp_35 = ldq_10_bits_order_fail;
      5'b01011:
        casez_tmp_35 = ldq_11_bits_order_fail;
      5'b01100:
        casez_tmp_35 = ldq_12_bits_order_fail;
      5'b01101:
        casez_tmp_35 = ldq_13_bits_order_fail;
      5'b01110:
        casez_tmp_35 = ldq_14_bits_order_fail;
      5'b01111:
        casez_tmp_35 = ldq_15_bits_order_fail;
      5'b10000:
        casez_tmp_35 = ldq_16_bits_order_fail;
      5'b10001:
        casez_tmp_35 = ldq_17_bits_order_fail;
      5'b10010:
        casez_tmp_35 = ldq_18_bits_order_fail;
      5'b10011:
        casez_tmp_35 = ldq_19_bits_order_fail;
      5'b10100:
        casez_tmp_35 = ldq_20_bits_order_fail;
      5'b10101:
        casez_tmp_35 = ldq_21_bits_order_fail;
      5'b10110:
        casez_tmp_35 = ldq_22_bits_order_fail;
      5'b10111:
        casez_tmp_35 = ldq_23_bits_order_fail;
      5'b11000:
        casez_tmp_35 = ldq_24_bits_order_fail;
      5'b11001:
        casez_tmp_35 = ldq_25_bits_order_fail;
      5'b11010:
        casez_tmp_35 = ldq_26_bits_order_fail;
      5'b11011:
        casez_tmp_35 = ldq_27_bits_order_fail;
      5'b11100:
        casez_tmp_35 = ldq_28_bits_order_fail;
      5'b11101:
        casez_tmp_35 = ldq_29_bits_order_fail;
      5'b11110:
        casez_tmp_35 = ldq_30_bits_order_fail;
      default:
        casez_tmp_35 = ldq_31_bits_order_fail;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_36 = p1_block_load_mask_0;
      5'b00001:
        casez_tmp_36 = p1_block_load_mask_1;
      5'b00010:
        casez_tmp_36 = p1_block_load_mask_2;
      5'b00011:
        casez_tmp_36 = p1_block_load_mask_3;
      5'b00100:
        casez_tmp_36 = p1_block_load_mask_4;
      5'b00101:
        casez_tmp_36 = p1_block_load_mask_5;
      5'b00110:
        casez_tmp_36 = p1_block_load_mask_6;
      5'b00111:
        casez_tmp_36 = p1_block_load_mask_7;
      5'b01000:
        casez_tmp_36 = p1_block_load_mask_8;
      5'b01001:
        casez_tmp_36 = p1_block_load_mask_9;
      5'b01010:
        casez_tmp_36 = p1_block_load_mask_10;
      5'b01011:
        casez_tmp_36 = p1_block_load_mask_11;
      5'b01100:
        casez_tmp_36 = p1_block_load_mask_12;
      5'b01101:
        casez_tmp_36 = p1_block_load_mask_13;
      5'b01110:
        casez_tmp_36 = p1_block_load_mask_14;
      5'b01111:
        casez_tmp_36 = p1_block_load_mask_15;
      5'b10000:
        casez_tmp_36 = p1_block_load_mask_16;
      5'b10001:
        casez_tmp_36 = p1_block_load_mask_17;
      5'b10010:
        casez_tmp_36 = p1_block_load_mask_18;
      5'b10011:
        casez_tmp_36 = p1_block_load_mask_19;
      5'b10100:
        casez_tmp_36 = p1_block_load_mask_20;
      5'b10101:
        casez_tmp_36 = p1_block_load_mask_21;
      5'b10110:
        casez_tmp_36 = p1_block_load_mask_22;
      5'b10111:
        casez_tmp_36 = p1_block_load_mask_23;
      5'b11000:
        casez_tmp_36 = p1_block_load_mask_24;
      5'b11001:
        casez_tmp_36 = p1_block_load_mask_25;
      5'b11010:
        casez_tmp_36 = p1_block_load_mask_26;
      5'b11011:
        casez_tmp_36 = p1_block_load_mask_27;
      5'b11100:
        casez_tmp_36 = p1_block_load_mask_28;
      5'b11101:
        casez_tmp_36 = p1_block_load_mask_29;
      5'b11110:
        casez_tmp_36 = p1_block_load_mask_30;
      default:
        casez_tmp_36 = p1_block_load_mask_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_37 = p2_block_load_mask_0;
      5'b00001:
        casez_tmp_37 = p2_block_load_mask_1;
      5'b00010:
        casez_tmp_37 = p2_block_load_mask_2;
      5'b00011:
        casez_tmp_37 = p2_block_load_mask_3;
      5'b00100:
        casez_tmp_37 = p2_block_load_mask_4;
      5'b00101:
        casez_tmp_37 = p2_block_load_mask_5;
      5'b00110:
        casez_tmp_37 = p2_block_load_mask_6;
      5'b00111:
        casez_tmp_37 = p2_block_load_mask_7;
      5'b01000:
        casez_tmp_37 = p2_block_load_mask_8;
      5'b01001:
        casez_tmp_37 = p2_block_load_mask_9;
      5'b01010:
        casez_tmp_37 = p2_block_load_mask_10;
      5'b01011:
        casez_tmp_37 = p2_block_load_mask_11;
      5'b01100:
        casez_tmp_37 = p2_block_load_mask_12;
      5'b01101:
        casez_tmp_37 = p2_block_load_mask_13;
      5'b01110:
        casez_tmp_37 = p2_block_load_mask_14;
      5'b01111:
        casez_tmp_37 = p2_block_load_mask_15;
      5'b10000:
        casez_tmp_37 = p2_block_load_mask_16;
      5'b10001:
        casez_tmp_37 = p2_block_load_mask_17;
      5'b10010:
        casez_tmp_37 = p2_block_load_mask_18;
      5'b10011:
        casez_tmp_37 = p2_block_load_mask_19;
      5'b10100:
        casez_tmp_37 = p2_block_load_mask_20;
      5'b10101:
        casez_tmp_37 = p2_block_load_mask_21;
      5'b10110:
        casez_tmp_37 = p2_block_load_mask_22;
      5'b10111:
        casez_tmp_37 = p2_block_load_mask_23;
      5'b11000:
        casez_tmp_37 = p2_block_load_mask_24;
      5'b11001:
        casez_tmp_37 = p2_block_load_mask_25;
      5'b11010:
        casez_tmp_37 = p2_block_load_mask_26;
      5'b11011:
        casez_tmp_37 = p2_block_load_mask_27;
      5'b11100:
        casez_tmp_37 = p2_block_load_mask_28;
      5'b11101:
        casez_tmp_37 = p2_block_load_mask_29;
      5'b11110:
        casez_tmp_37 = p2_block_load_mask_30;
      default:
        casez_tmp_37 = p2_block_load_mask_31;
    endcase
  end // always @(*)
  wire        _GEN_139807 = casez_tmp_2 & ~io_dmem_ordered;
  wire        store_needs_order = _GEN & _GEN_139807;
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_38 = ldq_0_bits_addr_is_uncacheable;
      5'b00001:
        casez_tmp_38 = ldq_1_bits_addr_is_uncacheable;
      5'b00010:
        casez_tmp_38 = ldq_2_bits_addr_is_uncacheable;
      5'b00011:
        casez_tmp_38 = ldq_3_bits_addr_is_uncacheable;
      5'b00100:
        casez_tmp_38 = ldq_4_bits_addr_is_uncacheable;
      5'b00101:
        casez_tmp_38 = ldq_5_bits_addr_is_uncacheable;
      5'b00110:
        casez_tmp_38 = ldq_6_bits_addr_is_uncacheable;
      5'b00111:
        casez_tmp_38 = ldq_7_bits_addr_is_uncacheable;
      5'b01000:
        casez_tmp_38 = ldq_8_bits_addr_is_uncacheable;
      5'b01001:
        casez_tmp_38 = ldq_9_bits_addr_is_uncacheable;
      5'b01010:
        casez_tmp_38 = ldq_10_bits_addr_is_uncacheable;
      5'b01011:
        casez_tmp_38 = ldq_11_bits_addr_is_uncacheable;
      5'b01100:
        casez_tmp_38 = ldq_12_bits_addr_is_uncacheable;
      5'b01101:
        casez_tmp_38 = ldq_13_bits_addr_is_uncacheable;
      5'b01110:
        casez_tmp_38 = ldq_14_bits_addr_is_uncacheable;
      5'b01111:
        casez_tmp_38 = ldq_15_bits_addr_is_uncacheable;
      5'b10000:
        casez_tmp_38 = ldq_16_bits_addr_is_uncacheable;
      5'b10001:
        casez_tmp_38 = ldq_17_bits_addr_is_uncacheable;
      5'b10010:
        casez_tmp_38 = ldq_18_bits_addr_is_uncacheable;
      5'b10011:
        casez_tmp_38 = ldq_19_bits_addr_is_uncacheable;
      5'b10100:
        casez_tmp_38 = ldq_20_bits_addr_is_uncacheable;
      5'b10101:
        casez_tmp_38 = ldq_21_bits_addr_is_uncacheable;
      5'b10110:
        casez_tmp_38 = ldq_22_bits_addr_is_uncacheable;
      5'b10111:
        casez_tmp_38 = ldq_23_bits_addr_is_uncacheable;
      5'b11000:
        casez_tmp_38 = ldq_24_bits_addr_is_uncacheable;
      5'b11001:
        casez_tmp_38 = ldq_25_bits_addr_is_uncacheable;
      5'b11010:
        casez_tmp_38 = ldq_26_bits_addr_is_uncacheable;
      5'b11011:
        casez_tmp_38 = ldq_27_bits_addr_is_uncacheable;
      5'b11100:
        casez_tmp_38 = ldq_28_bits_addr_is_uncacheable;
      5'b11101:
        casez_tmp_38 = ldq_29_bits_addr_is_uncacheable;
      5'b11110:
        casez_tmp_38 = ldq_30_bits_addr_is_uncacheable;
      default:
        casez_tmp_38 = ldq_31_bits_addr_is_uncacheable;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_39 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_39 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_39 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_39 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_39 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_39 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_39 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_39 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_39 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_39 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_39 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_39 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_39 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_39 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_39 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_39 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_39 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_39 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_39 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_39 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_39 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_39 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_39 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_39 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_39 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_39 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_39 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_39 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_39 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_39 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_39 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_39 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  wire        can_fire_load_incoming_1 = exe_req_1_valid & exe_req_1_bits_uop_ctrl_is_load;
  wire        _can_fire_sta_incoming_T_3 = exe_req_1_valid & exe_req_1_bits_uop_ctrl_is_sta;
  wire        will_fire_stad_incoming_1 = _can_fire_sta_incoming_T_3 & exe_req_1_bits_uop_ctrl_is_std & ~can_fire_load_incoming_1 & ~can_fire_load_incoming_1;
  wire        _will_fire_sta_incoming_1_will_fire_T_2 = ~can_fire_load_incoming_1 & ~will_fire_stad_incoming_1;
  wire        _will_fire_sta_incoming_1_will_fire_T_6 = ~can_fire_load_incoming_1 & ~will_fire_stad_incoming_1;
  wire        will_fire_sta_incoming_1 = _can_fire_sta_incoming_T_3 & ~exe_req_1_bits_uop_ctrl_is_std & _will_fire_sta_incoming_1_will_fire_T_2 & _will_fire_sta_incoming_1_will_fire_T_6 & ~will_fire_stad_incoming_1;
  wire        _will_fire_sfence_1_will_fire_T_2 = _will_fire_sta_incoming_1_will_fire_T_2 & ~will_fire_sta_incoming_1;
  wire        _will_fire_release_1_will_fire_T_6 = _will_fire_sta_incoming_1_will_fire_T_6 & ~will_fire_sta_incoming_1;
  wire        _will_fire_std_incoming_1_will_fire_T_14 = ~will_fire_stad_incoming_1 & ~will_fire_sta_incoming_1;
  wire        will_fire_std_incoming_1 = exe_req_1_valid & exe_req_1_bits_uop_ctrl_is_std & ~exe_req_1_bits_uop_ctrl_is_sta & _will_fire_std_incoming_1_will_fire_T_14;
  wire        _will_fire_sfence_1_will_fire_T_14 = _will_fire_std_incoming_1_will_fire_T_14 & ~will_fire_std_incoming_1;
  wire        will_fire_sfence_1 = exe_req_1_valid & exe_req_1_bits_sfence_valid & _will_fire_sfence_1_will_fire_T_2 & _will_fire_sfence_1_will_fire_T_14;
  wire        _will_fire_hella_incoming_1_will_fire_T_2 = _will_fire_sfence_1_will_fire_T_2 & ~will_fire_sfence_1;
  wire        will_fire_release_1 = io_dmem_release_valid & _will_fire_release_1_will_fire_T_6;
  wire        _GEN_140251 = hella_state == 3'h1;
  wire        _will_fire_load_retry_1_will_fire_T_6 = _will_fire_release_1_will_fire_T_6 & ~will_fire_release_1;
  wire        will_fire_hella_incoming_1 = (|hella_state) & _GEN_140251 & _will_fire_hella_incoming_1_will_fire_T_2 & ~can_fire_load_incoming_1;
  wire        _will_fire_load_retry_1_will_fire_T_2 = _will_fire_hella_incoming_1_will_fire_T_2 & ~will_fire_hella_incoming_1;
  wire        _GEN_140233 = hella_state == 3'h3;
  wire        _GEN_330 = hella_state == 3'h2;
  wire        _GEN_331 = hella_state == 3'h4;
  wire        _GEN_140205 = hella_state == 3'h5;
  wire        _will_fire_hella_wakeup_1_will_fire_T_10 = ~can_fire_load_incoming_1 & ~will_fire_hella_incoming_1;
  wire        will_fire_hella_wakeup_1 = ~(~(|hella_state) | _GEN_140251 | _GEN_140233 | _GEN_330 | _GEN_331) & _GEN_140205 & _will_fire_hella_wakeup_1_will_fire_T_10;
  reg  [4:0]  ldq_retry_idx;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_40 = ldq_0_valid;
      5'b00001:
        casez_tmp_40 = ldq_1_valid;
      5'b00010:
        casez_tmp_40 = ldq_2_valid;
      5'b00011:
        casez_tmp_40 = ldq_3_valid;
      5'b00100:
        casez_tmp_40 = ldq_4_valid;
      5'b00101:
        casez_tmp_40 = ldq_5_valid;
      5'b00110:
        casez_tmp_40 = ldq_6_valid;
      5'b00111:
        casez_tmp_40 = ldq_7_valid;
      5'b01000:
        casez_tmp_40 = ldq_8_valid;
      5'b01001:
        casez_tmp_40 = ldq_9_valid;
      5'b01010:
        casez_tmp_40 = ldq_10_valid;
      5'b01011:
        casez_tmp_40 = ldq_11_valid;
      5'b01100:
        casez_tmp_40 = ldq_12_valid;
      5'b01101:
        casez_tmp_40 = ldq_13_valid;
      5'b01110:
        casez_tmp_40 = ldq_14_valid;
      5'b01111:
        casez_tmp_40 = ldq_15_valid;
      5'b10000:
        casez_tmp_40 = ldq_16_valid;
      5'b10001:
        casez_tmp_40 = ldq_17_valid;
      5'b10010:
        casez_tmp_40 = ldq_18_valid;
      5'b10011:
        casez_tmp_40 = ldq_19_valid;
      5'b10100:
        casez_tmp_40 = ldq_20_valid;
      5'b10101:
        casez_tmp_40 = ldq_21_valid;
      5'b10110:
        casez_tmp_40 = ldq_22_valid;
      5'b10111:
        casez_tmp_40 = ldq_23_valid;
      5'b11000:
        casez_tmp_40 = ldq_24_valid;
      5'b11001:
        casez_tmp_40 = ldq_25_valid;
      5'b11010:
        casez_tmp_40 = ldq_26_valid;
      5'b11011:
        casez_tmp_40 = ldq_27_valid;
      5'b11100:
        casez_tmp_40 = ldq_28_valid;
      5'b11101:
        casez_tmp_40 = ldq_29_valid;
      5'b11110:
        casez_tmp_40 = ldq_30_valid;
      default:
        casez_tmp_40 = ldq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_41 = ldq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_41 = ldq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_41 = ldq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_41 = ldq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_41 = ldq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_41 = ldq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_41 = ldq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_41 = ldq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_41 = ldq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_41 = ldq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_41 = ldq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_41 = ldq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_41 = ldq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_41 = ldq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_41 = ldq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_41 = ldq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_41 = ldq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_41 = ldq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_41 = ldq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_41 = ldq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_41 = ldq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_41 = ldq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_41 = ldq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_41 = ldq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_41 = ldq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_41 = ldq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_41 = ldq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_41 = ldq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_41 = ldq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_41 = ldq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_41 = ldq_30_bits_addr_valid;
      default:
        casez_tmp_41 = ldq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_42 = ldq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_42 = ldq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_42 = ldq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_42 = ldq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_42 = ldq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_42 = ldq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_42 = ldq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_42 = ldq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_42 = ldq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_42 = ldq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_42 = ldq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_42 = ldq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_42 = ldq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_42 = ldq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_42 = ldq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_42 = ldq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_42 = ldq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_42 = ldq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_42 = ldq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_42 = ldq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_42 = ldq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_42 = ldq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_42 = ldq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_42 = ldq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_42 = ldq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_42 = ldq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_42 = ldq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_42 = ldq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_42 = ldq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_42 = ldq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_42 = ldq_30_bits_addr_is_virtual;
      default:
        casez_tmp_42 = ldq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_43 = p1_block_load_mask_0;
      5'b00001:
        casez_tmp_43 = p1_block_load_mask_1;
      5'b00010:
        casez_tmp_43 = p1_block_load_mask_2;
      5'b00011:
        casez_tmp_43 = p1_block_load_mask_3;
      5'b00100:
        casez_tmp_43 = p1_block_load_mask_4;
      5'b00101:
        casez_tmp_43 = p1_block_load_mask_5;
      5'b00110:
        casez_tmp_43 = p1_block_load_mask_6;
      5'b00111:
        casez_tmp_43 = p1_block_load_mask_7;
      5'b01000:
        casez_tmp_43 = p1_block_load_mask_8;
      5'b01001:
        casez_tmp_43 = p1_block_load_mask_9;
      5'b01010:
        casez_tmp_43 = p1_block_load_mask_10;
      5'b01011:
        casez_tmp_43 = p1_block_load_mask_11;
      5'b01100:
        casez_tmp_43 = p1_block_load_mask_12;
      5'b01101:
        casez_tmp_43 = p1_block_load_mask_13;
      5'b01110:
        casez_tmp_43 = p1_block_load_mask_14;
      5'b01111:
        casez_tmp_43 = p1_block_load_mask_15;
      5'b10000:
        casez_tmp_43 = p1_block_load_mask_16;
      5'b10001:
        casez_tmp_43 = p1_block_load_mask_17;
      5'b10010:
        casez_tmp_43 = p1_block_load_mask_18;
      5'b10011:
        casez_tmp_43 = p1_block_load_mask_19;
      5'b10100:
        casez_tmp_43 = p1_block_load_mask_20;
      5'b10101:
        casez_tmp_43 = p1_block_load_mask_21;
      5'b10110:
        casez_tmp_43 = p1_block_load_mask_22;
      5'b10111:
        casez_tmp_43 = p1_block_load_mask_23;
      5'b11000:
        casez_tmp_43 = p1_block_load_mask_24;
      5'b11001:
        casez_tmp_43 = p1_block_load_mask_25;
      5'b11010:
        casez_tmp_43 = p1_block_load_mask_26;
      5'b11011:
        casez_tmp_43 = p1_block_load_mask_27;
      5'b11100:
        casez_tmp_43 = p1_block_load_mask_28;
      5'b11101:
        casez_tmp_43 = p1_block_load_mask_29;
      5'b11110:
        casez_tmp_43 = p1_block_load_mask_30;
      default:
        casez_tmp_43 = p1_block_load_mask_31;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_44 = p2_block_load_mask_0;
      5'b00001:
        casez_tmp_44 = p2_block_load_mask_1;
      5'b00010:
        casez_tmp_44 = p2_block_load_mask_2;
      5'b00011:
        casez_tmp_44 = p2_block_load_mask_3;
      5'b00100:
        casez_tmp_44 = p2_block_load_mask_4;
      5'b00101:
        casez_tmp_44 = p2_block_load_mask_5;
      5'b00110:
        casez_tmp_44 = p2_block_load_mask_6;
      5'b00111:
        casez_tmp_44 = p2_block_load_mask_7;
      5'b01000:
        casez_tmp_44 = p2_block_load_mask_8;
      5'b01001:
        casez_tmp_44 = p2_block_load_mask_9;
      5'b01010:
        casez_tmp_44 = p2_block_load_mask_10;
      5'b01011:
        casez_tmp_44 = p2_block_load_mask_11;
      5'b01100:
        casez_tmp_44 = p2_block_load_mask_12;
      5'b01101:
        casez_tmp_44 = p2_block_load_mask_13;
      5'b01110:
        casez_tmp_44 = p2_block_load_mask_14;
      5'b01111:
        casez_tmp_44 = p2_block_load_mask_15;
      5'b10000:
        casez_tmp_44 = p2_block_load_mask_16;
      5'b10001:
        casez_tmp_44 = p2_block_load_mask_17;
      5'b10010:
        casez_tmp_44 = p2_block_load_mask_18;
      5'b10011:
        casez_tmp_44 = p2_block_load_mask_19;
      5'b10100:
        casez_tmp_44 = p2_block_load_mask_20;
      5'b10101:
        casez_tmp_44 = p2_block_load_mask_21;
      5'b10110:
        casez_tmp_44 = p2_block_load_mask_22;
      5'b10111:
        casez_tmp_44 = p2_block_load_mask_23;
      5'b11000:
        casez_tmp_44 = p2_block_load_mask_24;
      5'b11001:
        casez_tmp_44 = p2_block_load_mask_25;
      5'b11010:
        casez_tmp_44 = p2_block_load_mask_26;
      5'b11011:
        casez_tmp_44 = p2_block_load_mask_27;
      5'b11100:
        casez_tmp_44 = p2_block_load_mask_28;
      5'b11101:
        casez_tmp_44 = p2_block_load_mask_29;
      5'b11110:
        casez_tmp_44 = p2_block_load_mask_30;
      default:
        casez_tmp_44 = p2_block_load_mask_31;
    endcase
  end // always @(*)
  reg         can_fire_load_retry_REG_1;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_45 = ldq_0_bits_order_fail;
      5'b00001:
        casez_tmp_45 = ldq_1_bits_order_fail;
      5'b00010:
        casez_tmp_45 = ldq_2_bits_order_fail;
      5'b00011:
        casez_tmp_45 = ldq_3_bits_order_fail;
      5'b00100:
        casez_tmp_45 = ldq_4_bits_order_fail;
      5'b00101:
        casez_tmp_45 = ldq_5_bits_order_fail;
      5'b00110:
        casez_tmp_45 = ldq_6_bits_order_fail;
      5'b00111:
        casez_tmp_45 = ldq_7_bits_order_fail;
      5'b01000:
        casez_tmp_45 = ldq_8_bits_order_fail;
      5'b01001:
        casez_tmp_45 = ldq_9_bits_order_fail;
      5'b01010:
        casez_tmp_45 = ldq_10_bits_order_fail;
      5'b01011:
        casez_tmp_45 = ldq_11_bits_order_fail;
      5'b01100:
        casez_tmp_45 = ldq_12_bits_order_fail;
      5'b01101:
        casez_tmp_45 = ldq_13_bits_order_fail;
      5'b01110:
        casez_tmp_45 = ldq_14_bits_order_fail;
      5'b01111:
        casez_tmp_45 = ldq_15_bits_order_fail;
      5'b10000:
        casez_tmp_45 = ldq_16_bits_order_fail;
      5'b10001:
        casez_tmp_45 = ldq_17_bits_order_fail;
      5'b10010:
        casez_tmp_45 = ldq_18_bits_order_fail;
      5'b10011:
        casez_tmp_45 = ldq_19_bits_order_fail;
      5'b10100:
        casez_tmp_45 = ldq_20_bits_order_fail;
      5'b10101:
        casez_tmp_45 = ldq_21_bits_order_fail;
      5'b10110:
        casez_tmp_45 = ldq_22_bits_order_fail;
      5'b10111:
        casez_tmp_45 = ldq_23_bits_order_fail;
      5'b11000:
        casez_tmp_45 = ldq_24_bits_order_fail;
      5'b11001:
        casez_tmp_45 = ldq_25_bits_order_fail;
      5'b11010:
        casez_tmp_45 = ldq_26_bits_order_fail;
      5'b11011:
        casez_tmp_45 = ldq_27_bits_order_fail;
      5'b11100:
        casez_tmp_45 = ldq_28_bits_order_fail;
      5'b11101:
        casez_tmp_45 = ldq_29_bits_order_fail;
      5'b11110:
        casez_tmp_45 = ldq_30_bits_order_fail;
      default:
        casez_tmp_45 = ldq_31_bits_order_fail;
    endcase
  end // always @(*)
  wire        _will_fire_load_retry_1_will_fire_T_10 = _will_fire_hella_wakeup_1_will_fire_T_10 & ~will_fire_hella_wakeup_1;
  wire        will_fire_load_retry_1 = casez_tmp_40 & casez_tmp_41 & casez_tmp_42 & ~casez_tmp_43 & ~casez_tmp_44 & can_fire_load_retry_REG_1 & ~store_needs_order & ~casez_tmp_45 & _will_fire_load_retry_1_will_fire_T_2 & _will_fire_load_retry_1_will_fire_T_6 & _will_fire_load_retry_1_will_fire_T_10;
  wire        _will_fire_sta_retry_1_will_fire_T_2 = _will_fire_load_retry_1_will_fire_T_2 & ~will_fire_load_retry_1;
  reg  [4:0]  stq_retry_idx;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_46 = stq_0_valid;
      5'b00001:
        casez_tmp_46 = stq_1_valid;
      5'b00010:
        casez_tmp_46 = stq_2_valid;
      5'b00011:
        casez_tmp_46 = stq_3_valid;
      5'b00100:
        casez_tmp_46 = stq_4_valid;
      5'b00101:
        casez_tmp_46 = stq_5_valid;
      5'b00110:
        casez_tmp_46 = stq_6_valid;
      5'b00111:
        casez_tmp_46 = stq_7_valid;
      5'b01000:
        casez_tmp_46 = stq_8_valid;
      5'b01001:
        casez_tmp_46 = stq_9_valid;
      5'b01010:
        casez_tmp_46 = stq_10_valid;
      5'b01011:
        casez_tmp_46 = stq_11_valid;
      5'b01100:
        casez_tmp_46 = stq_12_valid;
      5'b01101:
        casez_tmp_46 = stq_13_valid;
      5'b01110:
        casez_tmp_46 = stq_14_valid;
      5'b01111:
        casez_tmp_46 = stq_15_valid;
      5'b10000:
        casez_tmp_46 = stq_16_valid;
      5'b10001:
        casez_tmp_46 = stq_17_valid;
      5'b10010:
        casez_tmp_46 = stq_18_valid;
      5'b10011:
        casez_tmp_46 = stq_19_valid;
      5'b10100:
        casez_tmp_46 = stq_20_valid;
      5'b10101:
        casez_tmp_46 = stq_21_valid;
      5'b10110:
        casez_tmp_46 = stq_22_valid;
      5'b10111:
        casez_tmp_46 = stq_23_valid;
      5'b11000:
        casez_tmp_46 = stq_24_valid;
      5'b11001:
        casez_tmp_46 = stq_25_valid;
      5'b11010:
        casez_tmp_46 = stq_26_valid;
      5'b11011:
        casez_tmp_46 = stq_27_valid;
      5'b11100:
        casez_tmp_46 = stq_28_valid;
      5'b11101:
        casez_tmp_46 = stq_29_valid;
      5'b11110:
        casez_tmp_46 = stq_30_valid;
      default:
        casez_tmp_46 = stq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_47 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_47 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_47 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_47 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_47 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_47 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_47 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_47 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_47 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_47 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_47 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_47 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_47 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_47 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_47 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_47 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_47 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_47 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_47 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_47 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_47 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_47 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_47 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_47 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_47 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_47 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_47 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_47 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_47 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_47 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_47 = stq_30_bits_addr_valid;
      default:
        casez_tmp_47 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_48 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_48 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_48 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_48 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_48 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_48 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_48 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_48 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_48 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_48 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_48 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_48 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_48 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_48 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_48 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_48 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_48 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_48 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_48 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_48 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_48 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_48 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_48 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_48 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_48 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_48 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_48 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_48 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_48 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_48 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_48 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_48 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  reg         can_fire_sta_retry_REG_1;
  wire        can_fire_std_incoming_0 = exe_req_0_valid & mem_incoming_uop_out_ctrl_is_std & ~mem_incoming_uop_out_ctrl_is_sta;
  wire        _will_fire_sta_retry_1_will_fire_T_6 = _will_fire_load_retry_1_will_fire_T_6 & ~will_fire_load_retry_1;
  wire        will_fire_sta_retry_1 = casez_tmp_46 & casez_tmp_47 & casez_tmp_48 & can_fire_sta_retry_REG_1 & ~(can_fire_std_incoming_0 & stq_incoming_idx_0 == stq_retry_idx) & _will_fire_sta_retry_1_will_fire_T_2 & _will_fire_sta_retry_1_will_fire_T_6 & _will_fire_sfence_1_will_fire_T_14 & ~will_fire_sfence_1;
  assign _will_fire_store_commit_1_T_2 = _will_fire_sta_retry_1_will_fire_T_2 & ~will_fire_sta_retry_1;
  wire        will_fire_load_wakeup_1 = casez_tmp_30 & casez_tmp_31 & ~casez_tmp_32 & ~casez_tmp_33 & ~casez_tmp_34 & ~casez_tmp_35 & ~casez_tmp_36 & ~casez_tmp_37 & ~store_needs_order & (~casez_tmp_38 | io_core_commit_load_at_rob_head & ldq_head == ldq_wakeup_idx & casez_tmp_39 == 32'h0) & _will_fire_sta_retry_1_will_fire_T_6 & ~will_fire_sta_retry_1 & _will_fire_load_retry_1_will_fire_T_10 & ~will_fire_load_retry_1;
  wire        can_fire_load_incoming_0 = exe_req_0_valid & mem_incoming_uop_out_ctrl_is_load;
  wire        _can_fire_sta_incoming_T = exe_req_0_valid & mem_incoming_uop_out_ctrl_is_sta;
  wire        will_fire_stad_incoming_0 = _can_fire_sta_incoming_T & mem_incoming_uop_out_ctrl_is_std & ~can_fire_load_incoming_0 & ~can_fire_load_incoming_0;
  wire        _will_fire_sta_incoming_0_will_fire_T_2 = ~can_fire_load_incoming_0 & ~will_fire_stad_incoming_0;
  wire        will_fire_sta_incoming_0 = _can_fire_sta_incoming_T & ~mem_incoming_uop_out_ctrl_is_std & _will_fire_sta_incoming_0_will_fire_T_2 & ~can_fire_load_incoming_0 & ~will_fire_stad_incoming_0 & ~will_fire_stad_incoming_0;
  wire        _will_fire_sfence_0_will_fire_T_2 = _will_fire_sta_incoming_0_will_fire_T_2 & ~will_fire_sta_incoming_0;
  wire        _will_fire_std_incoming_0_will_fire_T_14 = ~will_fire_stad_incoming_0 & ~will_fire_sta_incoming_0;
  wire        will_fire_std_incoming_0 = can_fire_std_incoming_0 & _will_fire_std_incoming_0_will_fire_T_14;
  wire        will_fire_sfence_0 = exe_req_0_valid & exe_req_0_bits_sfence_valid & _will_fire_sfence_0_will_fire_T_2 & _will_fire_std_incoming_0_will_fire_T_14 & ~will_fire_std_incoming_0;
  assign _will_fire_store_commit_0_T_2 = _will_fire_sfence_0_will_fire_T_2 & ~will_fire_sfence_0;
  wire        _temp_bits_T = ldq_head == 5'h0;
  wire        _temp_bits_T_2 = ldq_head < 5'h2;
  wire        _temp_bits_T_4 = ldq_head < 5'h3;
  wire        _temp_bits_T_6 = ldq_head < 5'h4;
  wire        _temp_bits_T_8 = ldq_head < 5'h5;
  wire        _temp_bits_T_10 = ldq_head < 5'h6;
  wire        _temp_bits_T_12 = ldq_head < 5'h7;
  wire        _temp_bits_T_14 = ldq_head < 5'h8;
  wire        _temp_bits_T_16 = ldq_head < 5'h9;
  wire        _temp_bits_T_18 = ldq_head < 5'hA;
  wire        _temp_bits_T_20 = ldq_head < 5'hB;
  wire        _temp_bits_T_22 = ldq_head < 5'hC;
  wire        _temp_bits_T_24 = ldq_head < 5'hD;
  wire        _temp_bits_T_26 = ldq_head < 5'hE;
  wire        _temp_bits_T_28 = ldq_head < 5'hF;
  wire        _temp_bits_T_32 = ldq_head < 5'h11;
  wire        _temp_bits_T_34 = ldq_head < 5'h12;
  wire        _temp_bits_T_36 = ldq_head < 5'h13;
  wire        _temp_bits_T_38 = ldq_head < 5'h14;
  wire        _temp_bits_T_40 = ldq_head < 5'h15;
  wire        _temp_bits_T_42 = ldq_head < 5'h16;
  wire        _temp_bits_T_44 = ldq_head < 5'h17;
  wire        _temp_bits_T_46 = ldq_head[4:3] != 2'h3;
  wire        _temp_bits_T_48 = ldq_head < 5'h19;
  wire        _temp_bits_T_50 = ldq_head < 5'h1A;
  wire        _temp_bits_T_52 = ldq_head < 5'h1B;
  wire        _temp_bits_T_54 = ldq_head[4:2] != 3'h7;
  wire        _temp_bits_T_56 = ldq_head < 5'h1D;
  wire        _temp_bits_T_58 = ldq_head[4:1] != 4'hF;
  wire        _temp_bits_T_60 = ldq_head != 5'h1F;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_49 = stq_0_bits_uop_is_fence;
      5'b00001:
        casez_tmp_49 = stq_1_bits_uop_is_fence;
      5'b00010:
        casez_tmp_49 = stq_2_bits_uop_is_fence;
      5'b00011:
        casez_tmp_49 = stq_3_bits_uop_is_fence;
      5'b00100:
        casez_tmp_49 = stq_4_bits_uop_is_fence;
      5'b00101:
        casez_tmp_49 = stq_5_bits_uop_is_fence;
      5'b00110:
        casez_tmp_49 = stq_6_bits_uop_is_fence;
      5'b00111:
        casez_tmp_49 = stq_7_bits_uop_is_fence;
      5'b01000:
        casez_tmp_49 = stq_8_bits_uop_is_fence;
      5'b01001:
        casez_tmp_49 = stq_9_bits_uop_is_fence;
      5'b01010:
        casez_tmp_49 = stq_10_bits_uop_is_fence;
      5'b01011:
        casez_tmp_49 = stq_11_bits_uop_is_fence;
      5'b01100:
        casez_tmp_49 = stq_12_bits_uop_is_fence;
      5'b01101:
        casez_tmp_49 = stq_13_bits_uop_is_fence;
      5'b01110:
        casez_tmp_49 = stq_14_bits_uop_is_fence;
      5'b01111:
        casez_tmp_49 = stq_15_bits_uop_is_fence;
      5'b10000:
        casez_tmp_49 = stq_16_bits_uop_is_fence;
      5'b10001:
        casez_tmp_49 = stq_17_bits_uop_is_fence;
      5'b10010:
        casez_tmp_49 = stq_18_bits_uop_is_fence;
      5'b10011:
        casez_tmp_49 = stq_19_bits_uop_is_fence;
      5'b10100:
        casez_tmp_49 = stq_20_bits_uop_is_fence;
      5'b10101:
        casez_tmp_49 = stq_21_bits_uop_is_fence;
      5'b10110:
        casez_tmp_49 = stq_22_bits_uop_is_fence;
      5'b10111:
        casez_tmp_49 = stq_23_bits_uop_is_fence;
      5'b11000:
        casez_tmp_49 = stq_24_bits_uop_is_fence;
      5'b11001:
        casez_tmp_49 = stq_25_bits_uop_is_fence;
      5'b11010:
        casez_tmp_49 = stq_26_bits_uop_is_fence;
      5'b11011:
        casez_tmp_49 = stq_27_bits_uop_is_fence;
      5'b11100:
        casez_tmp_49 = stq_28_bits_uop_is_fence;
      5'b11101:
        casez_tmp_49 = stq_29_bits_uop_is_fence;
      5'b11110:
        casez_tmp_49 = stq_30_bits_uop_is_fence;
      default:
        casez_tmp_49 = stq_31_bits_uop_is_fence;
    endcase
  end // always @(*)
  reg         mem_xcpt_valids_0;
  reg         mem_xcpt_valids_1;
  wire        mem_xcpt_valid = mem_xcpt_valids_0 | mem_xcpt_valids_1;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_50 = stq_0_bits_uop_exception;
      5'b00001:
        casez_tmp_50 = stq_1_bits_uop_exception;
      5'b00010:
        casez_tmp_50 = stq_2_bits_uop_exception;
      5'b00011:
        casez_tmp_50 = stq_3_bits_uop_exception;
      5'b00100:
        casez_tmp_50 = stq_4_bits_uop_exception;
      5'b00101:
        casez_tmp_50 = stq_5_bits_uop_exception;
      5'b00110:
        casez_tmp_50 = stq_6_bits_uop_exception;
      5'b00111:
        casez_tmp_50 = stq_7_bits_uop_exception;
      5'b01000:
        casez_tmp_50 = stq_8_bits_uop_exception;
      5'b01001:
        casez_tmp_50 = stq_9_bits_uop_exception;
      5'b01010:
        casez_tmp_50 = stq_10_bits_uop_exception;
      5'b01011:
        casez_tmp_50 = stq_11_bits_uop_exception;
      5'b01100:
        casez_tmp_50 = stq_12_bits_uop_exception;
      5'b01101:
        casez_tmp_50 = stq_13_bits_uop_exception;
      5'b01110:
        casez_tmp_50 = stq_14_bits_uop_exception;
      5'b01111:
        casez_tmp_50 = stq_15_bits_uop_exception;
      5'b10000:
        casez_tmp_50 = stq_16_bits_uop_exception;
      5'b10001:
        casez_tmp_50 = stq_17_bits_uop_exception;
      5'b10010:
        casez_tmp_50 = stq_18_bits_uop_exception;
      5'b10011:
        casez_tmp_50 = stq_19_bits_uop_exception;
      5'b10100:
        casez_tmp_50 = stq_20_bits_uop_exception;
      5'b10101:
        casez_tmp_50 = stq_21_bits_uop_exception;
      5'b10110:
        casez_tmp_50 = stq_22_bits_uop_exception;
      5'b10111:
        casez_tmp_50 = stq_23_bits_uop_exception;
      5'b11000:
        casez_tmp_50 = stq_24_bits_uop_exception;
      5'b11001:
        casez_tmp_50 = stq_25_bits_uop_exception;
      5'b11010:
        casez_tmp_50 = stq_26_bits_uop_exception;
      5'b11011:
        casez_tmp_50 = stq_27_bits_uop_exception;
      5'b11100:
        casez_tmp_50 = stq_28_bits_uop_exception;
      5'b11101:
        casez_tmp_50 = stq_29_bits_uop_exception;
      5'b11110:
        casez_tmp_50 = stq_30_bits_uop_exception;
      default:
        casez_tmp_50 = stq_31_bits_uop_exception;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_51 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_51 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_51 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_51 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_51 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_51 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_51 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_51 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_51 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_51 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_51 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_51 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_51 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_51 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_51 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_51 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_51 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_51 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_51 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_51 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_51 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_51 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_51 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_51 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_51 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_51 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_51 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_51 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_51 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_51 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_51 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_51 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_52 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_52 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_52 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_52 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_52 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_52 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_52 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_52 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_52 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_52 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_52 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_52 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_52 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_52 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_52 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_52 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_52 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_52 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_52 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_52 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_52 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_52 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_52 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_52 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_52 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_52 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_52 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_52 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_52 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_52 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_52 = stq_30_bits_addr_valid;
      default:
        casez_tmp_52 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_53 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_53 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_53 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_53 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_53 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_53 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_53 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_53 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_53 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_53 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_53 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_53 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_53 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_53 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_53 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_53 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_53 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_53 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_53 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_53 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_53 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_53 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_53 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_53 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_53 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_53 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_53 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_53 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_53 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_53 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_53 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_53 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_54 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_54 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_54 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_54 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_54 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_54 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_54 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_54 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_54 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_54 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_54 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_54 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_54 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_54 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_54 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_54 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_54 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_54 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_54 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_54 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_54 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_54 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_54 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_54 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_54 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_54 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_54 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_54 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_54 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_54 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_54 = stq_30_bits_data_valid;
      default:
        casez_tmp_54 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_55 = stq_0_bits_committed;
      5'b00001:
        casez_tmp_55 = stq_1_bits_committed;
      5'b00010:
        casez_tmp_55 = stq_2_bits_committed;
      5'b00011:
        casez_tmp_55 = stq_3_bits_committed;
      5'b00100:
        casez_tmp_55 = stq_4_bits_committed;
      5'b00101:
        casez_tmp_55 = stq_5_bits_committed;
      5'b00110:
        casez_tmp_55 = stq_6_bits_committed;
      5'b00111:
        casez_tmp_55 = stq_7_bits_committed;
      5'b01000:
        casez_tmp_55 = stq_8_bits_committed;
      5'b01001:
        casez_tmp_55 = stq_9_bits_committed;
      5'b01010:
        casez_tmp_55 = stq_10_bits_committed;
      5'b01011:
        casez_tmp_55 = stq_11_bits_committed;
      5'b01100:
        casez_tmp_55 = stq_12_bits_committed;
      5'b01101:
        casez_tmp_55 = stq_13_bits_committed;
      5'b01110:
        casez_tmp_55 = stq_14_bits_committed;
      5'b01111:
        casez_tmp_55 = stq_15_bits_committed;
      5'b10000:
        casez_tmp_55 = stq_16_bits_committed;
      5'b10001:
        casez_tmp_55 = stq_17_bits_committed;
      5'b10010:
        casez_tmp_55 = stq_18_bits_committed;
      5'b10011:
        casez_tmp_55 = stq_19_bits_committed;
      5'b10100:
        casez_tmp_55 = stq_20_bits_committed;
      5'b10101:
        casez_tmp_55 = stq_21_bits_committed;
      5'b10110:
        casez_tmp_55 = stq_22_bits_committed;
      5'b10111:
        casez_tmp_55 = stq_23_bits_committed;
      5'b11000:
        casez_tmp_55 = stq_24_bits_committed;
      5'b11001:
        casez_tmp_55 = stq_25_bits_committed;
      5'b11010:
        casez_tmp_55 = stq_26_bits_committed;
      5'b11011:
        casez_tmp_55 = stq_27_bits_committed;
      5'b11100:
        casez_tmp_55 = stq_28_bits_committed;
      5'b11101:
        casez_tmp_55 = stq_29_bits_committed;
      5'b11110:
        casez_tmp_55 = stq_30_bits_committed;
      default:
        casez_tmp_55 = stq_31_bits_committed;
    endcase
  end // always @(*)
  wire        will_fire_store_commit_0 = casez_tmp & ~casez_tmp_49 & ~mem_xcpt_valid & ~casez_tmp_50 & (casez_tmp_55 | casez_tmp_51 & casez_tmp_52 & ~casez_tmp_53 & casez_tmp_54) & ~can_fire_load_incoming_0;
  wire        _exe_cmd_T = can_fire_load_incoming_0 | will_fire_stad_incoming_0;
  wire        _exe_cmd_T_7 = can_fire_load_incoming_1 | will_fire_stad_incoming_1;
  wire        _exe_tlb_uop_T_2 = _exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_56 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_56 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_56 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_56 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_56 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_56 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_56 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_56 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_56 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_56 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_56 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_56 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_56 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_56 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_56 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_56 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_56 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_56 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_56 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_56 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_56 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_56 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_56 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_56 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_56 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_56 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_56 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_56 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_56 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_56 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_56 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_56 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_57 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_57 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_57 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_57 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_57 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_57 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_57 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_57 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_57 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_57 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_57 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_57 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_57 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_57 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_57 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_57 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_57 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_57 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_57 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_57 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_57 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_57 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_57 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_57 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_57 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_57 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_57 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_57 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_57 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_57 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_57 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_57 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_58 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_58 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_58 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_58 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_58 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_58 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_58 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_58 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_58 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_58 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_58 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_58 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_58 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_58 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_58 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_58 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_58 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_58 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_58 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_58 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_58 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_58 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_58 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_58 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_58 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_58 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_58 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_58 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_58 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_58 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_58 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_58 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_59 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_59 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_59 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_59 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_59 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_59 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_59 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_59 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_59 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_59 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_59 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_59 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_59 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_59 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_59 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_59 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_59 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_59 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_59 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_59 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_59 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_59 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_59 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_59 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_59 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_59 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_59 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_59 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_59 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_59 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_59 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_59 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_60 = stq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_60 = stq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_60 = stq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_60 = stq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_60 = stq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_60 = stq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_60 = stq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_60 = stq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_60 = stq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_60 = stq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_60 = stq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_60 = stq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_60 = stq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_60 = stq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_60 = stq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_60 = stq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_60 = stq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_60 = stq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_60 = stq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_60 = stq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_60 = stq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_60 = stq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_60 = stq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_60 = stq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_60 = stq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_60 = stq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_60 = stq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_60 = stq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_60 = stq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_60 = stq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_60 = stq_30_bits_uop_pdst;
      default:
        casez_tmp_60 = stq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_61 = stq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_61 = stq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_61 = stq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_61 = stq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_61 = stq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_61 = stq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_61 = stq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_61 = stq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_61 = stq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_61 = stq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_61 = stq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_61 = stq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_61 = stq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_61 = stq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_61 = stq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_61 = stq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_61 = stq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_61 = stq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_61 = stq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_61 = stq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_61 = stq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_61 = stq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_61 = stq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_61 = stq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_61 = stq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_61 = stq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_61 = stq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_61 = stq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_61 = stq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_61 = stq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_61 = stq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_61 = stq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_62 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_62 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_62 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_62 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_62 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_62 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_62 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_62 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_62 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_62 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_62 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_62 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_62 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_62 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_62 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_62 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_62 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_62 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_62 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_62 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_62 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_62 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_62 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_62 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_62 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_62 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_62 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_62 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_62 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_62 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_62 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_62 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_63 = stq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_63 = stq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_63 = stq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_63 = stq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_63 = stq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_63 = stq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_63 = stq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_63 = stq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_63 = stq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_63 = stq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_63 = stq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_63 = stq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_63 = stq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_63 = stq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_63 = stq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_63 = stq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_63 = stq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_63 = stq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_63 = stq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_63 = stq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_63 = stq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_63 = stq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_63 = stq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_63 = stq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_63 = stq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_63 = stq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_63 = stq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_63 = stq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_63 = stq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_63 = stq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_63 = stq_30_bits_uop_mem_signed;
      default:
        casez_tmp_63 = stq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_64 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_64 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_64 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_64 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_64 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_64 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_64 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_64 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_64 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_64 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_64 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_64 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_64 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_64 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_64 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_64 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_64 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_64 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_64 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_64 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_64 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_64 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_64 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_64 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_64 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_64 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_64 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_64 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_64 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_64 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_64 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_64 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_65 = stq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_65 = stq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_65 = stq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_65 = stq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_65 = stq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_65 = stq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_65 = stq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_65 = stq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_65 = stq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_65 = stq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_65 = stq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_65 = stq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_65 = stq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_65 = stq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_65 = stq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_65 = stq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_65 = stq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_65 = stq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_65 = stq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_65 = stq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_65 = stq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_65 = stq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_65 = stq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_65 = stq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_65 = stq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_65 = stq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_65 = stq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_65 = stq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_65 = stq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_65 = stq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_65 = stq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_65 = stq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_66 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_66 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_66 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_66 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_66 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_66 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_66 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_66 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_66 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_66 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_66 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_66 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_66 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_66 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_66 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_66 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_66 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_66 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_66 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_66 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_66 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_66 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_66 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_66 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_66 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_66 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_66 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_66 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_66 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_66 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_66 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_66 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_67 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_67 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_67 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_67 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_67 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_67 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_67 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_67 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_67 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_67 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_67 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_67 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_67 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_67 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_67 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_67 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_67 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_67 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_67 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_67 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_67 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_67 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_67 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_67 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_67 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_67 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_67 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_67 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_67 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_67 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_67 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_67 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_68 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_68 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_68 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_68 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_68 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_68 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_68 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_68 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_68 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_68 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_68 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_68 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_68 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_68 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_68 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_68 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_68 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_68 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_68 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_68 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_68 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_68 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_68 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_68 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_68 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_68 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_68 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_68 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_68 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_68 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_68 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_68 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_69 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_69 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_69 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_69 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_69 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_69 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_69 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_69 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_69 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_69 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_69 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_69 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_69 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_69 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_69 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_69 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_69 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_69 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_69 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_69 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_69 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_69 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_69 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_69 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_69 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_69 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_69 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_69 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_69 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_69 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_69 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_69 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_70 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_70 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_70 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_70 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_70 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_70 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_70 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_70 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_70 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_70 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_70 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_70 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_70 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_70 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_70 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_70 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_70 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_70 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_70 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_70 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_70 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_70 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_70 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_70 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_70 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_70 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_70 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_70 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_70 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_70 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_70 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_70 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_71 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_71 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_71 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_71 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_71 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_71 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_71 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_71 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_71 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_71 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_71 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_71 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_71 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_71 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_71 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_71 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_71 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_71 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_71 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_71 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_71 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_71 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_71 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_71 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_71 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_71 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_71 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_71 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_71 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_71 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_71 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_71 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_72 = ldq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_72 = ldq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_72 = ldq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_72 = ldq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_72 = ldq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_72 = ldq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_72 = ldq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_72 = ldq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_72 = ldq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_72 = ldq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_72 = ldq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_72 = ldq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_72 = ldq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_72 = ldq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_72 = ldq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_72 = ldq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_72 = ldq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_72 = ldq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_72 = ldq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_72 = ldq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_72 = ldq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_72 = ldq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_72 = ldq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_72 = ldq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_72 = ldq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_72 = ldq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_72 = ldq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_72 = ldq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_72 = ldq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_72 = ldq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_72 = ldq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_72 = ldq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_73 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_73 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_73 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_73 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_73 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_73 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_73 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_73 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_73 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_73 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_73 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_73 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_73 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_73 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_73 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_73 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_73 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_73 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_73 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_73 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_73 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_73 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_73 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_73 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_73 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_73 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_73 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_73 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_73 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_73 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_73 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_73 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_74 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_74 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_74 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_74 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_74 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_74 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_74 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_74 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_74 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_74 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_74 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_74 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_74 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_74 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_74 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_74 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_74 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_74 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_74 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_74 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_74 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_74 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_74 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_74 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_74 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_74 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_74 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_74 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_74 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_74 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_74 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_74 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_75 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_75 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_75 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_75 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_75 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_75 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_75 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_75 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_75 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_75 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_75 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_75 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_75 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_75 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_75 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_75 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_75 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_75 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_75 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_75 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_75 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_75 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_75 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_75 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_75 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_75 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_75 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_75 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_75 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_75 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_75 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_75 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_76 = ldq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_76 = ldq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_76 = ldq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_76 = ldq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_76 = ldq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_76 = ldq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_76 = ldq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_76 = ldq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_76 = ldq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_76 = ldq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_76 = ldq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_76 = ldq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_76 = ldq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_76 = ldq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_76 = ldq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_76 = ldq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_76 = ldq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_76 = ldq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_76 = ldq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_76 = ldq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_76 = ldq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_76 = ldq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_76 = ldq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_76 = ldq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_76 = ldq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_76 = ldq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_76 = ldq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_76 = ldq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_76 = ldq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_76 = ldq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_76 = ldq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_76 = ldq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_77 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_77 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_77 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_77 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_77 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_77 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_77 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_77 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_77 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_77 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_77 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_77 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_77 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_77 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_77 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_77 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_77 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_77 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_77 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_77 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_77 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_77 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_77 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_77 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_77 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_77 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_77 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_77 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_77 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_77 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_77 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_77 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  wire [19:0] exe_tlb_uop_0_br_mask = _exe_tlb_uop_T_2 ? exe_req_0_bits_uop_br_mask : 20'h0;
  wire        exe_tlb_uop_0_uses_ldq = _exe_tlb_uop_T_2 & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_uses_ldq : io_core_exe_0_req_bits_uop_uses_ldq);
  wire        exe_tlb_uop_0_uses_stq = _exe_tlb_uop_T_2 & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_uses_stq : io_core_exe_0_req_bits_uop_uses_stq);
  wire        _exe_tlb_uop_T_9 = _exe_cmd_T_7 | will_fire_sta_incoming_1 | will_fire_sfence_1;
  wire        _exe_tlb_uop_T_11_uses_ldq = will_fire_sta_retry_1 & casez_tmp_65;
  wire [19:0] exe_tlb_uop_1_br_mask = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_br_mask : will_fire_load_retry_1 ? casez_tmp_67 : will_fire_sta_retry_1 ? casez_tmp_56 : 20'h0;
  wire [4:0]  exe_tlb_uop_1_mem_cmd = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_mem_cmd : will_fire_load_retry_1 ? casez_tmp_72 : will_fire_sta_retry_1 ? casez_tmp_61 : 5'h0;
  wire [1:0]  exe_tlb_uop_1_mem_size = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_mem_size : will_fire_load_retry_1 ? casez_tmp_73 : will_fire_sta_retry_1 ? casez_tmp_62 : 2'h0;
  wire        exe_tlb_uop_1_uses_ldq = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_uses_ldq : will_fire_load_retry_1 ? casez_tmp_76 : _exe_tlb_uop_T_11_uses_ldq;
  wire        exe_tlb_uop_1_uses_stq = _exe_tlb_uop_T_9 ? exe_req_1_bits_uop_uses_stq : will_fire_load_retry_1 ? casez_tmp_77 : will_fire_sta_retry_1 & casez_tmp_66;
  wire        _exe_tlb_vaddr_T_1 = _exe_cmd_T | will_fire_sta_incoming_0;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_78 = stq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_78 = stq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_78 = stq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_78 = stq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_78 = stq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_78 = stq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_78 = stq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_78 = stq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_78 = stq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_78 = stq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_78 = stq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_78 = stq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_78 = stq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_78 = stq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_78 = stq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_78 = stq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_78 = stq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_78 = stq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_78 = stq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_78 = stq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_78 = stq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_78 = stq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_78 = stq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_78 = stq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_78 = stq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_78 = stq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_78 = stq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_78 = stq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_78 = stq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_78 = stq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_78 = stq_30_bits_addr_bits;
      default:
        casez_tmp_78 = stq_31_bits_addr_bits;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_79 = ldq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_79 = ldq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_79 = ldq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_79 = ldq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_79 = ldq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_79 = ldq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_79 = ldq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_79 = ldq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_79 = ldq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_79 = ldq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_79 = ldq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_79 = ldq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_79 = ldq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_79 = ldq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_79 = ldq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_79 = ldq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_79 = ldq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_79 = ldq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_79 = ldq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_79 = ldq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_79 = ldq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_79 = ldq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_79 = ldq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_79 = ldq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_79 = ldq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_79 = ldq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_79 = ldq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_79 = ldq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_79 = ldq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_79 = ldq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_79 = ldq_30_bits_addr_bits;
      default:
        casez_tmp_79 = ldq_31_bits_addr_bits;
    endcase
  end // always @(*)
  wire [39:0] _GEN_332 = {1'h0, exe_req_0_bits_sfence_bits_addr};
  wire [39:0] exe_tlb_vaddr_0 = _exe_tlb_vaddr_T_1 ? (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_addr : io_core_exe_0_req_bits_addr) : will_fire_sfence_0 ? _GEN_332 : 40'h0;
  wire        _exe_tlb_vaddr_T_8 = _exe_cmd_T_7 | will_fire_sta_incoming_1;
  wire [39:0] _GEN_333 = {1'h0, exe_req_1_bits_sfence_bits_addr};
  wire [39:0] exe_tlb_vaddr_1 = _exe_tlb_vaddr_T_8 ? (_GEN_329 ? io_core_exe_1_req_bits_addr : io_core_exe_0_req_bits_addr) : will_fire_sfence_1 ? _GEN_333 : will_fire_load_retry_1 ? casez_tmp_79 : will_fire_sta_retry_1 ? casez_tmp_78 : will_fire_hella_incoming_1 ? hella_req_addr : 40'h0;
  wire        _stq_idx_T = will_fire_sta_incoming_0 | will_fire_stad_incoming_0;
  wire        _stq_idx_T_1 = will_fire_sta_incoming_1 | will_fire_stad_incoming_1;
  reg  [19:0] mem_xcpt_uops_0_br_mask;
  reg  [6:0]  mem_xcpt_uops_0_rob_idx;
  reg  [4:0]  mem_xcpt_uops_0_stq_idx;
  reg         mem_xcpt_uops_0_uses_ldq;
  reg  [19:0] mem_xcpt_uops_1_br_mask;
  reg  [6:0]  mem_xcpt_uops_1_rob_idx;
  reg  [4:0]  mem_xcpt_uops_1_stq_idx;
  reg         mem_xcpt_uops_1_uses_ldq;
  reg  [3:0]  mem_xcpt_causes_0;
  reg  [3:0]  mem_xcpt_causes_1;
  reg  [39:0] mem_xcpt_vaddrs_0;
  reg  [39:0] mem_xcpt_vaddrs_1;
  wire        exe_tlb_miss_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_miss;
  wire        exe_tlb_miss_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_miss;
  wire [31:0] exe_tlb_paddr_0 = {_dtlb_io_resp_0_paddr[31:12], exe_tlb_vaddr_0[11:0]};
  wire [31:0] exe_tlb_paddr_1 = {_dtlb_io_resp_1_paddr[31:12], exe_tlb_vaddr_1[11:0]};
  wire        dmem_req_0_valid = can_fire_load_incoming_0 ? ~exe_tlb_miss_0 & _dtlb_io_resp_0_cacheable : will_fire_store_commit_0;
  wire        dmem_req_1_valid = can_fire_load_incoming_1 ? ~exe_tlb_miss_1 & _dtlb_io_resp_1_cacheable : will_fire_load_retry_1 ? ~exe_tlb_miss_1 & _dtlb_io_resp_1_cacheable : will_fire_load_wakeup_1 | (will_fire_hella_incoming_1 ? ~io_hellacache_s1_kill & (~exe_tlb_miss_1 | hella_req_phys) : will_fire_hella_wakeup_1);
  wire        _io_dmem_req_valid_output = dmem_req_0_valid | dmem_req_1_valid;
  wire        _dmem_req_fire_T_2 = io_dmem_req_ready & _io_dmem_req_valid_output;
  wire        dmem_req_fire_1 = dmem_req_1_valid & _dmem_req_fire_T_2;
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_80 = stq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_80 = stq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_80 = stq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_80 = stq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_80 = stq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_80 = stq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_80 = stq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_80 = stq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_80 = stq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_80 = stq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_80 = stq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_80 = stq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_80 = stq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_80 = stq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_80 = stq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_80 = stq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_80 = stq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_80 = stq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_80 = stq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_80 = stq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_80 = stq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_80 = stq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_80 = stq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_80 = stq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_80 = stq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_80 = stq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_80 = stq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_80 = stq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_80 = stq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_80 = stq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_80 = stq_30_bits_addr_bits;
      default:
        casez_tmp_80 = stq_31_bits_addr_bits;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_81 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_81 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_81 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_81 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_81 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_81 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_81 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_81 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_81 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_81 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_81 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_81 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_81 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_81 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_81 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_81 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_81 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_81 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_81 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_81 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_81 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_81 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_81 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_81 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_81 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_81 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_81 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_81 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_81 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_81 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_81 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_81 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_82 = stq_0_bits_data_bits;
      5'b00001:
        casez_tmp_82 = stq_1_bits_data_bits;
      5'b00010:
        casez_tmp_82 = stq_2_bits_data_bits;
      5'b00011:
        casez_tmp_82 = stq_3_bits_data_bits;
      5'b00100:
        casez_tmp_82 = stq_4_bits_data_bits;
      5'b00101:
        casez_tmp_82 = stq_5_bits_data_bits;
      5'b00110:
        casez_tmp_82 = stq_6_bits_data_bits;
      5'b00111:
        casez_tmp_82 = stq_7_bits_data_bits;
      5'b01000:
        casez_tmp_82 = stq_8_bits_data_bits;
      5'b01001:
        casez_tmp_82 = stq_9_bits_data_bits;
      5'b01010:
        casez_tmp_82 = stq_10_bits_data_bits;
      5'b01011:
        casez_tmp_82 = stq_11_bits_data_bits;
      5'b01100:
        casez_tmp_82 = stq_12_bits_data_bits;
      5'b01101:
        casez_tmp_82 = stq_13_bits_data_bits;
      5'b01110:
        casez_tmp_82 = stq_14_bits_data_bits;
      5'b01111:
        casez_tmp_82 = stq_15_bits_data_bits;
      5'b10000:
        casez_tmp_82 = stq_16_bits_data_bits;
      5'b10001:
        casez_tmp_82 = stq_17_bits_data_bits;
      5'b10010:
        casez_tmp_82 = stq_18_bits_data_bits;
      5'b10011:
        casez_tmp_82 = stq_19_bits_data_bits;
      5'b10100:
        casez_tmp_82 = stq_20_bits_data_bits;
      5'b10101:
        casez_tmp_82 = stq_21_bits_data_bits;
      5'b10110:
        casez_tmp_82 = stq_22_bits_data_bits;
      5'b10111:
        casez_tmp_82 = stq_23_bits_data_bits;
      5'b11000:
        casez_tmp_82 = stq_24_bits_data_bits;
      5'b11001:
        casez_tmp_82 = stq_25_bits_data_bits;
      5'b11010:
        casez_tmp_82 = stq_26_bits_data_bits;
      5'b11011:
        casez_tmp_82 = stq_27_bits_data_bits;
      5'b11100:
        casez_tmp_82 = stq_28_bits_data_bits;
      5'b11101:
        casez_tmp_82 = stq_29_bits_data_bits;
      5'b11110:
        casez_tmp_82 = stq_30_bits_data_bits;
      default:
        casez_tmp_82 = stq_31_bits_data_bits;
    endcase
  end // always @(*)
  always @(*) begin
    casez (casez_tmp_81)
      2'b00:
        casez_tmp_83 = {2{{2{{2{casez_tmp_82[7:0]}}}}}};
      2'b01:
        casez_tmp_83 = {2{{2{casez_tmp_82[15:0]}}}};
      2'b10:
        casez_tmp_83 = {2{casez_tmp_82[31:0]}};
      default:
        casez_tmp_83 = casez_tmp_82;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_84 = stq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_84 = stq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_84 = stq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_84 = stq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_84 = stq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_84 = stq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_84 = stq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_84 = stq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_84 = stq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_84 = stq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_84 = stq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_84 = stq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_84 = stq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_84 = stq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_84 = stq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_84 = stq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_84 = stq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_84 = stq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_84 = stq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_84 = stq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_84 = stq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_84 = stq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_84 = stq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_84 = stq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_84 = stq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_84 = stq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_84 = stq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_84 = stq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_84 = stq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_84 = stq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_84 = stq_30_bits_uop_br_mask;
      default:
        casez_tmp_84 = stq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_85 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_85 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_85 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_85 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_85 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_85 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_85 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_85 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_85 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_85 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_85 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_85 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_85 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_85 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_85 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_85 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_85 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_85 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_85 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_85 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_85 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_85 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_85 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_85 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_85 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_85 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_85 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_85 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_85 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_85 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_85 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_85 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_86 = stq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_86 = stq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_86 = stq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_86 = stq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_86 = stq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_86 = stq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_86 = stq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_86 = stq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_86 = stq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_86 = stq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_86 = stq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_86 = stq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_86 = stq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_86 = stq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_86 = stq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_86 = stq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_86 = stq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_86 = stq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_86 = stq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_86 = stq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_86 = stq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_86 = stq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_86 = stq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_86 = stq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_86 = stq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_86 = stq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_86 = stq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_86 = stq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_86 = stq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_86 = stq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_86 = stq_30_bits_uop_stq_idx;
      default:
        casez_tmp_86 = stq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_87 = stq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_87 = stq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_87 = stq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_87 = stq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_87 = stq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_87 = stq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_87 = stq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_87 = stq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_87 = stq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_87 = stq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_87 = stq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_87 = stq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_87 = stq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_87 = stq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_87 = stq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_87 = stq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_87 = stq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_87 = stq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_87 = stq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_87 = stq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_87 = stq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_87 = stq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_87 = stq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_87 = stq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_87 = stq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_87 = stq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_87 = stq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_87 = stq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_87 = stq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_87 = stq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_87 = stq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_87 = stq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_88 = stq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_88 = stq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_88 = stq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_88 = stq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_88 = stq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_88 = stq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_88 = stq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_88 = stq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_88 = stq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_88 = stq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_88 = stq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_88 = stq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_88 = stq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_88 = stq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_88 = stq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_88 = stq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_88 = stq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_88 = stq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_88 = stq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_88 = stq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_88 = stq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_88 = stq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_88 = stq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_88 = stq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_88 = stq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_88 = stq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_88 = stq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_88 = stq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_88 = stq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_88 = stq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_88 = stq_30_bits_uop_mem_signed;
      default:
        casez_tmp_88 = stq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_89 = stq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_89 = stq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_89 = stq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_89 = stq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_89 = stq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_89 = stq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_89 = stq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_89 = stq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_89 = stq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_89 = stq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_89 = stq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_89 = stq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_89 = stq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_89 = stq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_89 = stq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_89 = stq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_89 = stq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_89 = stq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_89 = stq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_89 = stq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_89 = stq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_89 = stq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_89 = stq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_89 = stq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_89 = stq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_89 = stq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_89 = stq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_89 = stq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_89 = stq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_89 = stq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_89 = stq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_89 = stq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (stq_execute_head)
      5'b00000:
        casez_tmp_90 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_90 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_90 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_90 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_90 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_90 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_90 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_90 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_90 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_90 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_90 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_90 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_90 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_90 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_90 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_90 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_90 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_90 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_90 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_90 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_90 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_90 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_90 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_90 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_90 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_90 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_90 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_90 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_90 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_90 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_90 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_90 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_91 = ldq_0_bits_addr_bits;
      5'b00001:
        casez_tmp_91 = ldq_1_bits_addr_bits;
      5'b00010:
        casez_tmp_91 = ldq_2_bits_addr_bits;
      5'b00011:
        casez_tmp_91 = ldq_3_bits_addr_bits;
      5'b00100:
        casez_tmp_91 = ldq_4_bits_addr_bits;
      5'b00101:
        casez_tmp_91 = ldq_5_bits_addr_bits;
      5'b00110:
        casez_tmp_91 = ldq_6_bits_addr_bits;
      5'b00111:
        casez_tmp_91 = ldq_7_bits_addr_bits;
      5'b01000:
        casez_tmp_91 = ldq_8_bits_addr_bits;
      5'b01001:
        casez_tmp_91 = ldq_9_bits_addr_bits;
      5'b01010:
        casez_tmp_91 = ldq_10_bits_addr_bits;
      5'b01011:
        casez_tmp_91 = ldq_11_bits_addr_bits;
      5'b01100:
        casez_tmp_91 = ldq_12_bits_addr_bits;
      5'b01101:
        casez_tmp_91 = ldq_13_bits_addr_bits;
      5'b01110:
        casez_tmp_91 = ldq_14_bits_addr_bits;
      5'b01111:
        casez_tmp_91 = ldq_15_bits_addr_bits;
      5'b10000:
        casez_tmp_91 = ldq_16_bits_addr_bits;
      5'b10001:
        casez_tmp_91 = ldq_17_bits_addr_bits;
      5'b10010:
        casez_tmp_91 = ldq_18_bits_addr_bits;
      5'b10011:
        casez_tmp_91 = ldq_19_bits_addr_bits;
      5'b10100:
        casez_tmp_91 = ldq_20_bits_addr_bits;
      5'b10101:
        casez_tmp_91 = ldq_21_bits_addr_bits;
      5'b10110:
        casez_tmp_91 = ldq_22_bits_addr_bits;
      5'b10111:
        casez_tmp_91 = ldq_23_bits_addr_bits;
      5'b11000:
        casez_tmp_91 = ldq_24_bits_addr_bits;
      5'b11001:
        casez_tmp_91 = ldq_25_bits_addr_bits;
      5'b11010:
        casez_tmp_91 = ldq_26_bits_addr_bits;
      5'b11011:
        casez_tmp_91 = ldq_27_bits_addr_bits;
      5'b11100:
        casez_tmp_91 = ldq_28_bits_addr_bits;
      5'b11101:
        casez_tmp_91 = ldq_29_bits_addr_bits;
      5'b11110:
        casez_tmp_91 = ldq_30_bits_addr_bits;
      default:
        casez_tmp_91 = ldq_31_bits_addr_bits;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_92 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_92 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_92 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_92 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_92 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_92 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_92 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_92 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_92 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_92 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_92 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_92 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_92 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_92 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_92 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_92 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_92 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_92 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_92 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_92 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_92 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_92 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_92 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_92 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_92 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_92 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_92 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_92 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_92 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_92 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_92 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_92 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_93 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_93 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_93 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_93 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_93 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_93 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_93 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_93 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_93 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_93 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_93 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_93 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_93 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_93 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_93 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_93 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_93 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_93 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_93 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_93 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_93 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_93 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_93 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_93 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_93 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_93 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_93 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_93 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_93 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_93 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_93 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_93 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_94 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_94 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_94 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_94 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_94 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_94 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_94 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_94 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_94 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_94 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_94 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_94 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_94 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_94 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_94 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_94 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_94 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_94 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_94 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_94 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_94 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_94 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_94 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_94 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_94 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_94 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_94 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_94 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_94 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_94 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_94 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_94 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_95 = ldq_0_bits_uop_mem_cmd;
      5'b00001:
        casez_tmp_95 = ldq_1_bits_uop_mem_cmd;
      5'b00010:
        casez_tmp_95 = ldq_2_bits_uop_mem_cmd;
      5'b00011:
        casez_tmp_95 = ldq_3_bits_uop_mem_cmd;
      5'b00100:
        casez_tmp_95 = ldq_4_bits_uop_mem_cmd;
      5'b00101:
        casez_tmp_95 = ldq_5_bits_uop_mem_cmd;
      5'b00110:
        casez_tmp_95 = ldq_6_bits_uop_mem_cmd;
      5'b00111:
        casez_tmp_95 = ldq_7_bits_uop_mem_cmd;
      5'b01000:
        casez_tmp_95 = ldq_8_bits_uop_mem_cmd;
      5'b01001:
        casez_tmp_95 = ldq_9_bits_uop_mem_cmd;
      5'b01010:
        casez_tmp_95 = ldq_10_bits_uop_mem_cmd;
      5'b01011:
        casez_tmp_95 = ldq_11_bits_uop_mem_cmd;
      5'b01100:
        casez_tmp_95 = ldq_12_bits_uop_mem_cmd;
      5'b01101:
        casez_tmp_95 = ldq_13_bits_uop_mem_cmd;
      5'b01110:
        casez_tmp_95 = ldq_14_bits_uop_mem_cmd;
      5'b01111:
        casez_tmp_95 = ldq_15_bits_uop_mem_cmd;
      5'b10000:
        casez_tmp_95 = ldq_16_bits_uop_mem_cmd;
      5'b10001:
        casez_tmp_95 = ldq_17_bits_uop_mem_cmd;
      5'b10010:
        casez_tmp_95 = ldq_18_bits_uop_mem_cmd;
      5'b10011:
        casez_tmp_95 = ldq_19_bits_uop_mem_cmd;
      5'b10100:
        casez_tmp_95 = ldq_20_bits_uop_mem_cmd;
      5'b10101:
        casez_tmp_95 = ldq_21_bits_uop_mem_cmd;
      5'b10110:
        casez_tmp_95 = ldq_22_bits_uop_mem_cmd;
      5'b10111:
        casez_tmp_95 = ldq_23_bits_uop_mem_cmd;
      5'b11000:
        casez_tmp_95 = ldq_24_bits_uop_mem_cmd;
      5'b11001:
        casez_tmp_95 = ldq_25_bits_uop_mem_cmd;
      5'b11010:
        casez_tmp_95 = ldq_26_bits_uop_mem_cmd;
      5'b11011:
        casez_tmp_95 = ldq_27_bits_uop_mem_cmd;
      5'b11100:
        casez_tmp_95 = ldq_28_bits_uop_mem_cmd;
      5'b11101:
        casez_tmp_95 = ldq_29_bits_uop_mem_cmd;
      5'b11110:
        casez_tmp_95 = ldq_30_bits_uop_mem_cmd;
      default:
        casez_tmp_95 = ldq_31_bits_uop_mem_cmd;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_96 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_96 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_96 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_96 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_96 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_96 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_96 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_96 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_96 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_96 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_96 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_96 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_96 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_96 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_96 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_96 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_96 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_96 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_96 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_96 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_96 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_96 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_96 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_96 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_96 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_96 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_96 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_96 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_96 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_96 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_96 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_96 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_97 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_97 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_97 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_97 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_97 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_97 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_97 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_97 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_97 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_97 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_97 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_97 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_97 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_97 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_97 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_97 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_97 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_97 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_97 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_97 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_97 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_97 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_97 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_97 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_97 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_97 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_97 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_97 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_97 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_97 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_97 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_97 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_98 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_98 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_98 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_98 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_98 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_98 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_98 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_98 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_98 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_98 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_98 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_98 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_98 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_98 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_98 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_98 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_98 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_98 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_98 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_98 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_98 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_98 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_98 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_98 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_98 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_98 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_98 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_98 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_98 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_98 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_98 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_98 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_99 = ldq_0_bits_uop_uses_ldq;
      5'b00001:
        casez_tmp_99 = ldq_1_bits_uop_uses_ldq;
      5'b00010:
        casez_tmp_99 = ldq_2_bits_uop_uses_ldq;
      5'b00011:
        casez_tmp_99 = ldq_3_bits_uop_uses_ldq;
      5'b00100:
        casez_tmp_99 = ldq_4_bits_uop_uses_ldq;
      5'b00101:
        casez_tmp_99 = ldq_5_bits_uop_uses_ldq;
      5'b00110:
        casez_tmp_99 = ldq_6_bits_uop_uses_ldq;
      5'b00111:
        casez_tmp_99 = ldq_7_bits_uop_uses_ldq;
      5'b01000:
        casez_tmp_99 = ldq_8_bits_uop_uses_ldq;
      5'b01001:
        casez_tmp_99 = ldq_9_bits_uop_uses_ldq;
      5'b01010:
        casez_tmp_99 = ldq_10_bits_uop_uses_ldq;
      5'b01011:
        casez_tmp_99 = ldq_11_bits_uop_uses_ldq;
      5'b01100:
        casez_tmp_99 = ldq_12_bits_uop_uses_ldq;
      5'b01101:
        casez_tmp_99 = ldq_13_bits_uop_uses_ldq;
      5'b01110:
        casez_tmp_99 = ldq_14_bits_uop_uses_ldq;
      5'b01111:
        casez_tmp_99 = ldq_15_bits_uop_uses_ldq;
      5'b10000:
        casez_tmp_99 = ldq_16_bits_uop_uses_ldq;
      5'b10001:
        casez_tmp_99 = ldq_17_bits_uop_uses_ldq;
      5'b10010:
        casez_tmp_99 = ldq_18_bits_uop_uses_ldq;
      5'b10011:
        casez_tmp_99 = ldq_19_bits_uop_uses_ldq;
      5'b10100:
        casez_tmp_99 = ldq_20_bits_uop_uses_ldq;
      5'b10101:
        casez_tmp_99 = ldq_21_bits_uop_uses_ldq;
      5'b10110:
        casez_tmp_99 = ldq_22_bits_uop_uses_ldq;
      5'b10111:
        casez_tmp_99 = ldq_23_bits_uop_uses_ldq;
      5'b11000:
        casez_tmp_99 = ldq_24_bits_uop_uses_ldq;
      5'b11001:
        casez_tmp_99 = ldq_25_bits_uop_uses_ldq;
      5'b11010:
        casez_tmp_99 = ldq_26_bits_uop_uses_ldq;
      5'b11011:
        casez_tmp_99 = ldq_27_bits_uop_uses_ldq;
      5'b11100:
        casez_tmp_99 = ldq_28_bits_uop_uses_ldq;
      5'b11101:
        casez_tmp_99 = ldq_29_bits_uop_uses_ldq;
      5'b11110:
        casez_tmp_99 = ldq_30_bits_uop_uses_ldq;
      default:
        casez_tmp_99 = ldq_31_bits_uop_uses_ldq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (ldq_wakeup_idx)
      5'b00000:
        casez_tmp_100 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_100 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_100 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_100 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_100 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_100 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_100 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_100 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_100 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_100 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_100 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_100 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_100 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_100 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_100 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_100 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_100 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_100 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_100 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_100 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_100 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_100 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_100 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_100 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_100 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_100 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_100 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_100 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_100 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_100 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_100 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_100 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  wire [39:0] _GEN_334 = {8'h0, _dtlb_io_resp_0_paddr[31:12], exe_tlb_vaddr_0[11:0]};
  wire        _io_core_fp_stdata_ready_output = ~will_fire_std_incoming_0 & ~will_fire_stad_incoming_0;
  wire        fp_stdata_fire = _io_core_fp_stdata_ready_output & io_core_fp_stdata_valid;
  wire        _stq_bits_data_bits_T = will_fire_std_incoming_0 | will_fire_stad_incoming_0;
  wire        _GEN_335 = _stq_bits_data_bits_T | fp_stdata_fire;
  wire [4:0]  sidx = _stq_bits_data_bits_T ? stq_incoming_idx_0 : io_core_fp_stdata_bits_uop_stq_idx;
  always @(*) begin
    casez (hella_req_size)
      2'b00:
        casez_tmp_101 = {2{{2{{2{hella_data_data[7:0]}}}}}};
      2'b01:
        casez_tmp_101 = {2{{2{hella_data_data[15:0]}}}};
      2'b10:
        casez_tmp_101 = {2{hella_data_data[31:0]}};
      default:
        casez_tmp_101 = hella_data_data;
    endcase
  end // always @(*)
  wire        _GEN_336 = will_fire_hella_incoming_1 | will_fire_hella_wakeup_1;
  wire [39:0] _GEN_337 = {8'h0, will_fire_hella_incoming_1 ? exe_tlb_paddr_1 : will_fire_hella_wakeup_1 ? hella_paddr : 32'h0};
  wire [39:0] _GEN_338 = {8'h0, _dtlb_io_resp_1_paddr[31:12], exe_tlb_vaddr_1[11:0]};
  wire        _GEN_339 = can_fire_load_incoming_1 | will_fire_load_retry_1;
  wire        _GEN_340 = can_fire_load_incoming_1 | will_fire_load_retry_1 | will_fire_load_wakeup_1;
  wire        _GEN_341 = can_fire_load_incoming_1 | will_fire_load_retry_1;
  wire        _GEN_342 = _stq_idx_T_1 | will_fire_sta_retry_1;
  wire        _stq_bits_data_bits_T_2 = will_fire_std_incoming_1 | will_fire_stad_incoming_1;
  wire [4:0]  sidx_1 = _stq_bits_data_bits_T_2 ? stq_incoming_idx_1 : io_core_fp_stdata_bits_uop_stq_idx;
  reg         fired_load_incoming_0;
  reg         fired_load_incoming_1;
  reg         fired_stad_incoming_0;
  reg         fired_stad_incoming_1;
  reg         fired_sta_incoming_0;
  reg         fired_sta_incoming_1;
  reg         fired_std_incoming_0;
  reg         fired_std_incoming_1;
  reg         fired_stdf_incoming;
  reg         fired_sfence_0;
  reg         fired_sfence_1;
  reg         fired_release_1;
  reg         fired_load_retry_1;
  reg         fired_sta_retry_1;
  reg         fired_load_wakeup_1;
  reg  [19:0] mem_incoming_uop_0_br_mask;
  reg  [6:0]  mem_incoming_uop_0_rob_idx;
  reg  [4:0]  mem_incoming_uop_0_ldq_idx;
  reg  [4:0]  mem_incoming_uop_0_stq_idx;
  reg  [6:0]  mem_incoming_uop_0_pdst;
  reg         mem_incoming_uop_0_fp_val;
  reg  [19:0] mem_incoming_uop_1_br_mask;
  reg  [6:0]  mem_incoming_uop_1_rob_idx;
  reg  [4:0]  mem_incoming_uop_1_ldq_idx;
  reg  [4:0]  mem_incoming_uop_1_stq_idx;
  reg  [6:0]  mem_incoming_uop_1_pdst;
  reg         mem_incoming_uop_1_fp_val;
  reg  [19:0] mem_ldq_incoming_e_0_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_incoming_e_0_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_incoming_e_0_bits_uop_mem_size;
  reg  [31:0] mem_ldq_incoming_e_0_bits_st_dep_mask;
  reg  [19:0] mem_ldq_incoming_e_1_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_incoming_e_1_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_incoming_e_1_bits_uop_mem_size;
  reg  [31:0] mem_ldq_incoming_e_1_bits_st_dep_mask;
  reg         mem_stq_incoming_e_0_valid;
  reg  [19:0] mem_stq_incoming_e_0_bits_uop_br_mask;
  reg  [6:0]  mem_stq_incoming_e_0_bits_uop_rob_idx;
  reg  [4:0]  mem_stq_incoming_e_0_bits_uop_stq_idx;
  reg  [1:0]  mem_stq_incoming_e_0_bits_uop_mem_size;
  reg         mem_stq_incoming_e_0_bits_uop_is_amo;
  reg         mem_stq_incoming_e_0_bits_addr_valid;
  reg         mem_stq_incoming_e_0_bits_addr_is_virtual;
  reg         mem_stq_incoming_e_0_bits_data_valid;
  reg         mem_stq_incoming_e_1_valid;
  reg  [19:0] mem_stq_incoming_e_1_bits_uop_br_mask;
  reg  [6:0]  mem_stq_incoming_e_1_bits_uop_rob_idx;
  reg  [4:0]  mem_stq_incoming_e_1_bits_uop_stq_idx;
  reg  [1:0]  mem_stq_incoming_e_1_bits_uop_mem_size;
  reg         mem_stq_incoming_e_1_bits_uop_is_amo;
  reg         mem_stq_incoming_e_1_bits_addr_valid;
  reg         mem_stq_incoming_e_1_bits_addr_is_virtual;
  reg         mem_stq_incoming_e_1_bits_data_valid;
  reg  [19:0] mem_ldq_wakeup_e_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_wakeup_e_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_wakeup_e_bits_uop_mem_size;
  reg  [31:0] mem_ldq_wakeup_e_bits_st_dep_mask;
  always @(*) begin
    casez (ldq_retry_idx)
      5'b00000:
        casez_tmp_102 = ldq_0_bits_st_dep_mask;
      5'b00001:
        casez_tmp_102 = ldq_1_bits_st_dep_mask;
      5'b00010:
        casez_tmp_102 = ldq_2_bits_st_dep_mask;
      5'b00011:
        casez_tmp_102 = ldq_3_bits_st_dep_mask;
      5'b00100:
        casez_tmp_102 = ldq_4_bits_st_dep_mask;
      5'b00101:
        casez_tmp_102 = ldq_5_bits_st_dep_mask;
      5'b00110:
        casez_tmp_102 = ldq_6_bits_st_dep_mask;
      5'b00111:
        casez_tmp_102 = ldq_7_bits_st_dep_mask;
      5'b01000:
        casez_tmp_102 = ldq_8_bits_st_dep_mask;
      5'b01001:
        casez_tmp_102 = ldq_9_bits_st_dep_mask;
      5'b01010:
        casez_tmp_102 = ldq_10_bits_st_dep_mask;
      5'b01011:
        casez_tmp_102 = ldq_11_bits_st_dep_mask;
      5'b01100:
        casez_tmp_102 = ldq_12_bits_st_dep_mask;
      5'b01101:
        casez_tmp_102 = ldq_13_bits_st_dep_mask;
      5'b01110:
        casez_tmp_102 = ldq_14_bits_st_dep_mask;
      5'b01111:
        casez_tmp_102 = ldq_15_bits_st_dep_mask;
      5'b10000:
        casez_tmp_102 = ldq_16_bits_st_dep_mask;
      5'b10001:
        casez_tmp_102 = ldq_17_bits_st_dep_mask;
      5'b10010:
        casez_tmp_102 = ldq_18_bits_st_dep_mask;
      5'b10011:
        casez_tmp_102 = ldq_19_bits_st_dep_mask;
      5'b10100:
        casez_tmp_102 = ldq_20_bits_st_dep_mask;
      5'b10101:
        casez_tmp_102 = ldq_21_bits_st_dep_mask;
      5'b10110:
        casez_tmp_102 = ldq_22_bits_st_dep_mask;
      5'b10111:
        casez_tmp_102 = ldq_23_bits_st_dep_mask;
      5'b11000:
        casez_tmp_102 = ldq_24_bits_st_dep_mask;
      5'b11001:
        casez_tmp_102 = ldq_25_bits_st_dep_mask;
      5'b11010:
        casez_tmp_102 = ldq_26_bits_st_dep_mask;
      5'b11011:
        casez_tmp_102 = ldq_27_bits_st_dep_mask;
      5'b11100:
        casez_tmp_102 = ldq_28_bits_st_dep_mask;
      5'b11101:
        casez_tmp_102 = ldq_29_bits_st_dep_mask;
      5'b11110:
        casez_tmp_102 = ldq_30_bits_st_dep_mask;
      default:
        casez_tmp_102 = ldq_31_bits_st_dep_mask;
    endcase
  end // always @(*)
  reg  [19:0] mem_ldq_retry_e_bits_uop_br_mask;
  reg  [4:0]  mem_ldq_retry_e_bits_uop_stq_idx;
  reg  [1:0]  mem_ldq_retry_e_bits_uop_mem_size;
  reg  [31:0] mem_ldq_retry_e_bits_st_dep_mask;
  always @(*) begin
    casez (stq_retry_idx)
      5'b00000:
        casez_tmp_103 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_103 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_103 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_103 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_103 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_103 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_103 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_103 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_103 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_103 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_103 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_103 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_103 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_103 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_103 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_103 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_103 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_103 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_103 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_103 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_103 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_103 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_103 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_103 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_103 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_103 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_103 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_103 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_103 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_103 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_103 = stq_30_bits_data_valid;
      default:
        casez_tmp_103 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  reg         mem_stq_retry_e_valid;
  reg  [19:0] mem_stq_retry_e_bits_uop_br_mask;
  reg  [6:0]  mem_stq_retry_e_bits_uop_rob_idx;
  reg  [4:0]  mem_stq_retry_e_bits_uop_stq_idx;
  reg  [1:0]  mem_stq_retry_e_bits_uop_mem_size;
  reg         mem_stq_retry_e_bits_uop_is_amo;
  reg         mem_stq_retry_e_bits_data_valid;
  wire [31:0] lcam_st_dep_mask_0 = fired_load_incoming_0 ? mem_ldq_incoming_e_0_bits_st_dep_mask : 32'h0;
  wire [31:0] lcam_st_dep_mask_1 = fired_load_incoming_1 ? mem_ldq_incoming_e_1_bits_st_dep_mask : fired_load_retry_1 ? mem_ldq_retry_e_bits_st_dep_mask : fired_load_wakeup_1 ? mem_ldq_wakeup_e_bits_st_dep_mask : 32'h0;
  wire        _lcam_stq_idx_T = fired_stad_incoming_0 | fired_sta_incoming_0;
  wire        _lcam_stq_idx_T_3 = fired_stad_incoming_1 | fired_sta_incoming_1;
  reg  [19:0] mem_stdf_uop_br_mask;
  reg  [6:0]  mem_stdf_uop_rob_idx;
  reg  [4:0]  mem_stdf_uop_stq_idx;
  reg         mem_tlb_miss_0;
  reg         mem_tlb_miss_1;
  reg         mem_tlb_uncacheable_0;
  reg         mem_tlb_uncacheable_1;
  reg  [39:0] mem_paddr_0;
  reg  [39:0] mem_paddr_1;
  reg         clr_bsy_valid_0;
  reg         clr_bsy_valid_1;
  reg  [6:0]  clr_bsy_rob_idx_0;
  reg  [6:0]  clr_bsy_rob_idx_1;
  reg  [19:0] clr_bsy_brmask_0;
  reg  [19:0] clr_bsy_brmask_1;
  reg         io_core_clr_bsy_0_valid_REG;
  reg         io_core_clr_bsy_0_valid_REG_1;
  reg         io_core_clr_bsy_0_valid_REG_2;
  reg         io_core_clr_bsy_1_valid_REG;
  reg         io_core_clr_bsy_1_valid_REG_1;
  reg         io_core_clr_bsy_1_valid_REG_2;
  reg         stdf_clr_bsy_valid;
  reg  [6:0]  stdf_clr_bsy_rob_idx;
  reg  [19:0] stdf_clr_bsy_brmask;
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_104 = stq_0_valid;
      5'b00001:
        casez_tmp_104 = stq_1_valid;
      5'b00010:
        casez_tmp_104 = stq_2_valid;
      5'b00011:
        casez_tmp_104 = stq_3_valid;
      5'b00100:
        casez_tmp_104 = stq_4_valid;
      5'b00101:
        casez_tmp_104 = stq_5_valid;
      5'b00110:
        casez_tmp_104 = stq_6_valid;
      5'b00111:
        casez_tmp_104 = stq_7_valid;
      5'b01000:
        casez_tmp_104 = stq_8_valid;
      5'b01001:
        casez_tmp_104 = stq_9_valid;
      5'b01010:
        casez_tmp_104 = stq_10_valid;
      5'b01011:
        casez_tmp_104 = stq_11_valid;
      5'b01100:
        casez_tmp_104 = stq_12_valid;
      5'b01101:
        casez_tmp_104 = stq_13_valid;
      5'b01110:
        casez_tmp_104 = stq_14_valid;
      5'b01111:
        casez_tmp_104 = stq_15_valid;
      5'b10000:
        casez_tmp_104 = stq_16_valid;
      5'b10001:
        casez_tmp_104 = stq_17_valid;
      5'b10010:
        casez_tmp_104 = stq_18_valid;
      5'b10011:
        casez_tmp_104 = stq_19_valid;
      5'b10100:
        casez_tmp_104 = stq_20_valid;
      5'b10101:
        casez_tmp_104 = stq_21_valid;
      5'b10110:
        casez_tmp_104 = stq_22_valid;
      5'b10111:
        casez_tmp_104 = stq_23_valid;
      5'b11000:
        casez_tmp_104 = stq_24_valid;
      5'b11001:
        casez_tmp_104 = stq_25_valid;
      5'b11010:
        casez_tmp_104 = stq_26_valid;
      5'b11011:
        casez_tmp_104 = stq_27_valid;
      5'b11100:
        casez_tmp_104 = stq_28_valid;
      5'b11101:
        casez_tmp_104 = stq_29_valid;
      5'b11110:
        casez_tmp_104 = stq_30_valid;
      default:
        casez_tmp_104 = stq_31_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_105 = stq_0_bits_addr_valid;
      5'b00001:
        casez_tmp_105 = stq_1_bits_addr_valid;
      5'b00010:
        casez_tmp_105 = stq_2_bits_addr_valid;
      5'b00011:
        casez_tmp_105 = stq_3_bits_addr_valid;
      5'b00100:
        casez_tmp_105 = stq_4_bits_addr_valid;
      5'b00101:
        casez_tmp_105 = stq_5_bits_addr_valid;
      5'b00110:
        casez_tmp_105 = stq_6_bits_addr_valid;
      5'b00111:
        casez_tmp_105 = stq_7_bits_addr_valid;
      5'b01000:
        casez_tmp_105 = stq_8_bits_addr_valid;
      5'b01001:
        casez_tmp_105 = stq_9_bits_addr_valid;
      5'b01010:
        casez_tmp_105 = stq_10_bits_addr_valid;
      5'b01011:
        casez_tmp_105 = stq_11_bits_addr_valid;
      5'b01100:
        casez_tmp_105 = stq_12_bits_addr_valid;
      5'b01101:
        casez_tmp_105 = stq_13_bits_addr_valid;
      5'b01110:
        casez_tmp_105 = stq_14_bits_addr_valid;
      5'b01111:
        casez_tmp_105 = stq_15_bits_addr_valid;
      5'b10000:
        casez_tmp_105 = stq_16_bits_addr_valid;
      5'b10001:
        casez_tmp_105 = stq_17_bits_addr_valid;
      5'b10010:
        casez_tmp_105 = stq_18_bits_addr_valid;
      5'b10011:
        casez_tmp_105 = stq_19_bits_addr_valid;
      5'b10100:
        casez_tmp_105 = stq_20_bits_addr_valid;
      5'b10101:
        casez_tmp_105 = stq_21_bits_addr_valid;
      5'b10110:
        casez_tmp_105 = stq_22_bits_addr_valid;
      5'b10111:
        casez_tmp_105 = stq_23_bits_addr_valid;
      5'b11000:
        casez_tmp_105 = stq_24_bits_addr_valid;
      5'b11001:
        casez_tmp_105 = stq_25_bits_addr_valid;
      5'b11010:
        casez_tmp_105 = stq_26_bits_addr_valid;
      5'b11011:
        casez_tmp_105 = stq_27_bits_addr_valid;
      5'b11100:
        casez_tmp_105 = stq_28_bits_addr_valid;
      5'b11101:
        casez_tmp_105 = stq_29_bits_addr_valid;
      5'b11110:
        casez_tmp_105 = stq_30_bits_addr_valid;
      default:
        casez_tmp_105 = stq_31_bits_addr_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_106 = stq_0_bits_addr_is_virtual;
      5'b00001:
        casez_tmp_106 = stq_1_bits_addr_is_virtual;
      5'b00010:
        casez_tmp_106 = stq_2_bits_addr_is_virtual;
      5'b00011:
        casez_tmp_106 = stq_3_bits_addr_is_virtual;
      5'b00100:
        casez_tmp_106 = stq_4_bits_addr_is_virtual;
      5'b00101:
        casez_tmp_106 = stq_5_bits_addr_is_virtual;
      5'b00110:
        casez_tmp_106 = stq_6_bits_addr_is_virtual;
      5'b00111:
        casez_tmp_106 = stq_7_bits_addr_is_virtual;
      5'b01000:
        casez_tmp_106 = stq_8_bits_addr_is_virtual;
      5'b01001:
        casez_tmp_106 = stq_9_bits_addr_is_virtual;
      5'b01010:
        casez_tmp_106 = stq_10_bits_addr_is_virtual;
      5'b01011:
        casez_tmp_106 = stq_11_bits_addr_is_virtual;
      5'b01100:
        casez_tmp_106 = stq_12_bits_addr_is_virtual;
      5'b01101:
        casez_tmp_106 = stq_13_bits_addr_is_virtual;
      5'b01110:
        casez_tmp_106 = stq_14_bits_addr_is_virtual;
      5'b01111:
        casez_tmp_106 = stq_15_bits_addr_is_virtual;
      5'b10000:
        casez_tmp_106 = stq_16_bits_addr_is_virtual;
      5'b10001:
        casez_tmp_106 = stq_17_bits_addr_is_virtual;
      5'b10010:
        casez_tmp_106 = stq_18_bits_addr_is_virtual;
      5'b10011:
        casez_tmp_106 = stq_19_bits_addr_is_virtual;
      5'b10100:
        casez_tmp_106 = stq_20_bits_addr_is_virtual;
      5'b10101:
        casez_tmp_106 = stq_21_bits_addr_is_virtual;
      5'b10110:
        casez_tmp_106 = stq_22_bits_addr_is_virtual;
      5'b10111:
        casez_tmp_106 = stq_23_bits_addr_is_virtual;
      5'b11000:
        casez_tmp_106 = stq_24_bits_addr_is_virtual;
      5'b11001:
        casez_tmp_106 = stq_25_bits_addr_is_virtual;
      5'b11010:
        casez_tmp_106 = stq_26_bits_addr_is_virtual;
      5'b11011:
        casez_tmp_106 = stq_27_bits_addr_is_virtual;
      5'b11100:
        casez_tmp_106 = stq_28_bits_addr_is_virtual;
      5'b11101:
        casez_tmp_106 = stq_29_bits_addr_is_virtual;
      5'b11110:
        casez_tmp_106 = stq_30_bits_addr_is_virtual;
      default:
        casez_tmp_106 = stq_31_bits_addr_is_virtual;
    endcase
  end // always @(*)
  always @(*) begin
    casez (mem_stdf_uop_stq_idx)
      5'b00000:
        casez_tmp_107 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_107 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_107 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_107 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_107 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_107 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_107 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_107 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_107 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_107 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_107 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_107 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_107 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_107 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_107 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_107 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_107 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_107 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_107 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_107 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_107 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_107 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_107 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_107 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_107 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_107 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_107 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_107 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_107 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_107 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_107 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_107 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  reg         io_core_clr_bsy_2_valid_REG;
  reg         io_core_clr_bsy_2_valid_REG_1;
  reg         io_core_clr_bsy_2_valid_REG_2;
  wire        do_st_search_0 = _lcam_stq_idx_T & ~mem_tlb_miss_0;
  wire        do_st_search_1 = (_lcam_stq_idx_T_3 | fired_sta_retry_1) & ~mem_tlb_miss_1;
  wire        _do_ld_search_T_2 = fired_load_incoming_0 & ~mem_tlb_miss_0;
  wire        _can_forward_T_6 = fired_load_incoming_1 | fired_load_retry_1;
  wire        do_ld_search_1 = _can_forward_T_6 & ~mem_tlb_miss_1 | fired_load_wakeup_1;
  reg  [31:0] lcam_addr_REG;
  wire [39:0] _GEN_343 = {8'h0, lcam_addr_REG};
  wire [39:0] lcam_addr_0 = _lcam_stq_idx_T ? _GEN_343 : mem_paddr_0;
  wire        _lcam_addr_T_5 = _lcam_stq_idx_T_3 | fired_sta_retry_1;
  reg  [31:0] lcam_addr_REG_2;
  reg  [31:0] lcam_addr_REG_3;
  wire [39:0] _GEN_344 = {8'h0, lcam_addr_REG_3};
  wire [39:0] _GEN_345 = {8'h0, lcam_addr_REG_2};
  wire [39:0] lcam_addr_1 = _lcam_addr_T_5 ? _GEN_345 : fired_release_1 ? _GEN_344 : mem_paddr_1;
  wire        _GEN_346 = _do_ld_search_T_2 & fired_load_incoming_0;
  wire [14:0] _lcam_mask_mask_T_2 = 15'h1 << lcam_addr_0[2:0];
  wire [14:0] _lcam_mask_mask_T_6 = 15'h3 << {12'h0, lcam_addr_0[2:1], 1'h0};
  always @(*) begin
    casez (do_st_search_0 ? (_lcam_stq_idx_T ? mem_stq_incoming_e_0_bits_uop_mem_size : 2'h0) : _GEN_346 ? mem_ldq_incoming_e_0_bits_uop_mem_size : 2'h0)
      2'b00:
        casez_tmp_108 = _lcam_mask_mask_T_2[7:0];
      2'b01:
        casez_tmp_108 = _lcam_mask_mask_T_6[7:0];
      2'b10:
        casez_tmp_108 = lcam_addr_0[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_108 = 8'hFF;
    endcase
  end // always @(*)
  wire [14:0] _lcam_mask_mask_T_17 = 15'h1 << lcam_addr_1[2:0];
  wire [14:0] _lcam_mask_mask_T_21 = 15'h3 << {12'h0, lcam_addr_1[2:1], 1'h0};
  always @(*) begin
    casez (do_st_search_1 ? (_lcam_stq_idx_T_3 ? mem_stq_incoming_e_1_bits_uop_mem_size : fired_sta_retry_1 ? mem_stq_retry_e_bits_uop_mem_size : 2'h0) : do_ld_search_1 ? (fired_load_incoming_1 ? mem_ldq_incoming_e_1_bits_uop_mem_size : fired_load_retry_1 ? mem_ldq_retry_e_bits_uop_mem_size : fired_load_wakeup_1 ? mem_ldq_wakeup_e_bits_uop_mem_size : 2'h0) : 2'h0)
      2'b00:
        casez_tmp_109 = _lcam_mask_mask_T_17[7:0];
      2'b01:
        casez_tmp_109 = _lcam_mask_mask_T_21[7:0];
      2'b10:
        casez_tmp_109 = lcam_addr_1[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_109 = 8'hFF;
    endcase
  end // always @(*)
  wire [4:0]  lcam_ldq_idx_0 = fired_load_incoming_0 ? mem_incoming_uop_0_ldq_idx : 5'h0;
  reg  [4:0]  lcam_ldq_idx_REG_2;
  reg  [4:0]  lcam_ldq_idx_REG_3;
  wire [4:0]  lcam_ldq_idx_1 = fired_load_incoming_1 ? mem_incoming_uop_1_ldq_idx : fired_load_wakeup_1 ? lcam_ldq_idx_REG_2 : fired_load_retry_1 ? lcam_ldq_idx_REG_3 : 5'h0;
  wire [4:0]  lcam_stq_idx_0 = _lcam_stq_idx_T ? mem_incoming_uop_0_stq_idx : 5'h0;
  reg  [4:0]  lcam_stq_idx_REG_1;
  wire [4:0]  lcam_stq_idx_1 = _lcam_stq_idx_T_3 ? mem_incoming_uop_1_stq_idx : fired_sta_retry_1 ? lcam_stq_idx_REG_1 : 5'h0;
  always @(*) begin
    casez (lcam_ldq_idx_0)
      5'b00000:
        casez_tmp_110 = ldq_0_bits_addr_is_uncacheable;
      5'b00001:
        casez_tmp_110 = ldq_1_bits_addr_is_uncacheable;
      5'b00010:
        casez_tmp_110 = ldq_2_bits_addr_is_uncacheable;
      5'b00011:
        casez_tmp_110 = ldq_3_bits_addr_is_uncacheable;
      5'b00100:
        casez_tmp_110 = ldq_4_bits_addr_is_uncacheable;
      5'b00101:
        casez_tmp_110 = ldq_5_bits_addr_is_uncacheable;
      5'b00110:
        casez_tmp_110 = ldq_6_bits_addr_is_uncacheable;
      5'b00111:
        casez_tmp_110 = ldq_7_bits_addr_is_uncacheable;
      5'b01000:
        casez_tmp_110 = ldq_8_bits_addr_is_uncacheable;
      5'b01001:
        casez_tmp_110 = ldq_9_bits_addr_is_uncacheable;
      5'b01010:
        casez_tmp_110 = ldq_10_bits_addr_is_uncacheable;
      5'b01011:
        casez_tmp_110 = ldq_11_bits_addr_is_uncacheable;
      5'b01100:
        casez_tmp_110 = ldq_12_bits_addr_is_uncacheable;
      5'b01101:
        casez_tmp_110 = ldq_13_bits_addr_is_uncacheable;
      5'b01110:
        casez_tmp_110 = ldq_14_bits_addr_is_uncacheable;
      5'b01111:
        casez_tmp_110 = ldq_15_bits_addr_is_uncacheable;
      5'b10000:
        casez_tmp_110 = ldq_16_bits_addr_is_uncacheable;
      5'b10001:
        casez_tmp_110 = ldq_17_bits_addr_is_uncacheable;
      5'b10010:
        casez_tmp_110 = ldq_18_bits_addr_is_uncacheable;
      5'b10011:
        casez_tmp_110 = ldq_19_bits_addr_is_uncacheable;
      5'b10100:
        casez_tmp_110 = ldq_20_bits_addr_is_uncacheable;
      5'b10101:
        casez_tmp_110 = ldq_21_bits_addr_is_uncacheable;
      5'b10110:
        casez_tmp_110 = ldq_22_bits_addr_is_uncacheable;
      5'b10111:
        casez_tmp_110 = ldq_23_bits_addr_is_uncacheable;
      5'b11000:
        casez_tmp_110 = ldq_24_bits_addr_is_uncacheable;
      5'b11001:
        casez_tmp_110 = ldq_25_bits_addr_is_uncacheable;
      5'b11010:
        casez_tmp_110 = ldq_26_bits_addr_is_uncacheable;
      5'b11011:
        casez_tmp_110 = ldq_27_bits_addr_is_uncacheable;
      5'b11100:
        casez_tmp_110 = ldq_28_bits_addr_is_uncacheable;
      5'b11101:
        casez_tmp_110 = ldq_29_bits_addr_is_uncacheable;
      5'b11110:
        casez_tmp_110 = ldq_30_bits_addr_is_uncacheable;
      default:
        casez_tmp_110 = ldq_31_bits_addr_is_uncacheable;
    endcase
  end // always @(*)
  always @(*) begin
    casez (lcam_ldq_idx_1)
      5'b00000:
        casez_tmp_111 = ldq_0_bits_addr_is_uncacheable;
      5'b00001:
        casez_tmp_111 = ldq_1_bits_addr_is_uncacheable;
      5'b00010:
        casez_tmp_111 = ldq_2_bits_addr_is_uncacheable;
      5'b00011:
        casez_tmp_111 = ldq_3_bits_addr_is_uncacheable;
      5'b00100:
        casez_tmp_111 = ldq_4_bits_addr_is_uncacheable;
      5'b00101:
        casez_tmp_111 = ldq_5_bits_addr_is_uncacheable;
      5'b00110:
        casez_tmp_111 = ldq_6_bits_addr_is_uncacheable;
      5'b00111:
        casez_tmp_111 = ldq_7_bits_addr_is_uncacheable;
      5'b01000:
        casez_tmp_111 = ldq_8_bits_addr_is_uncacheable;
      5'b01001:
        casez_tmp_111 = ldq_9_bits_addr_is_uncacheable;
      5'b01010:
        casez_tmp_111 = ldq_10_bits_addr_is_uncacheable;
      5'b01011:
        casez_tmp_111 = ldq_11_bits_addr_is_uncacheable;
      5'b01100:
        casez_tmp_111 = ldq_12_bits_addr_is_uncacheable;
      5'b01101:
        casez_tmp_111 = ldq_13_bits_addr_is_uncacheable;
      5'b01110:
        casez_tmp_111 = ldq_14_bits_addr_is_uncacheable;
      5'b01111:
        casez_tmp_111 = ldq_15_bits_addr_is_uncacheable;
      5'b10000:
        casez_tmp_111 = ldq_16_bits_addr_is_uncacheable;
      5'b10001:
        casez_tmp_111 = ldq_17_bits_addr_is_uncacheable;
      5'b10010:
        casez_tmp_111 = ldq_18_bits_addr_is_uncacheable;
      5'b10011:
        casez_tmp_111 = ldq_19_bits_addr_is_uncacheable;
      5'b10100:
        casez_tmp_111 = ldq_20_bits_addr_is_uncacheable;
      5'b10101:
        casez_tmp_111 = ldq_21_bits_addr_is_uncacheable;
      5'b10110:
        casez_tmp_111 = ldq_22_bits_addr_is_uncacheable;
      5'b10111:
        casez_tmp_111 = ldq_23_bits_addr_is_uncacheable;
      5'b11000:
        casez_tmp_111 = ldq_24_bits_addr_is_uncacheable;
      5'b11001:
        casez_tmp_111 = ldq_25_bits_addr_is_uncacheable;
      5'b11010:
        casez_tmp_111 = ldq_26_bits_addr_is_uncacheable;
      5'b11011:
        casez_tmp_111 = ldq_27_bits_addr_is_uncacheable;
      5'b11100:
        casez_tmp_111 = ldq_28_bits_addr_is_uncacheable;
      5'b11101:
        casez_tmp_111 = ldq_29_bits_addr_is_uncacheable;
      5'b11110:
        casez_tmp_111 = ldq_30_bits_addr_is_uncacheable;
      default:
        casez_tmp_111 = ldq_31_bits_addr_is_uncacheable;
    endcase
  end // always @(*)
  reg         s1_executing_loads_0;
  reg         s1_executing_loads_1;
  reg         s1_executing_loads_2;
  reg         s1_executing_loads_3;
  reg         s1_executing_loads_4;
  reg         s1_executing_loads_5;
  reg         s1_executing_loads_6;
  reg         s1_executing_loads_7;
  reg         s1_executing_loads_8;
  reg         s1_executing_loads_9;
  reg         s1_executing_loads_10;
  reg         s1_executing_loads_11;
  reg         s1_executing_loads_12;
  reg         s1_executing_loads_13;
  reg         s1_executing_loads_14;
  reg         s1_executing_loads_15;
  reg         s1_executing_loads_16;
  reg         s1_executing_loads_17;
  reg         s1_executing_loads_18;
  reg         s1_executing_loads_19;
  reg         s1_executing_loads_20;
  reg         s1_executing_loads_21;
  reg         s1_executing_loads_22;
  reg         s1_executing_loads_23;
  reg         s1_executing_loads_24;
  reg         s1_executing_loads_25;
  reg         s1_executing_loads_26;
  reg         s1_executing_loads_27;
  reg         s1_executing_loads_28;
  reg         s1_executing_loads_29;
  reg         s1_executing_loads_30;
  reg         s1_executing_loads_31;
  reg         wb_forward_valid_0;
  reg         wb_forward_valid_1;
  reg  [4:0]  wb_forward_ldq_idx_0;
  reg  [4:0]  wb_forward_ldq_idx_1;
  reg  [39:0] wb_forward_ld_addr_0;
  reg  [39:0] wb_forward_ld_addr_1;
  reg  [4:0]  wb_forward_stq_idx_0;
  reg  [4:0]  wb_forward_stq_idx_1;
  wire [14:0] _l_mask_mask_T_2 = 15'h1 << ldq_0_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_6 = 15'h3 << {12'h0, ldq_0_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_0_bits_uop_mem_size)
      2'b00:
        casez_tmp_112 = _l_mask_mask_T_2[7:0];
      2'b01:
        casez_tmp_112 = _l_mask_mask_T_6[7:0];
      2'b10:
        casez_tmp_112 = ldq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_112 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders__0 = wb_forward_valid_0 & ~(|wb_forward_ldq_idx_0);
  wire        l_forwarders__1 = wb_forward_valid_1 & ~(|wb_forward_ldq_idx_1);
  wire        l_is_forwarding = l_forwarders__0 | l_forwarders__1;
  wire [4:0]  l_forward_stq_idx = l_is_forwarding ? (l_forwarders__0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders__1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_0_bits_forward_stq_idx;
  wire        block_addr_matches__1 = lcam_addr_1[39:6] == ldq_0_bits_addr_bits[39:6];
  wire        dword_addr_matches__0 = lcam_addr_0[39:6] == ldq_0_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_0_bits_addr_bits[5:3];
  wire        dword_addr_matches__1 = block_addr_matches__1 & lcam_addr_1[5:3] == ldq_0_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T = casez_tmp_112 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_2 = casez_tmp_112 & casez_tmp_109;
  wire        _GEN_347 = ldq_0_bits_executed | ldq_0_bits_succeeded;
  wire        _GEN_348 = _GEN_347 | l_is_forwarding;
  wire [31:0] _GEN_349 = {27'h0, lcam_stq_idx_0};
  wire [31:0] _GEN_350 = ldq_0_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_351 = do_st_search_0 & ldq_0_valid & ldq_0_bits_addr_valid & _GEN_348 & ~ldq_0_bits_addr_is_virtual & _GEN_350[0] & dword_addr_matches__0 & (|_mask_overlap_T);
  wire        _forwarded_is_older_T_5 = l_forward_stq_idx < ldq_0_bits_youngest_stq_idx;
  wire        _GEN_83096 = ~ldq_0_bits_forward_std_val | l_forward_stq_idx != lcam_stq_idx_0 & (l_forward_stq_idx < lcam_stq_idx_0 ^ _forwarded_is_older_T_5 ^ lcam_stq_idx_0 < ldq_0_bits_youngest_stq_idx);
  wire        _GEN_352 = _do_ld_search_T_2 & ldq_0_valid & ldq_0_bits_addr_valid & ~ldq_0_bits_addr_is_virtual & dword_addr_matches__0 & (|_mask_overlap_T);
  wire        _searcher_is_older_T_249 = lcam_ldq_idx_0 < ldq_head;
  wire        searcher_is_older = _searcher_is_older_T_249 ^ (|ldq_head);
  wire        _GEN_353 = _GEN_348 & ~s1_executing_loads_0;
  wire        _GEN_83098 = _GEN_353 & ldq_0_bits_observed;
  reg         older_nacked_REG;
  wire        _GEN_116695 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h0;
  wire        _GEN_354 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h0;
  wire        nacking_loads_0 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_354 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116695;
  wire        _GEN_355 = ~_GEN_347 | nacking_loads_0 | older_nacked_REG;
  reg         io_dmem_s1_kill_0_REG;
  wire        _GEN_356 = (|lcam_ldq_idx_0) & _GEN_355;
  wire        _GEN_83272 = _GEN_351 ? _GEN_83096 : _GEN_352 & searcher_is_older & _GEN_83098;
  wire        _GEN_357 = fired_release_1 & ldq_0_valid & ldq_0_bits_addr_valid & block_addr_matches__1;
  wire [31:0] _GEN_358 = {27'h0, lcam_stq_idx_1};
  wire [31:0] _GEN_359 = ldq_0_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_360 = do_st_search_1 & ldq_0_valid & ldq_0_bits_addr_valid & _GEN_348 & ~ldq_0_bits_addr_is_virtual & _GEN_359[0] & dword_addr_matches__1 & (|_mask_overlap_T_2);
  wire        _GEN_361 = ~ldq_0_bits_forward_std_val | l_forward_stq_idx != lcam_stq_idx_1 & (l_forward_stq_idx < lcam_stq_idx_1 ^ _forwarded_is_older_T_5 ^ lcam_stq_idx_1 < ldq_0_bits_youngest_stq_idx);
  wire        _GEN_362 = do_ld_search_1 & ldq_0_valid & ldq_0_bits_addr_valid & ~ldq_0_bits_addr_is_virtual & dword_addr_matches__1 & (|_mask_overlap_T_2);
  wire        _searcher_is_older_T_253 = lcam_ldq_idx_1 < ldq_head;
  wire        searcher_is_older_1 = _searcher_is_older_T_253 ^ (|ldq_head);
  reg         older_nacked_REG_1;
  wire        _GEN_363 = ~_GEN_347 | nacking_loads_0 | older_nacked_REG_1;
  reg         io_dmem_s1_kill_1_REG;
  wire        _GEN_364 = (|lcam_ldq_idx_1) & _GEN_363;
  wire        _GEN_365 = _GEN_362 & searcher_is_older_1 & _GEN_353 & ldq_0_bits_observed;
  wire        failed_loads_0 = _GEN_357 ? _GEN_83272 : _GEN_360 ? _GEN_361 | _GEN_83272 : _GEN_365 | _GEN_83272;
  wire        _GEN_366 = _GEN_357 | _GEN_360;
  wire [14:0] _l_mask_mask_T_17 = 15'h1 << ldq_1_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_21 = 15'h3 << {12'h0, ldq_1_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_1_bits_uop_mem_size)
      2'b00:
        casez_tmp_113 = _l_mask_mask_T_17[7:0];
      2'b01:
        casez_tmp_113 = _l_mask_mask_T_21[7:0];
      2'b10:
        casez_tmp_113 = ldq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_113 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_1_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1;
  wire        l_forwarders_1_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1;
  wire        l_is_forwarding_1 = l_forwarders_1_0 | l_forwarders_1_1;
  wire [4:0]  l_forward_stq_idx_1 = l_is_forwarding_1 ? (l_forwarders_1_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_1_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_1_bits_forward_stq_idx;
  wire        block_addr_matches_1_1 = lcam_addr_1[39:6] == ldq_1_bits_addr_bits[39:6];
  wire        dword_addr_matches_1_0 = lcam_addr_0[39:6] == ldq_1_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_1_bits_addr_bits[5:3];
  wire        dword_addr_matches_1_1 = block_addr_matches_1_1 & lcam_addr_1[5:3] == ldq_1_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_4 = casez_tmp_113 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_6 = casez_tmp_113 & casez_tmp_109;
  wire        _GEN_367 = ldq_1_bits_executed | ldq_1_bits_succeeded;
  wire        _GEN_368 = _GEN_367 | l_is_forwarding_1;
  wire [31:0] _GEN_369 = ldq_1_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_370 = do_st_search_0 & ldq_1_valid & ldq_1_bits_addr_valid & _GEN_368 & ~ldq_1_bits_addr_is_virtual & _GEN_369[0] & dword_addr_matches_1_0 & (|_mask_overlap_T_4);
  wire        _forwarded_is_older_T_13 = l_forward_stq_idx_1 < ldq_1_bits_youngest_stq_idx;
  wire        _GEN_83594 = ~ldq_1_bits_forward_std_val | l_forward_stq_idx_1 != lcam_stq_idx_0 & (l_forward_stq_idx_1 < lcam_stq_idx_0 ^ _forwarded_is_older_T_13 ^ lcam_stq_idx_0 < ldq_1_bits_youngest_stq_idx);
  wire        _GEN_371 = _do_ld_search_T_2 & ldq_1_valid & ldq_1_bits_addr_valid & ~ldq_1_bits_addr_is_virtual & dword_addr_matches_1_0 & (|_mask_overlap_T_4);
  wire        searcher_is_older_2 = lcam_ldq_idx_0 == 5'h0 ^ _searcher_is_older_T_249 ^ (|(ldq_head[4:1]));
  wire        _GEN_372 = _GEN_368 & ~s1_executing_loads_1;
  wire        _GEN_83596 = _GEN_372 & ldq_1_bits_observed;
  wire        _GEN_373 = lcam_ldq_idx_0 != 5'h1;
  reg         older_nacked_REG_2;
  wire        _GEN_116696 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1;
  wire        _GEN_374 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1;
  wire        nacking_loads_1 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_374 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116696;
  wire        _GEN_375 = ~_GEN_367 | nacking_loads_1 | older_nacked_REG_2;
  reg         io_dmem_s1_kill_0_REG_1;
  wire        _GEN_83770 = _GEN_370 ? _GEN_83594 : _GEN_371 & searcher_is_older_2 & _GEN_83596;
  wire        _GEN_376 = _GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375);
  wire        _GEN_377 = fired_release_1 & ldq_1_valid & ldq_1_bits_addr_valid & block_addr_matches_1_1;
  wire [31:0] _GEN_378 = ldq_1_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_379 = do_st_search_1 & ldq_1_valid & ldq_1_bits_addr_valid & _GEN_368 & ~ldq_1_bits_addr_is_virtual & _GEN_378[0] & dword_addr_matches_1_1 & (|_mask_overlap_T_6);
  wire        _GEN_380 = ~ldq_1_bits_forward_std_val | l_forward_stq_idx_1 != lcam_stq_idx_1 & (l_forward_stq_idx_1 < lcam_stq_idx_1 ^ _forwarded_is_older_T_13 ^ lcam_stq_idx_1 < ldq_1_bits_youngest_stq_idx);
  wire        _GEN_381 = do_ld_search_1 & ldq_1_valid & ldq_1_bits_addr_valid & ~ldq_1_bits_addr_is_virtual & dword_addr_matches_1_1 & (|_mask_overlap_T_6);
  wire        searcher_is_older_3 = lcam_ldq_idx_1 == 5'h0 ^ _searcher_is_older_T_253 ^ (|(ldq_head[4:1]));
  wire        _GEN_382 = lcam_ldq_idx_1 != 5'h1;
  reg         older_nacked_REG_3;
  wire        _GEN_383 = ~_GEN_367 | nacking_loads_1 | older_nacked_REG_3;
  reg         io_dmem_s1_kill_1_REG_1;
  wire        _GEN_384 = _GEN_381 & searcher_is_older_3 & _GEN_372 & ldq_1_bits_observed;
  wire        failed_loads_1 = _GEN_377 ? _GEN_83770 : _GEN_379 ? _GEN_380 | _GEN_83770 : _GEN_384 | _GEN_83770;
  wire        _GEN_385 = _GEN_377 | _GEN_379;
  wire        _GEN_386 = _GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383);
  wire [14:0] _l_mask_mask_T_32 = 15'h1 << ldq_2_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_36 = 15'h3 << {12'h0, ldq_2_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_2_bits_uop_mem_size)
      2'b00:
        casez_tmp_114 = _l_mask_mask_T_32[7:0];
      2'b01:
        casez_tmp_114 = _l_mask_mask_T_36[7:0];
      2'b10:
        casez_tmp_114 = ldq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_114 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_2_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h2;
  wire        l_forwarders_2_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h2;
  wire        l_is_forwarding_2 = l_forwarders_2_0 | l_forwarders_2_1;
  wire [4:0]  l_forward_stq_idx_2 = l_is_forwarding_2 ? (l_forwarders_2_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_2_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_2_bits_forward_stq_idx;
  wire        block_addr_matches_2_1 = lcam_addr_1[39:6] == ldq_2_bits_addr_bits[39:6];
  wire        dword_addr_matches_2_0 = lcam_addr_0[39:6] == ldq_2_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_2_bits_addr_bits[5:3];
  wire        dword_addr_matches_2_1 = block_addr_matches_2_1 & lcam_addr_1[5:3] == ldq_2_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_8 = casez_tmp_114 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_10 = casez_tmp_114 & casez_tmp_109;
  wire        _GEN_387 = ldq_2_bits_executed | ldq_2_bits_succeeded;
  wire        _GEN_388 = _GEN_387 | l_is_forwarding_2;
  wire [31:0] _GEN_389 = ldq_2_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_390 = do_st_search_0 & ldq_2_valid & ldq_2_bits_addr_valid & _GEN_388 & ~ldq_2_bits_addr_is_virtual & _GEN_389[0] & dword_addr_matches_2_0 & (|_mask_overlap_T_8);
  wire        _forwarded_is_older_T_21 = l_forward_stq_idx_2 < ldq_2_bits_youngest_stq_idx;
  wire        _GEN_84092 = ~ldq_2_bits_forward_std_val | l_forward_stq_idx_2 != lcam_stq_idx_0 & (l_forward_stq_idx_2 < lcam_stq_idx_0 ^ _forwarded_is_older_T_21 ^ lcam_stq_idx_0 < ldq_2_bits_youngest_stq_idx);
  wire        _GEN_391 = _do_ld_search_T_2 & ldq_2_valid & ldq_2_bits_addr_valid & ~ldq_2_bits_addr_is_virtual & dword_addr_matches_2_0 & (|_mask_overlap_T_8);
  wire        _searcher_is_older_T_23 = ldq_head > 5'h2;
  wire        searcher_is_older_4 = lcam_ldq_idx_0 < 5'h2 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_23;
  wire        _GEN_392 = _GEN_388 & ~s1_executing_loads_2;
  wire        _GEN_84094 = _GEN_392 & ldq_2_bits_observed;
  wire        _GEN_393 = lcam_ldq_idx_0 != 5'h2;
  reg         older_nacked_REG_4;
  wire        _GEN_116697 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h2;
  wire        _GEN_394 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h2;
  wire        nacking_loads_2 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_394 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116697;
  wire        _GEN_395 = ~_GEN_387 | nacking_loads_2 | older_nacked_REG_4;
  reg         io_dmem_s1_kill_0_REG_2;
  wire        _GEN_84268 = _GEN_390 ? _GEN_84092 : _GEN_391 & searcher_is_older_4 & _GEN_84094;
  wire        _GEN_396 = _GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395);
  wire        _GEN_397 = fired_release_1 & ldq_2_valid & ldq_2_bits_addr_valid & block_addr_matches_2_1;
  wire [31:0] _GEN_398 = ldq_2_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_399 = do_st_search_1 & ldq_2_valid & ldq_2_bits_addr_valid & _GEN_388 & ~ldq_2_bits_addr_is_virtual & _GEN_398[0] & dword_addr_matches_2_1 & (|_mask_overlap_T_10);
  wire        _GEN_400 = ~ldq_2_bits_forward_std_val | l_forward_stq_idx_2 != lcam_stq_idx_1 & (l_forward_stq_idx_2 < lcam_stq_idx_1 ^ _forwarded_is_older_T_21 ^ lcam_stq_idx_1 < ldq_2_bits_youngest_stq_idx);
  wire        _GEN_401 = do_ld_search_1 & ldq_2_valid & ldq_2_bits_addr_valid & ~ldq_2_bits_addr_is_virtual & dword_addr_matches_2_1 & (|_mask_overlap_T_10);
  wire        searcher_is_older_5 = lcam_ldq_idx_1 < 5'h2 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_23;
  wire        _GEN_402 = lcam_ldq_idx_1 != 5'h2;
  reg         older_nacked_REG_5;
  wire        _GEN_403 = ~_GEN_387 | nacking_loads_2 | older_nacked_REG_5;
  reg         io_dmem_s1_kill_1_REG_2;
  wire        _GEN_404 = _GEN_401 & searcher_is_older_5 & _GEN_392 & ldq_2_bits_observed;
  wire        failed_loads_2 = _GEN_397 ? _GEN_84268 : _GEN_399 ? _GEN_400 | _GEN_84268 : _GEN_404 | _GEN_84268;
  wire        _GEN_405 = _GEN_397 | _GEN_399;
  wire        _GEN_406 = _GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403);
  wire [14:0] _l_mask_mask_T_47 = 15'h1 << ldq_3_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_51 = 15'h3 << {12'h0, ldq_3_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_3_bits_uop_mem_size)
      2'b00:
        casez_tmp_115 = _l_mask_mask_T_47[7:0];
      2'b01:
        casez_tmp_115 = _l_mask_mask_T_51[7:0];
      2'b10:
        casez_tmp_115 = ldq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_115 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_3_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h3;
  wire        l_forwarders_3_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h3;
  wire        l_is_forwarding_3 = l_forwarders_3_0 | l_forwarders_3_1;
  wire [4:0]  l_forward_stq_idx_3 = l_is_forwarding_3 ? (l_forwarders_3_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_3_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_3_bits_forward_stq_idx;
  wire        block_addr_matches_3_1 = lcam_addr_1[39:6] == ldq_3_bits_addr_bits[39:6];
  wire        dword_addr_matches_3_0 = lcam_addr_0[39:6] == ldq_3_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_3_bits_addr_bits[5:3];
  wire        dword_addr_matches_3_1 = block_addr_matches_3_1 & lcam_addr_1[5:3] == ldq_3_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_12 = casez_tmp_115 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_14 = casez_tmp_115 & casez_tmp_109;
  wire        _GEN_407 = ldq_3_bits_executed | ldq_3_bits_succeeded;
  wire        _GEN_408 = _GEN_407 | l_is_forwarding_3;
  wire [31:0] _GEN_409 = ldq_3_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_410 = do_st_search_0 & ldq_3_valid & ldq_3_bits_addr_valid & _GEN_408 & ~ldq_3_bits_addr_is_virtual & _GEN_409[0] & dword_addr_matches_3_0 & (|_mask_overlap_T_12);
  wire        _forwarded_is_older_T_29 = l_forward_stq_idx_3 < ldq_3_bits_youngest_stq_idx;
  wire        _GEN_84590 = ~ldq_3_bits_forward_std_val | l_forward_stq_idx_3 != lcam_stq_idx_0 & (l_forward_stq_idx_3 < lcam_stq_idx_0 ^ _forwarded_is_older_T_29 ^ lcam_stq_idx_0 < ldq_3_bits_youngest_stq_idx);
  wire        _GEN_411 = _do_ld_search_T_2 & ldq_3_valid & ldq_3_bits_addr_valid & ~ldq_3_bits_addr_is_virtual & dword_addr_matches_3_0 & (|_mask_overlap_T_12);
  wire        searcher_is_older_6 = lcam_ldq_idx_0 < 5'h3 ^ _searcher_is_older_T_249 ^ (|(ldq_head[4:2]));
  wire        _GEN_412 = _GEN_408 & ~s1_executing_loads_3;
  wire        _GEN_84592 = _GEN_412 & ldq_3_bits_observed;
  wire        _GEN_413 = lcam_ldq_idx_0 != 5'h3;
  reg         older_nacked_REG_6;
  wire        _GEN_116698 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h3;
  wire        _GEN_414 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h3;
  wire        nacking_loads_3 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_414 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116698;
  wire        _GEN_415 = ~_GEN_407 | nacking_loads_3 | older_nacked_REG_6;
  reg         io_dmem_s1_kill_0_REG_3;
  wire        _GEN_84766 = _GEN_410 ? _GEN_84590 : _GEN_411 & searcher_is_older_6 & _GEN_84592;
  wire        _GEN_416 = _GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415);
  wire        _GEN_417 = fired_release_1 & ldq_3_valid & ldq_3_bits_addr_valid & block_addr_matches_3_1;
  wire [31:0] _GEN_418 = ldq_3_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_419 = do_st_search_1 & ldq_3_valid & ldq_3_bits_addr_valid & _GEN_408 & ~ldq_3_bits_addr_is_virtual & _GEN_418[0] & dword_addr_matches_3_1 & (|_mask_overlap_T_14);
  wire        _GEN_420 = ~ldq_3_bits_forward_std_val | l_forward_stq_idx_3 != lcam_stq_idx_1 & (l_forward_stq_idx_3 < lcam_stq_idx_1 ^ _forwarded_is_older_T_29 ^ lcam_stq_idx_1 < ldq_3_bits_youngest_stq_idx);
  wire        _GEN_421 = do_ld_search_1 & ldq_3_valid & ldq_3_bits_addr_valid & ~ldq_3_bits_addr_is_virtual & dword_addr_matches_3_1 & (|_mask_overlap_T_14);
  wire        searcher_is_older_7 = lcam_ldq_idx_1 < 5'h3 ^ _searcher_is_older_T_253 ^ (|(ldq_head[4:2]));
  wire        _GEN_422 = lcam_ldq_idx_1 != 5'h3;
  reg         older_nacked_REG_7;
  wire        _GEN_423 = ~_GEN_407 | nacking_loads_3 | older_nacked_REG_7;
  reg         io_dmem_s1_kill_1_REG_3;
  wire        _GEN_424 = _GEN_421 & searcher_is_older_7 & _GEN_412 & ldq_3_bits_observed;
  wire        failed_loads_3 = _GEN_417 ? _GEN_84766 : _GEN_419 ? _GEN_420 | _GEN_84766 : _GEN_424 | _GEN_84766;
  wire        _GEN_425 = _GEN_417 | _GEN_419;
  wire        _GEN_426 = _GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423);
  wire [14:0] _l_mask_mask_T_62 = 15'h1 << ldq_4_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_66 = 15'h3 << {12'h0, ldq_4_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_4_bits_uop_mem_size)
      2'b00:
        casez_tmp_116 = _l_mask_mask_T_62[7:0];
      2'b01:
        casez_tmp_116 = _l_mask_mask_T_66[7:0];
      2'b10:
        casez_tmp_116 = ldq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_116 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_4_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h4;
  wire        l_forwarders_4_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h4;
  wire        l_is_forwarding_4 = l_forwarders_4_0 | l_forwarders_4_1;
  wire [4:0]  l_forward_stq_idx_4 = l_is_forwarding_4 ? (l_forwarders_4_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_4_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_4_bits_forward_stq_idx;
  wire        block_addr_matches_4_1 = lcam_addr_1[39:6] == ldq_4_bits_addr_bits[39:6];
  wire        dword_addr_matches_4_0 = lcam_addr_0[39:6] == ldq_4_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_4_bits_addr_bits[5:3];
  wire        dword_addr_matches_4_1 = block_addr_matches_4_1 & lcam_addr_1[5:3] == ldq_4_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_16 = casez_tmp_116 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_18 = casez_tmp_116 & casez_tmp_109;
  wire        _GEN_427 = ldq_4_bits_executed | ldq_4_bits_succeeded;
  wire        _GEN_428 = _GEN_427 | l_is_forwarding_4;
  wire [31:0] _GEN_429 = ldq_4_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_430 = do_st_search_0 & ldq_4_valid & ldq_4_bits_addr_valid & _GEN_428 & ~ldq_4_bits_addr_is_virtual & _GEN_429[0] & dword_addr_matches_4_0 & (|_mask_overlap_T_16);
  wire        _forwarded_is_older_T_37 = l_forward_stq_idx_4 < ldq_4_bits_youngest_stq_idx;
  wire        _GEN_85088 = ~ldq_4_bits_forward_std_val | l_forward_stq_idx_4 != lcam_stq_idx_0 & (l_forward_stq_idx_4 < lcam_stq_idx_0 ^ _forwarded_is_older_T_37 ^ lcam_stq_idx_0 < ldq_4_bits_youngest_stq_idx);
  wire        _GEN_431 = _do_ld_search_T_2 & ldq_4_valid & ldq_4_bits_addr_valid & ~ldq_4_bits_addr_is_virtual & dword_addr_matches_4_0 & (|_mask_overlap_T_16);
  wire        _searcher_is_older_T_39 = ldq_head > 5'h4;
  wire        searcher_is_older_8 = lcam_ldq_idx_0 < 5'h4 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_39;
  wire        _GEN_432 = _GEN_428 & ~s1_executing_loads_4;
  wire        _GEN_85090 = _GEN_432 & ldq_4_bits_observed;
  wire        _GEN_433 = lcam_ldq_idx_0 != 5'h4;
  reg         older_nacked_REG_8;
  wire        _GEN_116699 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h4;
  wire        _GEN_434 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h4;
  wire        nacking_loads_4 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_434 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116699;
  wire        _GEN_435 = ~_GEN_427 | nacking_loads_4 | older_nacked_REG_8;
  reg         io_dmem_s1_kill_0_REG_4;
  wire        _GEN_85264 = _GEN_430 ? _GEN_85088 : _GEN_431 & searcher_is_older_8 & _GEN_85090;
  wire        _GEN_436 = _GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435);
  wire        _GEN_437 = fired_release_1 & ldq_4_valid & ldq_4_bits_addr_valid & block_addr_matches_4_1;
  wire [31:0] _GEN_438 = ldq_4_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_439 = do_st_search_1 & ldq_4_valid & ldq_4_bits_addr_valid & _GEN_428 & ~ldq_4_bits_addr_is_virtual & _GEN_438[0] & dword_addr_matches_4_1 & (|_mask_overlap_T_18);
  wire        _GEN_440 = ~ldq_4_bits_forward_std_val | l_forward_stq_idx_4 != lcam_stq_idx_1 & (l_forward_stq_idx_4 < lcam_stq_idx_1 ^ _forwarded_is_older_T_37 ^ lcam_stq_idx_1 < ldq_4_bits_youngest_stq_idx);
  wire        _GEN_441 = do_ld_search_1 & ldq_4_valid & ldq_4_bits_addr_valid & ~ldq_4_bits_addr_is_virtual & dword_addr_matches_4_1 & (|_mask_overlap_T_18);
  wire        searcher_is_older_9 = lcam_ldq_idx_1 < 5'h4 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_39;
  wire        _GEN_442 = lcam_ldq_idx_1 != 5'h4;
  reg         older_nacked_REG_9;
  wire        _GEN_443 = ~_GEN_427 | nacking_loads_4 | older_nacked_REG_9;
  reg         io_dmem_s1_kill_1_REG_4;
  wire        _GEN_444 = _GEN_441 & searcher_is_older_9 & _GEN_432 & ldq_4_bits_observed;
  wire        failed_loads_4 = _GEN_437 ? _GEN_85264 : _GEN_439 ? _GEN_440 | _GEN_85264 : _GEN_444 | _GEN_85264;
  wire        _GEN_445 = _GEN_437 | _GEN_439;
  wire        _GEN_446 = _GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443);
  wire [14:0] _l_mask_mask_T_77 = 15'h1 << ldq_5_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_81 = 15'h3 << {12'h0, ldq_5_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_5_bits_uop_mem_size)
      2'b00:
        casez_tmp_117 = _l_mask_mask_T_77[7:0];
      2'b01:
        casez_tmp_117 = _l_mask_mask_T_81[7:0];
      2'b10:
        casez_tmp_117 = ldq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_117 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_5_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h5;
  wire        l_forwarders_5_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h5;
  wire        l_is_forwarding_5 = l_forwarders_5_0 | l_forwarders_5_1;
  wire [4:0]  l_forward_stq_idx_5 = l_is_forwarding_5 ? (l_forwarders_5_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_5_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_5_bits_forward_stq_idx;
  wire        block_addr_matches_5_1 = lcam_addr_1[39:6] == ldq_5_bits_addr_bits[39:6];
  wire        dword_addr_matches_5_0 = lcam_addr_0[39:6] == ldq_5_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_5_bits_addr_bits[5:3];
  wire        dword_addr_matches_5_1 = block_addr_matches_5_1 & lcam_addr_1[5:3] == ldq_5_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_20 = casez_tmp_117 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_22 = casez_tmp_117 & casez_tmp_109;
  wire        _GEN_447 = ldq_5_bits_executed | ldq_5_bits_succeeded;
  wire        _GEN_448 = _GEN_447 | l_is_forwarding_5;
  wire [31:0] _GEN_449 = ldq_5_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_450 = do_st_search_0 & ldq_5_valid & ldq_5_bits_addr_valid & _GEN_448 & ~ldq_5_bits_addr_is_virtual & _GEN_449[0] & dword_addr_matches_5_0 & (|_mask_overlap_T_20);
  wire        _forwarded_is_older_T_45 = l_forward_stq_idx_5 < ldq_5_bits_youngest_stq_idx;
  wire        _GEN_85586 = ~ldq_5_bits_forward_std_val | l_forward_stq_idx_5 != lcam_stq_idx_0 & (l_forward_stq_idx_5 < lcam_stq_idx_0 ^ _forwarded_is_older_T_45 ^ lcam_stq_idx_0 < ldq_5_bits_youngest_stq_idx);
  wire        _GEN_451 = _do_ld_search_T_2 & ldq_5_valid & ldq_5_bits_addr_valid & ~ldq_5_bits_addr_is_virtual & dword_addr_matches_5_0 & (|_mask_overlap_T_20);
  wire        _searcher_is_older_T_47 = ldq_head > 5'h5;
  wire        searcher_is_older_10 = lcam_ldq_idx_0 < 5'h5 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_47;
  wire        _GEN_452 = _GEN_448 & ~s1_executing_loads_5;
  wire        _GEN_85588 = _GEN_452 & ldq_5_bits_observed;
  wire        _GEN_453 = lcam_ldq_idx_0 != 5'h5;
  reg         older_nacked_REG_10;
  wire        _GEN_116700 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h5;
  wire        _GEN_454 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h5;
  wire        nacking_loads_5 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_454 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116700;
  wire        _GEN_455 = ~_GEN_447 | nacking_loads_5 | older_nacked_REG_10;
  reg         io_dmem_s1_kill_0_REG_5;
  wire        _GEN_85762 = _GEN_450 ? _GEN_85586 : _GEN_451 & searcher_is_older_10 & _GEN_85588;
  wire        _GEN_456 = _GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455);
  wire        _GEN_457 = fired_release_1 & ldq_5_valid & ldq_5_bits_addr_valid & block_addr_matches_5_1;
  wire [31:0] _GEN_458 = ldq_5_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_459 = do_st_search_1 & ldq_5_valid & ldq_5_bits_addr_valid & _GEN_448 & ~ldq_5_bits_addr_is_virtual & _GEN_458[0] & dword_addr_matches_5_1 & (|_mask_overlap_T_22);
  wire        _GEN_460 = ~ldq_5_bits_forward_std_val | l_forward_stq_idx_5 != lcam_stq_idx_1 & (l_forward_stq_idx_5 < lcam_stq_idx_1 ^ _forwarded_is_older_T_45 ^ lcam_stq_idx_1 < ldq_5_bits_youngest_stq_idx);
  wire        _GEN_461 = do_ld_search_1 & ldq_5_valid & ldq_5_bits_addr_valid & ~ldq_5_bits_addr_is_virtual & dword_addr_matches_5_1 & (|_mask_overlap_T_22);
  wire        searcher_is_older_11 = lcam_ldq_idx_1 < 5'h5 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_47;
  wire        _GEN_462 = lcam_ldq_idx_1 != 5'h5;
  reg         older_nacked_REG_11;
  wire        _GEN_463 = ~_GEN_447 | nacking_loads_5 | older_nacked_REG_11;
  reg         io_dmem_s1_kill_1_REG_5;
  wire        _GEN_464 = _GEN_461 & searcher_is_older_11 & _GEN_452 & ldq_5_bits_observed;
  wire        failed_loads_5 = _GEN_457 ? _GEN_85762 : _GEN_459 ? _GEN_460 | _GEN_85762 : _GEN_464 | _GEN_85762;
  wire        _GEN_465 = _GEN_457 | _GEN_459;
  wire        _GEN_466 = _GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463);
  wire [14:0] _l_mask_mask_T_92 = 15'h1 << ldq_6_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_96 = 15'h3 << {12'h0, ldq_6_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_6_bits_uop_mem_size)
      2'b00:
        casez_tmp_118 = _l_mask_mask_T_92[7:0];
      2'b01:
        casez_tmp_118 = _l_mask_mask_T_96[7:0];
      2'b10:
        casez_tmp_118 = ldq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_118 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_6_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h6;
  wire        l_forwarders_6_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h6;
  wire        l_is_forwarding_6 = l_forwarders_6_0 | l_forwarders_6_1;
  wire [4:0]  l_forward_stq_idx_6 = l_is_forwarding_6 ? (l_forwarders_6_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_6_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_6_bits_forward_stq_idx;
  wire        block_addr_matches_6_1 = lcam_addr_1[39:6] == ldq_6_bits_addr_bits[39:6];
  wire        dword_addr_matches_6_0 = lcam_addr_0[39:6] == ldq_6_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_6_bits_addr_bits[5:3];
  wire        dword_addr_matches_6_1 = block_addr_matches_6_1 & lcam_addr_1[5:3] == ldq_6_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_24 = casez_tmp_118 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_26 = casez_tmp_118 & casez_tmp_109;
  wire        _GEN_467 = ldq_6_bits_executed | ldq_6_bits_succeeded;
  wire        _GEN_468 = _GEN_467 | l_is_forwarding_6;
  wire [31:0] _GEN_469 = ldq_6_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_470 = do_st_search_0 & ldq_6_valid & ldq_6_bits_addr_valid & _GEN_468 & ~ldq_6_bits_addr_is_virtual & _GEN_469[0] & dword_addr_matches_6_0 & (|_mask_overlap_T_24);
  wire        _forwarded_is_older_T_53 = l_forward_stq_idx_6 < ldq_6_bits_youngest_stq_idx;
  wire        _GEN_86084 = ~ldq_6_bits_forward_std_val | l_forward_stq_idx_6 != lcam_stq_idx_0 & (l_forward_stq_idx_6 < lcam_stq_idx_0 ^ _forwarded_is_older_T_53 ^ lcam_stq_idx_0 < ldq_6_bits_youngest_stq_idx);
  wire        _GEN_471 = _do_ld_search_T_2 & ldq_6_valid & ldq_6_bits_addr_valid & ~ldq_6_bits_addr_is_virtual & dword_addr_matches_6_0 & (|_mask_overlap_T_24);
  wire        _searcher_is_older_T_55 = ldq_head > 5'h6;
  wire        searcher_is_older_12 = lcam_ldq_idx_0 < 5'h6 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_55;
  wire        _GEN_472 = _GEN_468 & ~s1_executing_loads_6;
  wire        _GEN_86086 = _GEN_472 & ldq_6_bits_observed;
  wire        _GEN_473 = lcam_ldq_idx_0 != 5'h6;
  reg         older_nacked_REG_12;
  wire        _GEN_116701 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h6;
  wire        _GEN_474 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h6;
  wire        nacking_loads_6 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_474 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116701;
  wire        _GEN_475 = ~_GEN_467 | nacking_loads_6 | older_nacked_REG_12;
  reg         io_dmem_s1_kill_0_REG_6;
  wire        _GEN_86260 = _GEN_470 ? _GEN_86084 : _GEN_471 & searcher_is_older_12 & _GEN_86086;
  wire        _GEN_476 = _GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475);
  wire        _GEN_477 = fired_release_1 & ldq_6_valid & ldq_6_bits_addr_valid & block_addr_matches_6_1;
  wire [31:0] _GEN_478 = ldq_6_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_479 = do_st_search_1 & ldq_6_valid & ldq_6_bits_addr_valid & _GEN_468 & ~ldq_6_bits_addr_is_virtual & _GEN_478[0] & dword_addr_matches_6_1 & (|_mask_overlap_T_26);
  wire        _GEN_480 = ~ldq_6_bits_forward_std_val | l_forward_stq_idx_6 != lcam_stq_idx_1 & (l_forward_stq_idx_6 < lcam_stq_idx_1 ^ _forwarded_is_older_T_53 ^ lcam_stq_idx_1 < ldq_6_bits_youngest_stq_idx);
  wire        _GEN_481 = do_ld_search_1 & ldq_6_valid & ldq_6_bits_addr_valid & ~ldq_6_bits_addr_is_virtual & dword_addr_matches_6_1 & (|_mask_overlap_T_26);
  wire        searcher_is_older_13 = lcam_ldq_idx_1 < 5'h6 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_55;
  wire        _GEN_482 = lcam_ldq_idx_1 != 5'h6;
  reg         older_nacked_REG_13;
  wire        _GEN_483 = ~_GEN_467 | nacking_loads_6 | older_nacked_REG_13;
  reg         io_dmem_s1_kill_1_REG_6;
  wire        _GEN_484 = _GEN_481 & searcher_is_older_13 & _GEN_472 & ldq_6_bits_observed;
  wire        failed_loads_6 = _GEN_477 ? _GEN_86260 : _GEN_479 ? _GEN_480 | _GEN_86260 : _GEN_484 | _GEN_86260;
  wire        _GEN_485 = _GEN_477 | _GEN_479;
  wire        _GEN_486 = _GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483);
  wire [14:0] _l_mask_mask_T_107 = 15'h1 << ldq_7_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_111 = 15'h3 << {12'h0, ldq_7_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_7_bits_uop_mem_size)
      2'b00:
        casez_tmp_119 = _l_mask_mask_T_107[7:0];
      2'b01:
        casez_tmp_119 = _l_mask_mask_T_111[7:0];
      2'b10:
        casez_tmp_119 = ldq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_119 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_7_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h7;
  wire        l_forwarders_7_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h7;
  wire        l_is_forwarding_7 = l_forwarders_7_0 | l_forwarders_7_1;
  wire [4:0]  l_forward_stq_idx_7 = l_is_forwarding_7 ? (l_forwarders_7_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_7_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_7_bits_forward_stq_idx;
  wire        block_addr_matches_7_1 = lcam_addr_1[39:6] == ldq_7_bits_addr_bits[39:6];
  wire        dword_addr_matches_7_0 = lcam_addr_0[39:6] == ldq_7_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_7_bits_addr_bits[5:3];
  wire        dword_addr_matches_7_1 = block_addr_matches_7_1 & lcam_addr_1[5:3] == ldq_7_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_28 = casez_tmp_119 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_30 = casez_tmp_119 & casez_tmp_109;
  wire        _GEN_487 = ldq_7_bits_executed | ldq_7_bits_succeeded;
  wire        _GEN_488 = _GEN_487 | l_is_forwarding_7;
  wire [31:0] _GEN_489 = ldq_7_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_490 = do_st_search_0 & ldq_7_valid & ldq_7_bits_addr_valid & _GEN_488 & ~ldq_7_bits_addr_is_virtual & _GEN_489[0] & dword_addr_matches_7_0 & (|_mask_overlap_T_28);
  wire        _forwarded_is_older_T_61 = l_forward_stq_idx_7 < ldq_7_bits_youngest_stq_idx;
  wire        _GEN_86582 = ~ldq_7_bits_forward_std_val | l_forward_stq_idx_7 != lcam_stq_idx_0 & (l_forward_stq_idx_7 < lcam_stq_idx_0 ^ _forwarded_is_older_T_61 ^ lcam_stq_idx_0 < ldq_7_bits_youngest_stq_idx);
  wire        _GEN_491 = _do_ld_search_T_2 & ldq_7_valid & ldq_7_bits_addr_valid & ~ldq_7_bits_addr_is_virtual & dword_addr_matches_7_0 & (|_mask_overlap_T_28);
  wire        searcher_is_older_14 = lcam_ldq_idx_0 < 5'h7 ^ _searcher_is_older_T_249 ^ (|(ldq_head[4:3]));
  wire        _GEN_492 = _GEN_488 & ~s1_executing_loads_7;
  wire        _GEN_86584 = _GEN_492 & ldq_7_bits_observed;
  wire        _GEN_493 = lcam_ldq_idx_0 != 5'h7;
  reg         older_nacked_REG_14;
  wire        _GEN_116702 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h7;
  wire        _GEN_494 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h7;
  wire        nacking_loads_7 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_494 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116702;
  wire        _GEN_495 = ~_GEN_487 | nacking_loads_7 | older_nacked_REG_14;
  reg         io_dmem_s1_kill_0_REG_7;
  wire        _GEN_86758 = _GEN_490 ? _GEN_86582 : _GEN_491 & searcher_is_older_14 & _GEN_86584;
  wire        _GEN_496 = _GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495);
  wire        _GEN_497 = fired_release_1 & ldq_7_valid & ldq_7_bits_addr_valid & block_addr_matches_7_1;
  wire [31:0] _GEN_498 = ldq_7_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_499 = do_st_search_1 & ldq_7_valid & ldq_7_bits_addr_valid & _GEN_488 & ~ldq_7_bits_addr_is_virtual & _GEN_498[0] & dword_addr_matches_7_1 & (|_mask_overlap_T_30);
  wire        _GEN_500 = ~ldq_7_bits_forward_std_val | l_forward_stq_idx_7 != lcam_stq_idx_1 & (l_forward_stq_idx_7 < lcam_stq_idx_1 ^ _forwarded_is_older_T_61 ^ lcam_stq_idx_1 < ldq_7_bits_youngest_stq_idx);
  wire        _GEN_501 = do_ld_search_1 & ldq_7_valid & ldq_7_bits_addr_valid & ~ldq_7_bits_addr_is_virtual & dword_addr_matches_7_1 & (|_mask_overlap_T_30);
  wire        searcher_is_older_15 = lcam_ldq_idx_1 < 5'h7 ^ _searcher_is_older_T_253 ^ (|(ldq_head[4:3]));
  wire        _GEN_502 = lcam_ldq_idx_1 != 5'h7;
  reg         older_nacked_REG_15;
  wire        _GEN_503 = ~_GEN_487 | nacking_loads_7 | older_nacked_REG_15;
  reg         io_dmem_s1_kill_1_REG_7;
  wire        _GEN_504 = _GEN_501 & searcher_is_older_15 & _GEN_492 & ldq_7_bits_observed;
  wire        failed_loads_7 = _GEN_497 ? _GEN_86758 : _GEN_499 ? _GEN_500 | _GEN_86758 : _GEN_504 | _GEN_86758;
  wire        _GEN_505 = _GEN_497 | _GEN_499;
  wire        _GEN_506 = _GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503);
  wire [14:0] _l_mask_mask_T_122 = 15'h1 << ldq_8_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_126 = 15'h3 << {12'h0, ldq_8_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_8_bits_uop_mem_size)
      2'b00:
        casez_tmp_120 = _l_mask_mask_T_122[7:0];
      2'b01:
        casez_tmp_120 = _l_mask_mask_T_126[7:0];
      2'b10:
        casez_tmp_120 = ldq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_120 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_8_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h8;
  wire        l_forwarders_8_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h8;
  wire        l_is_forwarding_8 = l_forwarders_8_0 | l_forwarders_8_1;
  wire [4:0]  l_forward_stq_idx_8 = l_is_forwarding_8 ? (l_forwarders_8_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_8_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_8_bits_forward_stq_idx;
  wire        block_addr_matches_8_1 = lcam_addr_1[39:6] == ldq_8_bits_addr_bits[39:6];
  wire        dword_addr_matches_8_0 = lcam_addr_0[39:6] == ldq_8_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_8_bits_addr_bits[5:3];
  wire        dword_addr_matches_8_1 = block_addr_matches_8_1 & lcam_addr_1[5:3] == ldq_8_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_32 = casez_tmp_120 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_34 = casez_tmp_120 & casez_tmp_109;
  wire        _GEN_507 = ldq_8_bits_executed | ldq_8_bits_succeeded;
  wire        _GEN_508 = _GEN_507 | l_is_forwarding_8;
  wire [31:0] _GEN_509 = ldq_8_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_510 = do_st_search_0 & ldq_8_valid & ldq_8_bits_addr_valid & _GEN_508 & ~ldq_8_bits_addr_is_virtual & _GEN_509[0] & dword_addr_matches_8_0 & (|_mask_overlap_T_32);
  wire        _forwarded_is_older_T_69 = l_forward_stq_idx_8 < ldq_8_bits_youngest_stq_idx;
  wire        _GEN_87080 = ~ldq_8_bits_forward_std_val | l_forward_stq_idx_8 != lcam_stq_idx_0 & (l_forward_stq_idx_8 < lcam_stq_idx_0 ^ _forwarded_is_older_T_69 ^ lcam_stq_idx_0 < ldq_8_bits_youngest_stq_idx);
  wire        _GEN_511 = _do_ld_search_T_2 & ldq_8_valid & ldq_8_bits_addr_valid & ~ldq_8_bits_addr_is_virtual & dword_addr_matches_8_0 & (|_mask_overlap_T_32);
  wire        _searcher_is_older_T_71 = ldq_head > 5'h8;
  wire        searcher_is_older_16 = lcam_ldq_idx_0 < 5'h8 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_71;
  wire        _GEN_512 = _GEN_508 & ~s1_executing_loads_8;
  wire        _GEN_87082 = _GEN_512 & ldq_8_bits_observed;
  wire        _GEN_513 = lcam_ldq_idx_0 != 5'h8;
  reg         older_nacked_REG_16;
  wire        _GEN_116703 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h8;
  wire        _GEN_514 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h8;
  wire        nacking_loads_8 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_514 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116703;
  wire        _GEN_515 = ~_GEN_507 | nacking_loads_8 | older_nacked_REG_16;
  reg         io_dmem_s1_kill_0_REG_8;
  wire        _GEN_87256 = _GEN_510 ? _GEN_87080 : _GEN_511 & searcher_is_older_16 & _GEN_87082;
  wire        _GEN_516 = _GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515);
  wire        _GEN_517 = fired_release_1 & ldq_8_valid & ldq_8_bits_addr_valid & block_addr_matches_8_1;
  wire [31:0] _GEN_518 = ldq_8_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_519 = do_st_search_1 & ldq_8_valid & ldq_8_bits_addr_valid & _GEN_508 & ~ldq_8_bits_addr_is_virtual & _GEN_518[0] & dword_addr_matches_8_1 & (|_mask_overlap_T_34);
  wire        _GEN_520 = ~ldq_8_bits_forward_std_val | l_forward_stq_idx_8 != lcam_stq_idx_1 & (l_forward_stq_idx_8 < lcam_stq_idx_1 ^ _forwarded_is_older_T_69 ^ lcam_stq_idx_1 < ldq_8_bits_youngest_stq_idx);
  wire        _GEN_521 = do_ld_search_1 & ldq_8_valid & ldq_8_bits_addr_valid & ~ldq_8_bits_addr_is_virtual & dword_addr_matches_8_1 & (|_mask_overlap_T_34);
  wire        searcher_is_older_17 = lcam_ldq_idx_1 < 5'h8 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_71;
  wire        _GEN_522 = lcam_ldq_idx_1 != 5'h8;
  reg         older_nacked_REG_17;
  wire        _GEN_523 = ~_GEN_507 | nacking_loads_8 | older_nacked_REG_17;
  reg         io_dmem_s1_kill_1_REG_8;
  wire        _GEN_524 = _GEN_521 & searcher_is_older_17 & _GEN_512 & ldq_8_bits_observed;
  wire        failed_loads_8 = _GEN_517 ? _GEN_87256 : _GEN_519 ? _GEN_520 | _GEN_87256 : _GEN_524 | _GEN_87256;
  wire        _GEN_525 = _GEN_517 | _GEN_519;
  wire        _GEN_526 = _GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523);
  wire [14:0] _l_mask_mask_T_137 = 15'h1 << ldq_9_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_141 = 15'h3 << {12'h0, ldq_9_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_9_bits_uop_mem_size)
      2'b00:
        casez_tmp_121 = _l_mask_mask_T_137[7:0];
      2'b01:
        casez_tmp_121 = _l_mask_mask_T_141[7:0];
      2'b10:
        casez_tmp_121 = ldq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_121 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_9_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h9;
  wire        l_forwarders_9_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h9;
  wire        l_is_forwarding_9 = l_forwarders_9_0 | l_forwarders_9_1;
  wire [4:0]  l_forward_stq_idx_9 = l_is_forwarding_9 ? (l_forwarders_9_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_9_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_9_bits_forward_stq_idx;
  wire        block_addr_matches_9_1 = lcam_addr_1[39:6] == ldq_9_bits_addr_bits[39:6];
  wire        dword_addr_matches_9_0 = lcam_addr_0[39:6] == ldq_9_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_9_bits_addr_bits[5:3];
  wire        dword_addr_matches_9_1 = block_addr_matches_9_1 & lcam_addr_1[5:3] == ldq_9_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_36 = casez_tmp_121 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_38 = casez_tmp_121 & casez_tmp_109;
  wire        _GEN_527 = ldq_9_bits_executed | ldq_9_bits_succeeded;
  wire        _GEN_528 = _GEN_527 | l_is_forwarding_9;
  wire [31:0] _GEN_529 = ldq_9_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_530 = do_st_search_0 & ldq_9_valid & ldq_9_bits_addr_valid & _GEN_528 & ~ldq_9_bits_addr_is_virtual & _GEN_529[0] & dword_addr_matches_9_0 & (|_mask_overlap_T_36);
  wire        _forwarded_is_older_T_77 = l_forward_stq_idx_9 < ldq_9_bits_youngest_stq_idx;
  wire        _GEN_87578 = ~ldq_9_bits_forward_std_val | l_forward_stq_idx_9 != lcam_stq_idx_0 & (l_forward_stq_idx_9 < lcam_stq_idx_0 ^ _forwarded_is_older_T_77 ^ lcam_stq_idx_0 < ldq_9_bits_youngest_stq_idx);
  wire        _GEN_531 = _do_ld_search_T_2 & ldq_9_valid & ldq_9_bits_addr_valid & ~ldq_9_bits_addr_is_virtual & dword_addr_matches_9_0 & (|_mask_overlap_T_36);
  wire        _searcher_is_older_T_79 = ldq_head > 5'h9;
  wire        searcher_is_older_18 = lcam_ldq_idx_0 < 5'h9 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_79;
  wire        _GEN_532 = _GEN_528 & ~s1_executing_loads_9;
  wire        _GEN_87580 = _GEN_532 & ldq_9_bits_observed;
  wire        _GEN_533 = lcam_ldq_idx_0 != 5'h9;
  reg         older_nacked_REG_18;
  wire        _GEN_116704 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h9;
  wire        _GEN_534 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h9;
  wire        nacking_loads_9 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_534 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116704;
  wire        _GEN_535 = ~_GEN_527 | nacking_loads_9 | older_nacked_REG_18;
  reg         io_dmem_s1_kill_0_REG_9;
  wire        _GEN_87754 = _GEN_530 ? _GEN_87578 : _GEN_531 & searcher_is_older_18 & _GEN_87580;
  wire        _GEN_536 = _GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535);
  wire        _GEN_537 = fired_release_1 & ldq_9_valid & ldq_9_bits_addr_valid & block_addr_matches_9_1;
  wire [31:0] _GEN_538 = ldq_9_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_539 = do_st_search_1 & ldq_9_valid & ldq_9_bits_addr_valid & _GEN_528 & ~ldq_9_bits_addr_is_virtual & _GEN_538[0] & dword_addr_matches_9_1 & (|_mask_overlap_T_38);
  wire        _GEN_540 = ~ldq_9_bits_forward_std_val | l_forward_stq_idx_9 != lcam_stq_idx_1 & (l_forward_stq_idx_9 < lcam_stq_idx_1 ^ _forwarded_is_older_T_77 ^ lcam_stq_idx_1 < ldq_9_bits_youngest_stq_idx);
  wire        _GEN_541 = do_ld_search_1 & ldq_9_valid & ldq_9_bits_addr_valid & ~ldq_9_bits_addr_is_virtual & dword_addr_matches_9_1 & (|_mask_overlap_T_38);
  wire        searcher_is_older_19 = lcam_ldq_idx_1 < 5'h9 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_79;
  wire        _GEN_542 = lcam_ldq_idx_1 != 5'h9;
  reg         older_nacked_REG_19;
  wire        _GEN_543 = ~_GEN_527 | nacking_loads_9 | older_nacked_REG_19;
  reg         io_dmem_s1_kill_1_REG_9;
  wire        _GEN_544 = _GEN_541 & searcher_is_older_19 & _GEN_532 & ldq_9_bits_observed;
  wire        failed_loads_9 = _GEN_537 ? _GEN_87754 : _GEN_539 ? _GEN_540 | _GEN_87754 : _GEN_544 | _GEN_87754;
  wire        _GEN_545 = _GEN_537 | _GEN_539;
  wire        _GEN_546 = _GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543);
  wire [14:0] _l_mask_mask_T_152 = 15'h1 << ldq_10_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_156 = 15'h3 << {12'h0, ldq_10_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_10_bits_uop_mem_size)
      2'b00:
        casez_tmp_122 = _l_mask_mask_T_152[7:0];
      2'b01:
        casez_tmp_122 = _l_mask_mask_T_156[7:0];
      2'b10:
        casez_tmp_122 = ldq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_122 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_10_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hA;
  wire        l_forwarders_10_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hA;
  wire        l_is_forwarding_10 = l_forwarders_10_0 | l_forwarders_10_1;
  wire [4:0]  l_forward_stq_idx_10 = l_is_forwarding_10 ? (l_forwarders_10_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_10_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_10_bits_forward_stq_idx;
  wire        block_addr_matches_10_1 = lcam_addr_1[39:6] == ldq_10_bits_addr_bits[39:6];
  wire        dword_addr_matches_10_0 = lcam_addr_0[39:6] == ldq_10_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_10_bits_addr_bits[5:3];
  wire        dword_addr_matches_10_1 = block_addr_matches_10_1 & lcam_addr_1[5:3] == ldq_10_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_40 = casez_tmp_122 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_42 = casez_tmp_122 & casez_tmp_109;
  wire        _GEN_547 = ldq_10_bits_executed | ldq_10_bits_succeeded;
  wire        _GEN_548 = _GEN_547 | l_is_forwarding_10;
  wire [31:0] _GEN_549 = ldq_10_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_550 = do_st_search_0 & ldq_10_valid & ldq_10_bits_addr_valid & _GEN_548 & ~ldq_10_bits_addr_is_virtual & _GEN_549[0] & dword_addr_matches_10_0 & (|_mask_overlap_T_40);
  wire        _forwarded_is_older_T_85 = l_forward_stq_idx_10 < ldq_10_bits_youngest_stq_idx;
  wire        _GEN_88076 = ~ldq_10_bits_forward_std_val | l_forward_stq_idx_10 != lcam_stq_idx_0 & (l_forward_stq_idx_10 < lcam_stq_idx_0 ^ _forwarded_is_older_T_85 ^ lcam_stq_idx_0 < ldq_10_bits_youngest_stq_idx);
  wire        _GEN_551 = _do_ld_search_T_2 & ldq_10_valid & ldq_10_bits_addr_valid & ~ldq_10_bits_addr_is_virtual & dword_addr_matches_10_0 & (|_mask_overlap_T_40);
  wire        _searcher_is_older_T_87 = ldq_head > 5'hA;
  wire        searcher_is_older_20 = lcam_ldq_idx_0 < 5'hA ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_87;
  wire        _GEN_552 = _GEN_548 & ~s1_executing_loads_10;
  wire        _GEN_88078 = _GEN_552 & ldq_10_bits_observed;
  wire        _GEN_553 = lcam_ldq_idx_0 != 5'hA;
  reg         older_nacked_REG_20;
  wire        _GEN_116705 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hA;
  wire        _GEN_554 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hA;
  wire        nacking_loads_10 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_554 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116705;
  wire        _GEN_555 = ~_GEN_547 | nacking_loads_10 | older_nacked_REG_20;
  reg         io_dmem_s1_kill_0_REG_10;
  wire        _GEN_88252 = _GEN_550 ? _GEN_88076 : _GEN_551 & searcher_is_older_20 & _GEN_88078;
  wire        _GEN_556 = _GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555);
  wire        _GEN_557 = fired_release_1 & ldq_10_valid & ldq_10_bits_addr_valid & block_addr_matches_10_1;
  wire [31:0] _GEN_558 = ldq_10_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_559 = do_st_search_1 & ldq_10_valid & ldq_10_bits_addr_valid & _GEN_548 & ~ldq_10_bits_addr_is_virtual & _GEN_558[0] & dword_addr_matches_10_1 & (|_mask_overlap_T_42);
  wire        _GEN_560 = ~ldq_10_bits_forward_std_val | l_forward_stq_idx_10 != lcam_stq_idx_1 & (l_forward_stq_idx_10 < lcam_stq_idx_1 ^ _forwarded_is_older_T_85 ^ lcam_stq_idx_1 < ldq_10_bits_youngest_stq_idx);
  wire        _GEN_561 = do_ld_search_1 & ldq_10_valid & ldq_10_bits_addr_valid & ~ldq_10_bits_addr_is_virtual & dword_addr_matches_10_1 & (|_mask_overlap_T_42);
  wire        searcher_is_older_21 = lcam_ldq_idx_1 < 5'hA ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_87;
  wire        _GEN_562 = lcam_ldq_idx_1 != 5'hA;
  reg         older_nacked_REG_21;
  wire        _GEN_563 = ~_GEN_547 | nacking_loads_10 | older_nacked_REG_21;
  reg         io_dmem_s1_kill_1_REG_10;
  wire        _GEN_564 = _GEN_561 & searcher_is_older_21 & _GEN_552 & ldq_10_bits_observed;
  wire        failed_loads_10 = _GEN_557 ? _GEN_88252 : _GEN_559 ? _GEN_560 | _GEN_88252 : _GEN_564 | _GEN_88252;
  wire        _GEN_565 = _GEN_557 | _GEN_559;
  wire        _GEN_566 = _GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563);
  wire [14:0] _l_mask_mask_T_167 = 15'h1 << ldq_11_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_171 = 15'h3 << {12'h0, ldq_11_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_11_bits_uop_mem_size)
      2'b00:
        casez_tmp_123 = _l_mask_mask_T_167[7:0];
      2'b01:
        casez_tmp_123 = _l_mask_mask_T_171[7:0];
      2'b10:
        casez_tmp_123 = ldq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_123 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_11_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hB;
  wire        l_forwarders_11_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hB;
  wire        l_is_forwarding_11 = l_forwarders_11_0 | l_forwarders_11_1;
  wire [4:0]  l_forward_stq_idx_11 = l_is_forwarding_11 ? (l_forwarders_11_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_11_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_11_bits_forward_stq_idx;
  wire        block_addr_matches_11_1 = lcam_addr_1[39:6] == ldq_11_bits_addr_bits[39:6];
  wire        dword_addr_matches_11_0 = lcam_addr_0[39:6] == ldq_11_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_11_bits_addr_bits[5:3];
  wire        dword_addr_matches_11_1 = block_addr_matches_11_1 & lcam_addr_1[5:3] == ldq_11_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_44 = casez_tmp_123 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_46 = casez_tmp_123 & casez_tmp_109;
  wire        _GEN_567 = ldq_11_bits_executed | ldq_11_bits_succeeded;
  wire        _GEN_568 = _GEN_567 | l_is_forwarding_11;
  wire [31:0] _GEN_569 = ldq_11_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_570 = do_st_search_0 & ldq_11_valid & ldq_11_bits_addr_valid & _GEN_568 & ~ldq_11_bits_addr_is_virtual & _GEN_569[0] & dword_addr_matches_11_0 & (|_mask_overlap_T_44);
  wire        _forwarded_is_older_T_93 = l_forward_stq_idx_11 < ldq_11_bits_youngest_stq_idx;
  wire        _GEN_88574 = ~ldq_11_bits_forward_std_val | l_forward_stq_idx_11 != lcam_stq_idx_0 & (l_forward_stq_idx_11 < lcam_stq_idx_0 ^ _forwarded_is_older_T_93 ^ lcam_stq_idx_0 < ldq_11_bits_youngest_stq_idx);
  wire        _GEN_571 = _do_ld_search_T_2 & ldq_11_valid & ldq_11_bits_addr_valid & ~ldq_11_bits_addr_is_virtual & dword_addr_matches_11_0 & (|_mask_overlap_T_44);
  wire        _searcher_is_older_T_95 = ldq_head > 5'hB;
  wire        searcher_is_older_22 = lcam_ldq_idx_0 < 5'hB ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_95;
  wire        _GEN_572 = _GEN_568 & ~s1_executing_loads_11;
  wire        _GEN_88576 = _GEN_572 & ldq_11_bits_observed;
  wire        _GEN_573 = lcam_ldq_idx_0 != 5'hB;
  reg         older_nacked_REG_22;
  wire        _GEN_116706 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hB;
  wire        _GEN_574 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hB;
  wire        nacking_loads_11 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_574 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116706;
  wire        _GEN_575 = ~_GEN_567 | nacking_loads_11 | older_nacked_REG_22;
  reg         io_dmem_s1_kill_0_REG_11;
  wire        _GEN_88750 = _GEN_570 ? _GEN_88574 : _GEN_571 & searcher_is_older_22 & _GEN_88576;
  wire        _GEN_576 = _GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575);
  wire        _GEN_577 = fired_release_1 & ldq_11_valid & ldq_11_bits_addr_valid & block_addr_matches_11_1;
  wire [31:0] _GEN_578 = ldq_11_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_579 = do_st_search_1 & ldq_11_valid & ldq_11_bits_addr_valid & _GEN_568 & ~ldq_11_bits_addr_is_virtual & _GEN_578[0] & dword_addr_matches_11_1 & (|_mask_overlap_T_46);
  wire        _GEN_580 = ~ldq_11_bits_forward_std_val | l_forward_stq_idx_11 != lcam_stq_idx_1 & (l_forward_stq_idx_11 < lcam_stq_idx_1 ^ _forwarded_is_older_T_93 ^ lcam_stq_idx_1 < ldq_11_bits_youngest_stq_idx);
  wire        _GEN_581 = do_ld_search_1 & ldq_11_valid & ldq_11_bits_addr_valid & ~ldq_11_bits_addr_is_virtual & dword_addr_matches_11_1 & (|_mask_overlap_T_46);
  wire        searcher_is_older_23 = lcam_ldq_idx_1 < 5'hB ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_95;
  wire        _GEN_582 = lcam_ldq_idx_1 != 5'hB;
  reg         older_nacked_REG_23;
  wire        _GEN_583 = ~_GEN_567 | nacking_loads_11 | older_nacked_REG_23;
  reg         io_dmem_s1_kill_1_REG_11;
  wire        _GEN_584 = _GEN_581 & searcher_is_older_23 & _GEN_572 & ldq_11_bits_observed;
  wire        failed_loads_11 = _GEN_577 ? _GEN_88750 : _GEN_579 ? _GEN_580 | _GEN_88750 : _GEN_584 | _GEN_88750;
  wire        _GEN_585 = _GEN_577 | _GEN_579;
  wire        _GEN_586 = _GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583);
  wire [14:0] _l_mask_mask_T_182 = 15'h1 << ldq_12_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_186 = 15'h3 << {12'h0, ldq_12_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_12_bits_uop_mem_size)
      2'b00:
        casez_tmp_124 = _l_mask_mask_T_182[7:0];
      2'b01:
        casez_tmp_124 = _l_mask_mask_T_186[7:0];
      2'b10:
        casez_tmp_124 = ldq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_124 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_12_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hC;
  wire        l_forwarders_12_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hC;
  wire        l_is_forwarding_12 = l_forwarders_12_0 | l_forwarders_12_1;
  wire [4:0]  l_forward_stq_idx_12 = l_is_forwarding_12 ? (l_forwarders_12_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_12_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_12_bits_forward_stq_idx;
  wire        block_addr_matches_12_1 = lcam_addr_1[39:6] == ldq_12_bits_addr_bits[39:6];
  wire        dword_addr_matches_12_0 = lcam_addr_0[39:6] == ldq_12_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_12_bits_addr_bits[5:3];
  wire        dword_addr_matches_12_1 = block_addr_matches_12_1 & lcam_addr_1[5:3] == ldq_12_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_48 = casez_tmp_124 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_50 = casez_tmp_124 & casez_tmp_109;
  wire        _GEN_587 = ldq_12_bits_executed | ldq_12_bits_succeeded;
  wire        _GEN_588 = _GEN_587 | l_is_forwarding_12;
  wire [31:0] _GEN_589 = ldq_12_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_590 = do_st_search_0 & ldq_12_valid & ldq_12_bits_addr_valid & _GEN_588 & ~ldq_12_bits_addr_is_virtual & _GEN_589[0] & dword_addr_matches_12_0 & (|_mask_overlap_T_48);
  wire        _forwarded_is_older_T_101 = l_forward_stq_idx_12 < ldq_12_bits_youngest_stq_idx;
  wire        _GEN_89072 = ~ldq_12_bits_forward_std_val | l_forward_stq_idx_12 != lcam_stq_idx_0 & (l_forward_stq_idx_12 < lcam_stq_idx_0 ^ _forwarded_is_older_T_101 ^ lcam_stq_idx_0 < ldq_12_bits_youngest_stq_idx);
  wire        _GEN_591 = _do_ld_search_T_2 & ldq_12_valid & ldq_12_bits_addr_valid & ~ldq_12_bits_addr_is_virtual & dword_addr_matches_12_0 & (|_mask_overlap_T_48);
  wire        _searcher_is_older_T_103 = ldq_head > 5'hC;
  wire        searcher_is_older_24 = lcam_ldq_idx_0 < 5'hC ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_103;
  wire        _GEN_592 = _GEN_588 & ~s1_executing_loads_12;
  wire        _GEN_89074 = _GEN_592 & ldq_12_bits_observed;
  wire        _GEN_593 = lcam_ldq_idx_0 != 5'hC;
  reg         older_nacked_REG_24;
  wire        _GEN_116707 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hC;
  wire        _GEN_594 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hC;
  wire        nacking_loads_12 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_594 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116707;
  wire        _GEN_595 = ~_GEN_587 | nacking_loads_12 | older_nacked_REG_24;
  reg         io_dmem_s1_kill_0_REG_12;
  wire        _GEN_89248 = _GEN_590 ? _GEN_89072 : _GEN_591 & searcher_is_older_24 & _GEN_89074;
  wire        _GEN_596 = _GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595);
  wire        _GEN_597 = fired_release_1 & ldq_12_valid & ldq_12_bits_addr_valid & block_addr_matches_12_1;
  wire [31:0] _GEN_598 = ldq_12_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_599 = do_st_search_1 & ldq_12_valid & ldq_12_bits_addr_valid & _GEN_588 & ~ldq_12_bits_addr_is_virtual & _GEN_598[0] & dword_addr_matches_12_1 & (|_mask_overlap_T_50);
  wire        _GEN_600 = ~ldq_12_bits_forward_std_val | l_forward_stq_idx_12 != lcam_stq_idx_1 & (l_forward_stq_idx_12 < lcam_stq_idx_1 ^ _forwarded_is_older_T_101 ^ lcam_stq_idx_1 < ldq_12_bits_youngest_stq_idx);
  wire        _GEN_601 = do_ld_search_1 & ldq_12_valid & ldq_12_bits_addr_valid & ~ldq_12_bits_addr_is_virtual & dword_addr_matches_12_1 & (|_mask_overlap_T_50);
  wire        searcher_is_older_25 = lcam_ldq_idx_1 < 5'hC ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_103;
  wire        _GEN_602 = lcam_ldq_idx_1 != 5'hC;
  reg         older_nacked_REG_25;
  wire        _GEN_603 = ~_GEN_587 | nacking_loads_12 | older_nacked_REG_25;
  reg         io_dmem_s1_kill_1_REG_12;
  wire        _GEN_604 = _GEN_601 & searcher_is_older_25 & _GEN_592 & ldq_12_bits_observed;
  wire        failed_loads_12 = _GEN_597 ? _GEN_89248 : _GEN_599 ? _GEN_600 | _GEN_89248 : _GEN_604 | _GEN_89248;
  wire        _GEN_605 = _GEN_597 | _GEN_599;
  wire        _GEN_606 = _GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603);
  wire [14:0] _l_mask_mask_T_197 = 15'h1 << ldq_13_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_201 = 15'h3 << {12'h0, ldq_13_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_13_bits_uop_mem_size)
      2'b00:
        casez_tmp_125 = _l_mask_mask_T_197[7:0];
      2'b01:
        casez_tmp_125 = _l_mask_mask_T_201[7:0];
      2'b10:
        casez_tmp_125 = ldq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_125 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_13_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hD;
  wire        l_forwarders_13_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hD;
  wire        l_is_forwarding_13 = l_forwarders_13_0 | l_forwarders_13_1;
  wire [4:0]  l_forward_stq_idx_13 = l_is_forwarding_13 ? (l_forwarders_13_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_13_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_13_bits_forward_stq_idx;
  wire        block_addr_matches_13_1 = lcam_addr_1[39:6] == ldq_13_bits_addr_bits[39:6];
  wire        dword_addr_matches_13_0 = lcam_addr_0[39:6] == ldq_13_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_13_bits_addr_bits[5:3];
  wire        dword_addr_matches_13_1 = block_addr_matches_13_1 & lcam_addr_1[5:3] == ldq_13_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_52 = casez_tmp_125 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_54 = casez_tmp_125 & casez_tmp_109;
  wire        _GEN_607 = ldq_13_bits_executed | ldq_13_bits_succeeded;
  wire        _GEN_608 = _GEN_607 | l_is_forwarding_13;
  wire [31:0] _GEN_609 = ldq_13_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_610 = do_st_search_0 & ldq_13_valid & ldq_13_bits_addr_valid & _GEN_608 & ~ldq_13_bits_addr_is_virtual & _GEN_609[0] & dword_addr_matches_13_0 & (|_mask_overlap_T_52);
  wire        _forwarded_is_older_T_109 = l_forward_stq_idx_13 < ldq_13_bits_youngest_stq_idx;
  wire        _GEN_89570 = ~ldq_13_bits_forward_std_val | l_forward_stq_idx_13 != lcam_stq_idx_0 & (l_forward_stq_idx_13 < lcam_stq_idx_0 ^ _forwarded_is_older_T_109 ^ lcam_stq_idx_0 < ldq_13_bits_youngest_stq_idx);
  wire        _GEN_611 = _do_ld_search_T_2 & ldq_13_valid & ldq_13_bits_addr_valid & ~ldq_13_bits_addr_is_virtual & dword_addr_matches_13_0 & (|_mask_overlap_T_52);
  wire        _searcher_is_older_T_111 = ldq_head > 5'hD;
  wire        searcher_is_older_26 = lcam_ldq_idx_0 < 5'hD ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_111;
  wire        _GEN_612 = _GEN_608 & ~s1_executing_loads_13;
  wire        _GEN_89572 = _GEN_612 & ldq_13_bits_observed;
  wire        _GEN_613 = lcam_ldq_idx_0 != 5'hD;
  reg         older_nacked_REG_26;
  wire        _GEN_116708 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hD;
  wire        _GEN_614 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hD;
  wire        nacking_loads_13 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_614 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116708;
  wire        _GEN_615 = ~_GEN_607 | nacking_loads_13 | older_nacked_REG_26;
  reg         io_dmem_s1_kill_0_REG_13;
  wire        _GEN_89746 = _GEN_610 ? _GEN_89570 : _GEN_611 & searcher_is_older_26 & _GEN_89572;
  wire        _GEN_616 = _GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615);
  wire        _GEN_617 = fired_release_1 & ldq_13_valid & ldq_13_bits_addr_valid & block_addr_matches_13_1;
  wire [31:0] _GEN_618 = ldq_13_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_619 = do_st_search_1 & ldq_13_valid & ldq_13_bits_addr_valid & _GEN_608 & ~ldq_13_bits_addr_is_virtual & _GEN_618[0] & dword_addr_matches_13_1 & (|_mask_overlap_T_54);
  wire        _GEN_620 = ~ldq_13_bits_forward_std_val | l_forward_stq_idx_13 != lcam_stq_idx_1 & (l_forward_stq_idx_13 < lcam_stq_idx_1 ^ _forwarded_is_older_T_109 ^ lcam_stq_idx_1 < ldq_13_bits_youngest_stq_idx);
  wire        _GEN_621 = do_ld_search_1 & ldq_13_valid & ldq_13_bits_addr_valid & ~ldq_13_bits_addr_is_virtual & dword_addr_matches_13_1 & (|_mask_overlap_T_54);
  wire        searcher_is_older_27 = lcam_ldq_idx_1 < 5'hD ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_111;
  wire        _GEN_622 = lcam_ldq_idx_1 != 5'hD;
  reg         older_nacked_REG_27;
  wire        _GEN_623 = ~_GEN_607 | nacking_loads_13 | older_nacked_REG_27;
  reg         io_dmem_s1_kill_1_REG_13;
  wire        _GEN_624 = _GEN_621 & searcher_is_older_27 & _GEN_612 & ldq_13_bits_observed;
  wire        failed_loads_13 = _GEN_617 ? _GEN_89746 : _GEN_619 ? _GEN_620 | _GEN_89746 : _GEN_624 | _GEN_89746;
  wire        _GEN_625 = _GEN_617 | _GEN_619;
  wire        _GEN_626 = _GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623);
  wire [14:0] _l_mask_mask_T_212 = 15'h1 << ldq_14_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_216 = 15'h3 << {12'h0, ldq_14_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_14_bits_uop_mem_size)
      2'b00:
        casez_tmp_126 = _l_mask_mask_T_212[7:0];
      2'b01:
        casez_tmp_126 = _l_mask_mask_T_216[7:0];
      2'b10:
        casez_tmp_126 = ldq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_126 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_14_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hE;
  wire        l_forwarders_14_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hE;
  wire        l_is_forwarding_14 = l_forwarders_14_0 | l_forwarders_14_1;
  wire [4:0]  l_forward_stq_idx_14 = l_is_forwarding_14 ? (l_forwarders_14_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_14_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_14_bits_forward_stq_idx;
  wire        block_addr_matches_14_1 = lcam_addr_1[39:6] == ldq_14_bits_addr_bits[39:6];
  wire        dword_addr_matches_14_0 = lcam_addr_0[39:6] == ldq_14_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_14_bits_addr_bits[5:3];
  wire        dword_addr_matches_14_1 = block_addr_matches_14_1 & lcam_addr_1[5:3] == ldq_14_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_56 = casez_tmp_126 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_58 = casez_tmp_126 & casez_tmp_109;
  wire        _GEN_627 = ldq_14_bits_executed | ldq_14_bits_succeeded;
  wire        _GEN_628 = _GEN_627 | l_is_forwarding_14;
  wire [31:0] _GEN_629 = ldq_14_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_630 = do_st_search_0 & ldq_14_valid & ldq_14_bits_addr_valid & _GEN_628 & ~ldq_14_bits_addr_is_virtual & _GEN_629[0] & dword_addr_matches_14_0 & (|_mask_overlap_T_56);
  wire        _forwarded_is_older_T_117 = l_forward_stq_idx_14 < ldq_14_bits_youngest_stq_idx;
  wire        _GEN_90068 = ~ldq_14_bits_forward_std_val | l_forward_stq_idx_14 != lcam_stq_idx_0 & (l_forward_stq_idx_14 < lcam_stq_idx_0 ^ _forwarded_is_older_T_117 ^ lcam_stq_idx_0 < ldq_14_bits_youngest_stq_idx);
  wire        _GEN_631 = _do_ld_search_T_2 & ldq_14_valid & ldq_14_bits_addr_valid & ~ldq_14_bits_addr_is_virtual & dword_addr_matches_14_0 & (|_mask_overlap_T_56);
  wire        _searcher_is_older_T_119 = ldq_head > 5'hE;
  wire        searcher_is_older_28 = lcam_ldq_idx_0 < 5'hE ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_119;
  wire        _GEN_632 = _GEN_628 & ~s1_executing_loads_14;
  wire        _GEN_90070 = _GEN_632 & ldq_14_bits_observed;
  wire        _GEN_633 = lcam_ldq_idx_0 != 5'hE;
  reg         older_nacked_REG_28;
  wire        _GEN_116709 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hE;
  wire        _GEN_634 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hE;
  wire        nacking_loads_14 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_634 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116709;
  wire        _GEN_635 = ~_GEN_627 | nacking_loads_14 | older_nacked_REG_28;
  reg         io_dmem_s1_kill_0_REG_14;
  wire        _GEN_90244 = _GEN_630 ? _GEN_90068 : _GEN_631 & searcher_is_older_28 & _GEN_90070;
  wire        _GEN_636 = _GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635);
  wire        _GEN_637 = fired_release_1 & ldq_14_valid & ldq_14_bits_addr_valid & block_addr_matches_14_1;
  wire [31:0] _GEN_638 = ldq_14_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_639 = do_st_search_1 & ldq_14_valid & ldq_14_bits_addr_valid & _GEN_628 & ~ldq_14_bits_addr_is_virtual & _GEN_638[0] & dword_addr_matches_14_1 & (|_mask_overlap_T_58);
  wire        _GEN_640 = ~ldq_14_bits_forward_std_val | l_forward_stq_idx_14 != lcam_stq_idx_1 & (l_forward_stq_idx_14 < lcam_stq_idx_1 ^ _forwarded_is_older_T_117 ^ lcam_stq_idx_1 < ldq_14_bits_youngest_stq_idx);
  wire        _GEN_641 = do_ld_search_1 & ldq_14_valid & ldq_14_bits_addr_valid & ~ldq_14_bits_addr_is_virtual & dword_addr_matches_14_1 & (|_mask_overlap_T_58);
  wire        searcher_is_older_29 = lcam_ldq_idx_1 < 5'hE ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_119;
  wire        _GEN_642 = lcam_ldq_idx_1 != 5'hE;
  reg         older_nacked_REG_29;
  wire        _GEN_643 = ~_GEN_627 | nacking_loads_14 | older_nacked_REG_29;
  reg         io_dmem_s1_kill_1_REG_14;
  wire        _GEN_644 = _GEN_641 & searcher_is_older_29 & _GEN_632 & ldq_14_bits_observed;
  wire        failed_loads_14 = _GEN_637 ? _GEN_90244 : _GEN_639 ? _GEN_640 | _GEN_90244 : _GEN_644 | _GEN_90244;
  wire        _GEN_645 = _GEN_637 | _GEN_639;
  wire        _GEN_646 = _GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643);
  wire [14:0] _l_mask_mask_T_227 = 15'h1 << ldq_15_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_231 = 15'h3 << {12'h0, ldq_15_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_15_bits_uop_mem_size)
      2'b00:
        casez_tmp_127 = _l_mask_mask_T_227[7:0];
      2'b01:
        casez_tmp_127 = _l_mask_mask_T_231[7:0];
      2'b10:
        casez_tmp_127 = ldq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_127 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_15_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'hF;
  wire        l_forwarders_15_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'hF;
  wire        l_is_forwarding_15 = l_forwarders_15_0 | l_forwarders_15_1;
  wire [4:0]  l_forward_stq_idx_15 = l_is_forwarding_15 ? (l_forwarders_15_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_15_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_15_bits_forward_stq_idx;
  wire        block_addr_matches_15_1 = lcam_addr_1[39:6] == ldq_15_bits_addr_bits[39:6];
  wire        dword_addr_matches_15_0 = lcam_addr_0[39:6] == ldq_15_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_15_bits_addr_bits[5:3];
  wire        dword_addr_matches_15_1 = block_addr_matches_15_1 & lcam_addr_1[5:3] == ldq_15_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_60 = casez_tmp_127 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_62 = casez_tmp_127 & casez_tmp_109;
  wire        _GEN_647 = ldq_15_bits_executed | ldq_15_bits_succeeded;
  wire        _GEN_648 = _GEN_647 | l_is_forwarding_15;
  wire [31:0] _GEN_649 = ldq_15_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_650 = do_st_search_0 & ldq_15_valid & ldq_15_bits_addr_valid & _GEN_648 & ~ldq_15_bits_addr_is_virtual & _GEN_649[0] & dword_addr_matches_15_0 & (|_mask_overlap_T_60);
  wire        _forwarded_is_older_T_125 = l_forward_stq_idx_15 < ldq_15_bits_youngest_stq_idx;
  wire        _GEN_90566 = ~ldq_15_bits_forward_std_val | l_forward_stq_idx_15 != lcam_stq_idx_0 & (l_forward_stq_idx_15 < lcam_stq_idx_0 ^ _forwarded_is_older_T_125 ^ lcam_stq_idx_0 < ldq_15_bits_youngest_stq_idx);
  wire        _GEN_651 = _do_ld_search_T_2 & ldq_15_valid & ldq_15_bits_addr_valid & ~ldq_15_bits_addr_is_virtual & dword_addr_matches_15_0 & (|_mask_overlap_T_60);
  wire        searcher_is_older_30 = lcam_ldq_idx_0 < 5'hF ^ _searcher_is_older_T_249 ^ ldq_head[4];
  wire        _GEN_652 = _GEN_648 & ~s1_executing_loads_15;
  wire        _GEN_90568 = _GEN_652 & ldq_15_bits_observed;
  wire        _GEN_653 = lcam_ldq_idx_0 != 5'hF;
  reg         older_nacked_REG_30;
  wire        _GEN_116710 = io_dmem_nack_0_bits_uop_ldq_idx == 5'hF;
  wire        _GEN_654 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'hF;
  wire        nacking_loads_15 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_654 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116710;
  wire        _GEN_655 = ~_GEN_647 | nacking_loads_15 | older_nacked_REG_30;
  reg         io_dmem_s1_kill_0_REG_15;
  wire        _GEN_90742 = _GEN_650 ? _GEN_90566 : _GEN_651 & searcher_is_older_30 & _GEN_90568;
  wire        _GEN_656 = _GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655);
  wire        _GEN_657 = fired_release_1 & ldq_15_valid & ldq_15_bits_addr_valid & block_addr_matches_15_1;
  wire [31:0] _GEN_658 = ldq_15_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_659 = do_st_search_1 & ldq_15_valid & ldq_15_bits_addr_valid & _GEN_648 & ~ldq_15_bits_addr_is_virtual & _GEN_658[0] & dword_addr_matches_15_1 & (|_mask_overlap_T_62);
  wire        _GEN_660 = ~ldq_15_bits_forward_std_val | l_forward_stq_idx_15 != lcam_stq_idx_1 & (l_forward_stq_idx_15 < lcam_stq_idx_1 ^ _forwarded_is_older_T_125 ^ lcam_stq_idx_1 < ldq_15_bits_youngest_stq_idx);
  wire        _GEN_661 = do_ld_search_1 & ldq_15_valid & ldq_15_bits_addr_valid & ~ldq_15_bits_addr_is_virtual & dword_addr_matches_15_1 & (|_mask_overlap_T_62);
  wire        searcher_is_older_31 = lcam_ldq_idx_1 < 5'hF ^ _searcher_is_older_T_253 ^ ldq_head[4];
  wire        _GEN_662 = lcam_ldq_idx_1 != 5'hF;
  reg         older_nacked_REG_31;
  wire        _GEN_663 = ~_GEN_647 | nacking_loads_15 | older_nacked_REG_31;
  reg         io_dmem_s1_kill_1_REG_15;
  wire        _GEN_664 = _GEN_661 & searcher_is_older_31 & _GEN_652 & ldq_15_bits_observed;
  wire        failed_loads_15 = _GEN_657 ? _GEN_90742 : _GEN_659 ? _GEN_660 | _GEN_90742 : _GEN_664 | _GEN_90742;
  wire        _GEN_665 = _GEN_657 | _GEN_659;
  wire        _GEN_666 = _GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663);
  wire [14:0] _l_mask_mask_T_242 = 15'h1 << ldq_16_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_246 = 15'h3 << {12'h0, ldq_16_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_16_bits_uop_mem_size)
      2'b00:
        casez_tmp_128 = _l_mask_mask_T_242[7:0];
      2'b01:
        casez_tmp_128 = _l_mask_mask_T_246[7:0];
      2'b10:
        casez_tmp_128 = ldq_16_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_128 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_16_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h10;
  wire        l_forwarders_16_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h10;
  wire        l_is_forwarding_16 = l_forwarders_16_0 | l_forwarders_16_1;
  wire [4:0]  l_forward_stq_idx_16 = l_is_forwarding_16 ? (l_forwarders_16_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_16_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_16_bits_forward_stq_idx;
  wire        block_addr_matches_16_1 = lcam_addr_1[39:6] == ldq_16_bits_addr_bits[39:6];
  wire        dword_addr_matches_16_0 = lcam_addr_0[39:6] == ldq_16_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_16_bits_addr_bits[5:3];
  wire        dword_addr_matches_16_1 = block_addr_matches_16_1 & lcam_addr_1[5:3] == ldq_16_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_64 = casez_tmp_128 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_66 = casez_tmp_128 & casez_tmp_109;
  wire        _GEN_667 = ldq_16_bits_executed | ldq_16_bits_succeeded;
  wire        _GEN_668 = _GEN_667 | l_is_forwarding_16;
  wire [31:0] _GEN_669 = ldq_16_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_670 = do_st_search_0 & ldq_16_valid & ldq_16_bits_addr_valid & _GEN_668 & ~ldq_16_bits_addr_is_virtual & _GEN_669[0] & dword_addr_matches_16_0 & (|_mask_overlap_T_64);
  wire        _forwarded_is_older_T_133 = l_forward_stq_idx_16 < ldq_16_bits_youngest_stq_idx;
  wire        _GEN_91064 = ~ldq_16_bits_forward_std_val | l_forward_stq_idx_16 != lcam_stq_idx_0 & (l_forward_stq_idx_16 < lcam_stq_idx_0 ^ _forwarded_is_older_T_133 ^ lcam_stq_idx_0 < ldq_16_bits_youngest_stq_idx);
  wire        _GEN_671 = _do_ld_search_T_2 & ldq_16_valid & ldq_16_bits_addr_valid & ~ldq_16_bits_addr_is_virtual & dword_addr_matches_16_0 & (|_mask_overlap_T_64);
  wire        _searcher_is_older_T_135 = ldq_head > 5'h10;
  wire        searcher_is_older_32 = lcam_ldq_idx_0[4] ^ _searcher_is_older_T_249 ^ ~_searcher_is_older_T_135;
  wire        _GEN_672 = _GEN_668 & ~s1_executing_loads_16;
  wire        _GEN_91066 = _GEN_672 & ldq_16_bits_observed;
  wire        _GEN_673 = lcam_ldq_idx_0 != 5'h10;
  reg         older_nacked_REG_32;
  wire        _GEN_116711 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h10;
  wire        _GEN_674 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h10;
  wire        nacking_loads_16 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_674 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116711;
  wire        _GEN_675 = ~_GEN_667 | nacking_loads_16 | older_nacked_REG_32;
  reg         io_dmem_s1_kill_0_REG_16;
  wire        _GEN_91240 = _GEN_670 ? _GEN_91064 : _GEN_671 & searcher_is_older_32 & _GEN_91066;
  wire        _GEN_676 = _GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675);
  wire        _GEN_677 = fired_release_1 & ldq_16_valid & ldq_16_bits_addr_valid & block_addr_matches_16_1;
  wire [31:0] _GEN_678 = ldq_16_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_679 = do_st_search_1 & ldq_16_valid & ldq_16_bits_addr_valid & _GEN_668 & ~ldq_16_bits_addr_is_virtual & _GEN_678[0] & dword_addr_matches_16_1 & (|_mask_overlap_T_66);
  wire        _GEN_680 = ~ldq_16_bits_forward_std_val | l_forward_stq_idx_16 != lcam_stq_idx_1 & (l_forward_stq_idx_16 < lcam_stq_idx_1 ^ _forwarded_is_older_T_133 ^ lcam_stq_idx_1 < ldq_16_bits_youngest_stq_idx);
  wire        _GEN_681 = do_ld_search_1 & ldq_16_valid & ldq_16_bits_addr_valid & ~ldq_16_bits_addr_is_virtual & dword_addr_matches_16_1 & (|_mask_overlap_T_66);
  wire        searcher_is_older_33 = lcam_ldq_idx_1[4] ^ _searcher_is_older_T_253 ^ ~_searcher_is_older_T_135;
  wire        _GEN_682 = lcam_ldq_idx_1 != 5'h10;
  reg         older_nacked_REG_33;
  wire        _GEN_683 = ~_GEN_667 | nacking_loads_16 | older_nacked_REG_33;
  reg         io_dmem_s1_kill_1_REG_16;
  wire        _GEN_684 = _GEN_681 & searcher_is_older_33 & _GEN_672 & ldq_16_bits_observed;
  wire        failed_loads_16 = _GEN_677 ? _GEN_91240 : _GEN_679 ? _GEN_680 | _GEN_91240 : _GEN_684 | _GEN_91240;
  wire        _GEN_685 = _GEN_677 | _GEN_679;
  wire        _GEN_686 = _GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683);
  wire [14:0] _l_mask_mask_T_257 = 15'h1 << ldq_17_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_261 = 15'h3 << {12'h0, ldq_17_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_17_bits_uop_mem_size)
      2'b00:
        casez_tmp_129 = _l_mask_mask_T_257[7:0];
      2'b01:
        casez_tmp_129 = _l_mask_mask_T_261[7:0];
      2'b10:
        casez_tmp_129 = ldq_17_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_129 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_17_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h11;
  wire        l_forwarders_17_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h11;
  wire        l_is_forwarding_17 = l_forwarders_17_0 | l_forwarders_17_1;
  wire [4:0]  l_forward_stq_idx_17 = l_is_forwarding_17 ? (l_forwarders_17_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_17_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_17_bits_forward_stq_idx;
  wire        block_addr_matches_17_1 = lcam_addr_1[39:6] == ldq_17_bits_addr_bits[39:6];
  wire        dword_addr_matches_17_0 = lcam_addr_0[39:6] == ldq_17_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_17_bits_addr_bits[5:3];
  wire        dword_addr_matches_17_1 = block_addr_matches_17_1 & lcam_addr_1[5:3] == ldq_17_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_68 = casez_tmp_129 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_70 = casez_tmp_129 & casez_tmp_109;
  wire        _GEN_687 = ldq_17_bits_executed | ldq_17_bits_succeeded;
  wire        _GEN_688 = _GEN_687 | l_is_forwarding_17;
  wire [31:0] _GEN_689 = ldq_17_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_690 = do_st_search_0 & ldq_17_valid & ldq_17_bits_addr_valid & _GEN_688 & ~ldq_17_bits_addr_is_virtual & _GEN_689[0] & dword_addr_matches_17_0 & (|_mask_overlap_T_68);
  wire        _forwarded_is_older_T_141 = l_forward_stq_idx_17 < ldq_17_bits_youngest_stq_idx;
  wire        _GEN_91562 = ~ldq_17_bits_forward_std_val | l_forward_stq_idx_17 != lcam_stq_idx_0 & (l_forward_stq_idx_17 < lcam_stq_idx_0 ^ _forwarded_is_older_T_141 ^ lcam_stq_idx_0 < ldq_17_bits_youngest_stq_idx);
  wire        _GEN_691 = _do_ld_search_T_2 & ldq_17_valid & ldq_17_bits_addr_valid & ~ldq_17_bits_addr_is_virtual & dword_addr_matches_17_0 & (|_mask_overlap_T_68);
  wire        _searcher_is_older_T_143 = ldq_head > 5'h11;
  wire        searcher_is_older_34 = lcam_ldq_idx_0 < 5'h11 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_143;
  wire        _GEN_692 = _GEN_688 & ~s1_executing_loads_17;
  wire        _GEN_91564 = _GEN_692 & ldq_17_bits_observed;
  wire        _GEN_693 = lcam_ldq_idx_0 != 5'h11;
  reg         older_nacked_REG_34;
  wire        _GEN_116712 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h11;
  wire        _GEN_694 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h11;
  wire        nacking_loads_17 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_694 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116712;
  wire        _GEN_695 = ~_GEN_687 | nacking_loads_17 | older_nacked_REG_34;
  reg         io_dmem_s1_kill_0_REG_17;
  wire        _GEN_91738 = _GEN_690 ? _GEN_91562 : _GEN_691 & searcher_is_older_34 & _GEN_91564;
  wire        _GEN_696 = _GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695);
  wire        _GEN_697 = fired_release_1 & ldq_17_valid & ldq_17_bits_addr_valid & block_addr_matches_17_1;
  wire [31:0] _GEN_698 = ldq_17_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_699 = do_st_search_1 & ldq_17_valid & ldq_17_bits_addr_valid & _GEN_688 & ~ldq_17_bits_addr_is_virtual & _GEN_698[0] & dword_addr_matches_17_1 & (|_mask_overlap_T_70);
  wire        _GEN_700 = ~ldq_17_bits_forward_std_val | l_forward_stq_idx_17 != lcam_stq_idx_1 & (l_forward_stq_idx_17 < lcam_stq_idx_1 ^ _forwarded_is_older_T_141 ^ lcam_stq_idx_1 < ldq_17_bits_youngest_stq_idx);
  wire        _GEN_701 = do_ld_search_1 & ldq_17_valid & ldq_17_bits_addr_valid & ~ldq_17_bits_addr_is_virtual & dword_addr_matches_17_1 & (|_mask_overlap_T_70);
  wire        searcher_is_older_35 = lcam_ldq_idx_1 < 5'h11 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_143;
  wire        _GEN_702 = lcam_ldq_idx_1 != 5'h11;
  reg         older_nacked_REG_35;
  wire        _GEN_703 = ~_GEN_687 | nacking_loads_17 | older_nacked_REG_35;
  reg         io_dmem_s1_kill_1_REG_17;
  wire        _GEN_704 = _GEN_701 & searcher_is_older_35 & _GEN_692 & ldq_17_bits_observed;
  wire        failed_loads_17 = _GEN_697 ? _GEN_91738 : _GEN_699 ? _GEN_700 | _GEN_91738 : _GEN_704 | _GEN_91738;
  wire        _GEN_705 = _GEN_697 | _GEN_699;
  wire        _GEN_706 = _GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703);
  wire [14:0] _l_mask_mask_T_272 = 15'h1 << ldq_18_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_276 = 15'h3 << {12'h0, ldq_18_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_18_bits_uop_mem_size)
      2'b00:
        casez_tmp_130 = _l_mask_mask_T_272[7:0];
      2'b01:
        casez_tmp_130 = _l_mask_mask_T_276[7:0];
      2'b10:
        casez_tmp_130 = ldq_18_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_130 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_18_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h12;
  wire        l_forwarders_18_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h12;
  wire        l_is_forwarding_18 = l_forwarders_18_0 | l_forwarders_18_1;
  wire [4:0]  l_forward_stq_idx_18 = l_is_forwarding_18 ? (l_forwarders_18_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_18_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_18_bits_forward_stq_idx;
  wire        block_addr_matches_18_1 = lcam_addr_1[39:6] == ldq_18_bits_addr_bits[39:6];
  wire        dword_addr_matches_18_0 = lcam_addr_0[39:6] == ldq_18_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_18_bits_addr_bits[5:3];
  wire        dword_addr_matches_18_1 = block_addr_matches_18_1 & lcam_addr_1[5:3] == ldq_18_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_72 = casez_tmp_130 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_74 = casez_tmp_130 & casez_tmp_109;
  wire        _GEN_707 = ldq_18_bits_executed | ldq_18_bits_succeeded;
  wire        _GEN_708 = _GEN_707 | l_is_forwarding_18;
  wire [31:0] _GEN_709 = ldq_18_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_710 = do_st_search_0 & ldq_18_valid & ldq_18_bits_addr_valid & _GEN_708 & ~ldq_18_bits_addr_is_virtual & _GEN_709[0] & dword_addr_matches_18_0 & (|_mask_overlap_T_72);
  wire        _forwarded_is_older_T_149 = l_forward_stq_idx_18 < ldq_18_bits_youngest_stq_idx;
  wire        _GEN_92060 = ~ldq_18_bits_forward_std_val | l_forward_stq_idx_18 != lcam_stq_idx_0 & (l_forward_stq_idx_18 < lcam_stq_idx_0 ^ _forwarded_is_older_T_149 ^ lcam_stq_idx_0 < ldq_18_bits_youngest_stq_idx);
  wire        _GEN_711 = _do_ld_search_T_2 & ldq_18_valid & ldq_18_bits_addr_valid & ~ldq_18_bits_addr_is_virtual & dword_addr_matches_18_0 & (|_mask_overlap_T_72);
  wire        _searcher_is_older_T_151 = ldq_head > 5'h12;
  wire        searcher_is_older_36 = lcam_ldq_idx_0 < 5'h12 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_151;
  wire        _GEN_712 = _GEN_708 & ~s1_executing_loads_18;
  wire        _GEN_92062 = _GEN_712 & ldq_18_bits_observed;
  wire        _GEN_713 = lcam_ldq_idx_0 != 5'h12;
  reg         older_nacked_REG_36;
  wire        _GEN_116713 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h12;
  wire        _GEN_714 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h12;
  wire        nacking_loads_18 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_714 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116713;
  wire        _GEN_715 = ~_GEN_707 | nacking_loads_18 | older_nacked_REG_36;
  reg         io_dmem_s1_kill_0_REG_18;
  wire        _GEN_92236 = _GEN_710 ? _GEN_92060 : _GEN_711 & searcher_is_older_36 & _GEN_92062;
  wire        _GEN_716 = _GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715);
  wire        _GEN_717 = fired_release_1 & ldq_18_valid & ldq_18_bits_addr_valid & block_addr_matches_18_1;
  wire [31:0] _GEN_718 = ldq_18_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_719 = do_st_search_1 & ldq_18_valid & ldq_18_bits_addr_valid & _GEN_708 & ~ldq_18_bits_addr_is_virtual & _GEN_718[0] & dword_addr_matches_18_1 & (|_mask_overlap_T_74);
  wire        _GEN_720 = ~ldq_18_bits_forward_std_val | l_forward_stq_idx_18 != lcam_stq_idx_1 & (l_forward_stq_idx_18 < lcam_stq_idx_1 ^ _forwarded_is_older_T_149 ^ lcam_stq_idx_1 < ldq_18_bits_youngest_stq_idx);
  wire        _GEN_721 = do_ld_search_1 & ldq_18_valid & ldq_18_bits_addr_valid & ~ldq_18_bits_addr_is_virtual & dword_addr_matches_18_1 & (|_mask_overlap_T_74);
  wire        searcher_is_older_37 = lcam_ldq_idx_1 < 5'h12 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_151;
  wire        _GEN_722 = lcam_ldq_idx_1 != 5'h12;
  reg         older_nacked_REG_37;
  wire        _GEN_723 = ~_GEN_707 | nacking_loads_18 | older_nacked_REG_37;
  reg         io_dmem_s1_kill_1_REG_18;
  wire        _GEN_724 = _GEN_721 & searcher_is_older_37 & _GEN_712 & ldq_18_bits_observed;
  wire        failed_loads_18 = _GEN_717 ? _GEN_92236 : _GEN_719 ? _GEN_720 | _GEN_92236 : _GEN_724 | _GEN_92236;
  wire        _GEN_725 = _GEN_717 | _GEN_719;
  wire        _GEN_726 = _GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723);
  wire [14:0] _l_mask_mask_T_287 = 15'h1 << ldq_19_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_291 = 15'h3 << {12'h0, ldq_19_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_19_bits_uop_mem_size)
      2'b00:
        casez_tmp_131 = _l_mask_mask_T_287[7:0];
      2'b01:
        casez_tmp_131 = _l_mask_mask_T_291[7:0];
      2'b10:
        casez_tmp_131 = ldq_19_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_131 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_19_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h13;
  wire        l_forwarders_19_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h13;
  wire        l_is_forwarding_19 = l_forwarders_19_0 | l_forwarders_19_1;
  wire [4:0]  l_forward_stq_idx_19 = l_is_forwarding_19 ? (l_forwarders_19_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_19_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_19_bits_forward_stq_idx;
  wire        block_addr_matches_19_1 = lcam_addr_1[39:6] == ldq_19_bits_addr_bits[39:6];
  wire        dword_addr_matches_19_0 = lcam_addr_0[39:6] == ldq_19_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_19_bits_addr_bits[5:3];
  wire        dword_addr_matches_19_1 = block_addr_matches_19_1 & lcam_addr_1[5:3] == ldq_19_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_76 = casez_tmp_131 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_78 = casez_tmp_131 & casez_tmp_109;
  wire        _GEN_727 = ldq_19_bits_executed | ldq_19_bits_succeeded;
  wire        _GEN_728 = _GEN_727 | l_is_forwarding_19;
  wire [31:0] _GEN_729 = ldq_19_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_730 = do_st_search_0 & ldq_19_valid & ldq_19_bits_addr_valid & _GEN_728 & ~ldq_19_bits_addr_is_virtual & _GEN_729[0] & dword_addr_matches_19_0 & (|_mask_overlap_T_76);
  wire        _forwarded_is_older_T_157 = l_forward_stq_idx_19 < ldq_19_bits_youngest_stq_idx;
  wire        _GEN_92558 = ~ldq_19_bits_forward_std_val | l_forward_stq_idx_19 != lcam_stq_idx_0 & (l_forward_stq_idx_19 < lcam_stq_idx_0 ^ _forwarded_is_older_T_157 ^ lcam_stq_idx_0 < ldq_19_bits_youngest_stq_idx);
  wire        _GEN_731 = _do_ld_search_T_2 & ldq_19_valid & ldq_19_bits_addr_valid & ~ldq_19_bits_addr_is_virtual & dword_addr_matches_19_0 & (|_mask_overlap_T_76);
  wire        _searcher_is_older_T_159 = ldq_head > 5'h13;
  wire        searcher_is_older_38 = lcam_ldq_idx_0 < 5'h13 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_159;
  wire        _GEN_732 = _GEN_728 & ~s1_executing_loads_19;
  wire        _GEN_92560 = _GEN_732 & ldq_19_bits_observed;
  wire        _GEN_733 = lcam_ldq_idx_0 != 5'h13;
  reg         older_nacked_REG_38;
  wire        _GEN_116714 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h13;
  wire        _GEN_734 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h13;
  wire        nacking_loads_19 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_734 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116714;
  wire        _GEN_735 = ~_GEN_727 | nacking_loads_19 | older_nacked_REG_38;
  reg         io_dmem_s1_kill_0_REG_19;
  wire        _GEN_92734 = _GEN_730 ? _GEN_92558 : _GEN_731 & searcher_is_older_38 & _GEN_92560;
  wire        _GEN_736 = _GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735);
  wire        _GEN_737 = fired_release_1 & ldq_19_valid & ldq_19_bits_addr_valid & block_addr_matches_19_1;
  wire [31:0] _GEN_738 = ldq_19_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_739 = do_st_search_1 & ldq_19_valid & ldq_19_bits_addr_valid & _GEN_728 & ~ldq_19_bits_addr_is_virtual & _GEN_738[0] & dword_addr_matches_19_1 & (|_mask_overlap_T_78);
  wire        _GEN_740 = ~ldq_19_bits_forward_std_val | l_forward_stq_idx_19 != lcam_stq_idx_1 & (l_forward_stq_idx_19 < lcam_stq_idx_1 ^ _forwarded_is_older_T_157 ^ lcam_stq_idx_1 < ldq_19_bits_youngest_stq_idx);
  wire        _GEN_741 = do_ld_search_1 & ldq_19_valid & ldq_19_bits_addr_valid & ~ldq_19_bits_addr_is_virtual & dword_addr_matches_19_1 & (|_mask_overlap_T_78);
  wire        searcher_is_older_39 = lcam_ldq_idx_1 < 5'h13 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_159;
  wire        _GEN_742 = lcam_ldq_idx_1 != 5'h13;
  reg         older_nacked_REG_39;
  wire        _GEN_743 = ~_GEN_727 | nacking_loads_19 | older_nacked_REG_39;
  reg         io_dmem_s1_kill_1_REG_19;
  wire        _GEN_744 = _GEN_741 & searcher_is_older_39 & _GEN_732 & ldq_19_bits_observed;
  wire        failed_loads_19 = _GEN_737 ? _GEN_92734 : _GEN_739 ? _GEN_740 | _GEN_92734 : _GEN_744 | _GEN_92734;
  wire        _GEN_745 = _GEN_737 | _GEN_739;
  wire        _GEN_746 = _GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743);
  wire [14:0] _l_mask_mask_T_302 = 15'h1 << ldq_20_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_306 = 15'h3 << {12'h0, ldq_20_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_20_bits_uop_mem_size)
      2'b00:
        casez_tmp_132 = _l_mask_mask_T_302[7:0];
      2'b01:
        casez_tmp_132 = _l_mask_mask_T_306[7:0];
      2'b10:
        casez_tmp_132 = ldq_20_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_132 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_20_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h14;
  wire        l_forwarders_20_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h14;
  wire        l_is_forwarding_20 = l_forwarders_20_0 | l_forwarders_20_1;
  wire [4:0]  l_forward_stq_idx_20 = l_is_forwarding_20 ? (l_forwarders_20_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_20_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_20_bits_forward_stq_idx;
  wire        block_addr_matches_20_1 = lcam_addr_1[39:6] == ldq_20_bits_addr_bits[39:6];
  wire        dword_addr_matches_20_0 = lcam_addr_0[39:6] == ldq_20_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_20_bits_addr_bits[5:3];
  wire        dword_addr_matches_20_1 = block_addr_matches_20_1 & lcam_addr_1[5:3] == ldq_20_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_80 = casez_tmp_132 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_82 = casez_tmp_132 & casez_tmp_109;
  wire        _GEN_747 = ldq_20_bits_executed | ldq_20_bits_succeeded;
  wire        _GEN_748 = _GEN_747 | l_is_forwarding_20;
  wire [31:0] _GEN_749 = ldq_20_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_750 = do_st_search_0 & ldq_20_valid & ldq_20_bits_addr_valid & _GEN_748 & ~ldq_20_bits_addr_is_virtual & _GEN_749[0] & dword_addr_matches_20_0 & (|_mask_overlap_T_80);
  wire        _forwarded_is_older_T_165 = l_forward_stq_idx_20 < ldq_20_bits_youngest_stq_idx;
  wire        _GEN_93056 = ~ldq_20_bits_forward_std_val | l_forward_stq_idx_20 != lcam_stq_idx_0 & (l_forward_stq_idx_20 < lcam_stq_idx_0 ^ _forwarded_is_older_T_165 ^ lcam_stq_idx_0 < ldq_20_bits_youngest_stq_idx);
  wire        _GEN_751 = _do_ld_search_T_2 & ldq_20_valid & ldq_20_bits_addr_valid & ~ldq_20_bits_addr_is_virtual & dword_addr_matches_20_0 & (|_mask_overlap_T_80);
  wire        _searcher_is_older_T_167 = ldq_head > 5'h14;
  wire        searcher_is_older_40 = lcam_ldq_idx_0 < 5'h14 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_167;
  wire        _GEN_752 = _GEN_748 & ~s1_executing_loads_20;
  wire        _GEN_93058 = _GEN_752 & ldq_20_bits_observed;
  wire        _GEN_753 = lcam_ldq_idx_0 != 5'h14;
  reg         older_nacked_REG_40;
  wire        _GEN_116715 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h14;
  wire        _GEN_754 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h14;
  wire        nacking_loads_20 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_754 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116715;
  wire        _GEN_755 = ~_GEN_747 | nacking_loads_20 | older_nacked_REG_40;
  reg         io_dmem_s1_kill_0_REG_20;
  wire        _GEN_93232 = _GEN_750 ? _GEN_93056 : _GEN_751 & searcher_is_older_40 & _GEN_93058;
  wire        _GEN_756 = _GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755);
  wire        _GEN_757 = fired_release_1 & ldq_20_valid & ldq_20_bits_addr_valid & block_addr_matches_20_1;
  wire [31:0] _GEN_758 = ldq_20_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_759 = do_st_search_1 & ldq_20_valid & ldq_20_bits_addr_valid & _GEN_748 & ~ldq_20_bits_addr_is_virtual & _GEN_758[0] & dword_addr_matches_20_1 & (|_mask_overlap_T_82);
  wire        _GEN_760 = ~ldq_20_bits_forward_std_val | l_forward_stq_idx_20 != lcam_stq_idx_1 & (l_forward_stq_idx_20 < lcam_stq_idx_1 ^ _forwarded_is_older_T_165 ^ lcam_stq_idx_1 < ldq_20_bits_youngest_stq_idx);
  wire        _GEN_761 = do_ld_search_1 & ldq_20_valid & ldq_20_bits_addr_valid & ~ldq_20_bits_addr_is_virtual & dword_addr_matches_20_1 & (|_mask_overlap_T_82);
  wire        searcher_is_older_41 = lcam_ldq_idx_1 < 5'h14 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_167;
  wire        _GEN_762 = lcam_ldq_idx_1 != 5'h14;
  reg         older_nacked_REG_41;
  wire        _GEN_763 = ~_GEN_747 | nacking_loads_20 | older_nacked_REG_41;
  reg         io_dmem_s1_kill_1_REG_20;
  wire        _GEN_764 = _GEN_761 & searcher_is_older_41 & _GEN_752 & ldq_20_bits_observed;
  wire        failed_loads_20 = _GEN_757 ? _GEN_93232 : _GEN_759 ? _GEN_760 | _GEN_93232 : _GEN_764 | _GEN_93232;
  wire        _GEN_765 = _GEN_757 | _GEN_759;
  wire        _GEN_766 = _GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763);
  wire [14:0] _l_mask_mask_T_317 = 15'h1 << ldq_21_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_321 = 15'h3 << {12'h0, ldq_21_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_21_bits_uop_mem_size)
      2'b00:
        casez_tmp_133 = _l_mask_mask_T_317[7:0];
      2'b01:
        casez_tmp_133 = _l_mask_mask_T_321[7:0];
      2'b10:
        casez_tmp_133 = ldq_21_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_133 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_21_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h15;
  wire        l_forwarders_21_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h15;
  wire        l_is_forwarding_21 = l_forwarders_21_0 | l_forwarders_21_1;
  wire [4:0]  l_forward_stq_idx_21 = l_is_forwarding_21 ? (l_forwarders_21_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_21_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_21_bits_forward_stq_idx;
  wire        block_addr_matches_21_1 = lcam_addr_1[39:6] == ldq_21_bits_addr_bits[39:6];
  wire        dword_addr_matches_21_0 = lcam_addr_0[39:6] == ldq_21_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_21_bits_addr_bits[5:3];
  wire        dword_addr_matches_21_1 = block_addr_matches_21_1 & lcam_addr_1[5:3] == ldq_21_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_84 = casez_tmp_133 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_86 = casez_tmp_133 & casez_tmp_109;
  wire        _GEN_767 = ldq_21_bits_executed | ldq_21_bits_succeeded;
  wire        _GEN_768 = _GEN_767 | l_is_forwarding_21;
  wire [31:0] _GEN_769 = ldq_21_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_770 = do_st_search_0 & ldq_21_valid & ldq_21_bits_addr_valid & _GEN_768 & ~ldq_21_bits_addr_is_virtual & _GEN_769[0] & dword_addr_matches_21_0 & (|_mask_overlap_T_84);
  wire        _forwarded_is_older_T_173 = l_forward_stq_idx_21 < ldq_21_bits_youngest_stq_idx;
  wire        _GEN_93554 = ~ldq_21_bits_forward_std_val | l_forward_stq_idx_21 != lcam_stq_idx_0 & (l_forward_stq_idx_21 < lcam_stq_idx_0 ^ _forwarded_is_older_T_173 ^ lcam_stq_idx_0 < ldq_21_bits_youngest_stq_idx);
  wire        _GEN_771 = _do_ld_search_T_2 & ldq_21_valid & ldq_21_bits_addr_valid & ~ldq_21_bits_addr_is_virtual & dword_addr_matches_21_0 & (|_mask_overlap_T_84);
  wire        _searcher_is_older_T_175 = ldq_head > 5'h15;
  wire        searcher_is_older_42 = lcam_ldq_idx_0 < 5'h15 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_175;
  wire        _GEN_772 = _GEN_768 & ~s1_executing_loads_21;
  wire        _GEN_93556 = _GEN_772 & ldq_21_bits_observed;
  wire        _GEN_773 = lcam_ldq_idx_0 != 5'h15;
  reg         older_nacked_REG_42;
  wire        _GEN_116716 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h15;
  wire        _GEN_774 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h15;
  wire        nacking_loads_21 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_774 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116716;
  wire        _GEN_775 = ~_GEN_767 | nacking_loads_21 | older_nacked_REG_42;
  reg         io_dmem_s1_kill_0_REG_21;
  wire        _GEN_93730 = _GEN_770 ? _GEN_93554 : _GEN_771 & searcher_is_older_42 & _GEN_93556;
  wire        _GEN_776 = _GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775);
  wire        _GEN_777 = fired_release_1 & ldq_21_valid & ldq_21_bits_addr_valid & block_addr_matches_21_1;
  wire [31:0] _GEN_778 = ldq_21_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_779 = do_st_search_1 & ldq_21_valid & ldq_21_bits_addr_valid & _GEN_768 & ~ldq_21_bits_addr_is_virtual & _GEN_778[0] & dword_addr_matches_21_1 & (|_mask_overlap_T_86);
  wire        _GEN_780 = ~ldq_21_bits_forward_std_val | l_forward_stq_idx_21 != lcam_stq_idx_1 & (l_forward_stq_idx_21 < lcam_stq_idx_1 ^ _forwarded_is_older_T_173 ^ lcam_stq_idx_1 < ldq_21_bits_youngest_stq_idx);
  wire        _GEN_781 = do_ld_search_1 & ldq_21_valid & ldq_21_bits_addr_valid & ~ldq_21_bits_addr_is_virtual & dword_addr_matches_21_1 & (|_mask_overlap_T_86);
  wire        searcher_is_older_43 = lcam_ldq_idx_1 < 5'h15 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_175;
  wire        _GEN_782 = lcam_ldq_idx_1 != 5'h15;
  reg         older_nacked_REG_43;
  wire        _GEN_783 = ~_GEN_767 | nacking_loads_21 | older_nacked_REG_43;
  reg         io_dmem_s1_kill_1_REG_21;
  wire        _GEN_784 = _GEN_781 & searcher_is_older_43 & _GEN_772 & ldq_21_bits_observed;
  wire        failed_loads_21 = _GEN_777 ? _GEN_93730 : _GEN_779 ? _GEN_780 | _GEN_93730 : _GEN_784 | _GEN_93730;
  wire        _GEN_785 = _GEN_777 | _GEN_779;
  wire        _GEN_786 = _GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783);
  wire [14:0] _l_mask_mask_T_332 = 15'h1 << ldq_22_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_336 = 15'h3 << {12'h0, ldq_22_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_22_bits_uop_mem_size)
      2'b00:
        casez_tmp_134 = _l_mask_mask_T_332[7:0];
      2'b01:
        casez_tmp_134 = _l_mask_mask_T_336[7:0];
      2'b10:
        casez_tmp_134 = ldq_22_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_134 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_22_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h16;
  wire        l_forwarders_22_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h16;
  wire        l_is_forwarding_22 = l_forwarders_22_0 | l_forwarders_22_1;
  wire [4:0]  l_forward_stq_idx_22 = l_is_forwarding_22 ? (l_forwarders_22_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_22_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_22_bits_forward_stq_idx;
  wire        block_addr_matches_22_1 = lcam_addr_1[39:6] == ldq_22_bits_addr_bits[39:6];
  wire        dword_addr_matches_22_0 = lcam_addr_0[39:6] == ldq_22_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_22_bits_addr_bits[5:3];
  wire        dword_addr_matches_22_1 = block_addr_matches_22_1 & lcam_addr_1[5:3] == ldq_22_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_88 = casez_tmp_134 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_90 = casez_tmp_134 & casez_tmp_109;
  wire        _GEN_787 = ldq_22_bits_executed | ldq_22_bits_succeeded;
  wire        _GEN_788 = _GEN_787 | l_is_forwarding_22;
  wire [31:0] _GEN_789 = ldq_22_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_790 = do_st_search_0 & ldq_22_valid & ldq_22_bits_addr_valid & _GEN_788 & ~ldq_22_bits_addr_is_virtual & _GEN_789[0] & dword_addr_matches_22_0 & (|_mask_overlap_T_88);
  wire        _forwarded_is_older_T_181 = l_forward_stq_idx_22 < ldq_22_bits_youngest_stq_idx;
  wire        _GEN_94052 = ~ldq_22_bits_forward_std_val | l_forward_stq_idx_22 != lcam_stq_idx_0 & (l_forward_stq_idx_22 < lcam_stq_idx_0 ^ _forwarded_is_older_T_181 ^ lcam_stq_idx_0 < ldq_22_bits_youngest_stq_idx);
  wire        _GEN_791 = _do_ld_search_T_2 & ldq_22_valid & ldq_22_bits_addr_valid & ~ldq_22_bits_addr_is_virtual & dword_addr_matches_22_0 & (|_mask_overlap_T_88);
  wire        _searcher_is_older_T_183 = ldq_head > 5'h16;
  wire        searcher_is_older_44 = lcam_ldq_idx_0 < 5'h16 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_183;
  wire        _GEN_792 = _GEN_788 & ~s1_executing_loads_22;
  wire        _GEN_94054 = _GEN_792 & ldq_22_bits_observed;
  wire        _GEN_793 = lcam_ldq_idx_0 != 5'h16;
  reg         older_nacked_REG_44;
  wire        _GEN_116717 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h16;
  wire        _GEN_794 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h16;
  wire        nacking_loads_22 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_794 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116717;
  wire        _GEN_795 = ~_GEN_787 | nacking_loads_22 | older_nacked_REG_44;
  reg         io_dmem_s1_kill_0_REG_22;
  wire        _GEN_94228 = _GEN_790 ? _GEN_94052 : _GEN_791 & searcher_is_older_44 & _GEN_94054;
  wire        _GEN_796 = _GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795);
  wire        _GEN_797 = fired_release_1 & ldq_22_valid & ldq_22_bits_addr_valid & block_addr_matches_22_1;
  wire [31:0] _GEN_798 = ldq_22_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_799 = do_st_search_1 & ldq_22_valid & ldq_22_bits_addr_valid & _GEN_788 & ~ldq_22_bits_addr_is_virtual & _GEN_798[0] & dword_addr_matches_22_1 & (|_mask_overlap_T_90);
  wire        _GEN_800 = ~ldq_22_bits_forward_std_val | l_forward_stq_idx_22 != lcam_stq_idx_1 & (l_forward_stq_idx_22 < lcam_stq_idx_1 ^ _forwarded_is_older_T_181 ^ lcam_stq_idx_1 < ldq_22_bits_youngest_stq_idx);
  wire        _GEN_801 = do_ld_search_1 & ldq_22_valid & ldq_22_bits_addr_valid & ~ldq_22_bits_addr_is_virtual & dword_addr_matches_22_1 & (|_mask_overlap_T_90);
  wire        searcher_is_older_45 = lcam_ldq_idx_1 < 5'h16 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_183;
  wire        _GEN_802 = lcam_ldq_idx_1 != 5'h16;
  reg         older_nacked_REG_45;
  wire        _GEN_803 = ~_GEN_787 | nacking_loads_22 | older_nacked_REG_45;
  reg         io_dmem_s1_kill_1_REG_22;
  wire        _GEN_804 = _GEN_801 & searcher_is_older_45 & _GEN_792 & ldq_22_bits_observed;
  wire        failed_loads_22 = _GEN_797 ? _GEN_94228 : _GEN_799 ? _GEN_800 | _GEN_94228 : _GEN_804 | _GEN_94228;
  wire        _GEN_805 = _GEN_797 | _GEN_799;
  wire        _GEN_806 = _GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803);
  wire [14:0] _l_mask_mask_T_347 = 15'h1 << ldq_23_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_351 = 15'h3 << {12'h0, ldq_23_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_23_bits_uop_mem_size)
      2'b00:
        casez_tmp_135 = _l_mask_mask_T_347[7:0];
      2'b01:
        casez_tmp_135 = _l_mask_mask_T_351[7:0];
      2'b10:
        casez_tmp_135 = ldq_23_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_135 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_23_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h17;
  wire        l_forwarders_23_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h17;
  wire        l_is_forwarding_23 = l_forwarders_23_0 | l_forwarders_23_1;
  wire [4:0]  l_forward_stq_idx_23 = l_is_forwarding_23 ? (l_forwarders_23_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_23_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_23_bits_forward_stq_idx;
  wire        block_addr_matches_23_1 = lcam_addr_1[39:6] == ldq_23_bits_addr_bits[39:6];
  wire        dword_addr_matches_23_0 = lcam_addr_0[39:6] == ldq_23_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_23_bits_addr_bits[5:3];
  wire        dword_addr_matches_23_1 = block_addr_matches_23_1 & lcam_addr_1[5:3] == ldq_23_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_92 = casez_tmp_135 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_94 = casez_tmp_135 & casez_tmp_109;
  wire        _GEN_807 = ldq_23_bits_executed | ldq_23_bits_succeeded;
  wire        _GEN_808 = _GEN_807 | l_is_forwarding_23;
  wire [31:0] _GEN_809 = ldq_23_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_810 = do_st_search_0 & ldq_23_valid & ldq_23_bits_addr_valid & _GEN_808 & ~ldq_23_bits_addr_is_virtual & _GEN_809[0] & dword_addr_matches_23_0 & (|_mask_overlap_T_92);
  wire        _forwarded_is_older_T_189 = l_forward_stq_idx_23 < ldq_23_bits_youngest_stq_idx;
  wire        _GEN_94550 = ~ldq_23_bits_forward_std_val | l_forward_stq_idx_23 != lcam_stq_idx_0 & (l_forward_stq_idx_23 < lcam_stq_idx_0 ^ _forwarded_is_older_T_189 ^ lcam_stq_idx_0 < ldq_23_bits_youngest_stq_idx);
  wire        _GEN_811 = _do_ld_search_T_2 & ldq_23_valid & ldq_23_bits_addr_valid & ~ldq_23_bits_addr_is_virtual & dword_addr_matches_23_0 & (|_mask_overlap_T_92);
  wire        _searcher_is_older_T_191 = ldq_head > 5'h17;
  wire        searcher_is_older_46 = lcam_ldq_idx_0 < 5'h17 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_191;
  wire        _GEN_812 = _GEN_808 & ~s1_executing_loads_23;
  wire        _GEN_94552 = _GEN_812 & ldq_23_bits_observed;
  wire        _GEN_813 = lcam_ldq_idx_0 != 5'h17;
  reg         older_nacked_REG_46;
  wire        _GEN_116718 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h17;
  wire        _GEN_814 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h17;
  wire        nacking_loads_23 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_814 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116718;
  wire        _GEN_815 = ~_GEN_807 | nacking_loads_23 | older_nacked_REG_46;
  reg         io_dmem_s1_kill_0_REG_23;
  wire        _GEN_94726 = _GEN_810 ? _GEN_94550 : _GEN_811 & searcher_is_older_46 & _GEN_94552;
  wire        _GEN_816 = _GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815);
  wire        _GEN_817 = fired_release_1 & ldq_23_valid & ldq_23_bits_addr_valid & block_addr_matches_23_1;
  wire [31:0] _GEN_818 = ldq_23_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_819 = do_st_search_1 & ldq_23_valid & ldq_23_bits_addr_valid & _GEN_808 & ~ldq_23_bits_addr_is_virtual & _GEN_818[0] & dword_addr_matches_23_1 & (|_mask_overlap_T_94);
  wire        _GEN_820 = ~ldq_23_bits_forward_std_val | l_forward_stq_idx_23 != lcam_stq_idx_1 & (l_forward_stq_idx_23 < lcam_stq_idx_1 ^ _forwarded_is_older_T_189 ^ lcam_stq_idx_1 < ldq_23_bits_youngest_stq_idx);
  wire        _GEN_821 = do_ld_search_1 & ldq_23_valid & ldq_23_bits_addr_valid & ~ldq_23_bits_addr_is_virtual & dword_addr_matches_23_1 & (|_mask_overlap_T_94);
  wire        searcher_is_older_47 = lcam_ldq_idx_1 < 5'h17 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_191;
  wire        _GEN_822 = lcam_ldq_idx_1 != 5'h17;
  reg         older_nacked_REG_47;
  wire        _GEN_823 = ~_GEN_807 | nacking_loads_23 | older_nacked_REG_47;
  reg         io_dmem_s1_kill_1_REG_23;
  wire        _GEN_824 = _GEN_821 & searcher_is_older_47 & _GEN_812 & ldq_23_bits_observed;
  wire        failed_loads_23 = _GEN_817 ? _GEN_94726 : _GEN_819 ? _GEN_820 | _GEN_94726 : _GEN_824 | _GEN_94726;
  wire        _GEN_825 = _GEN_817 | _GEN_819;
  wire        _GEN_826 = _GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823);
  wire [14:0] _l_mask_mask_T_362 = 15'h1 << ldq_24_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_366 = 15'h3 << {12'h0, ldq_24_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_24_bits_uop_mem_size)
      2'b00:
        casez_tmp_136 = _l_mask_mask_T_362[7:0];
      2'b01:
        casez_tmp_136 = _l_mask_mask_T_366[7:0];
      2'b10:
        casez_tmp_136 = ldq_24_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_136 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_24_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h18;
  wire        l_forwarders_24_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h18;
  wire        l_is_forwarding_24 = l_forwarders_24_0 | l_forwarders_24_1;
  wire [4:0]  l_forward_stq_idx_24 = l_is_forwarding_24 ? (l_forwarders_24_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_24_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_24_bits_forward_stq_idx;
  wire        block_addr_matches_24_1 = lcam_addr_1[39:6] == ldq_24_bits_addr_bits[39:6];
  wire        dword_addr_matches_24_0 = lcam_addr_0[39:6] == ldq_24_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_24_bits_addr_bits[5:3];
  wire        dword_addr_matches_24_1 = block_addr_matches_24_1 & lcam_addr_1[5:3] == ldq_24_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_96 = casez_tmp_136 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_98 = casez_tmp_136 & casez_tmp_109;
  wire        _GEN_827 = ldq_24_bits_executed | ldq_24_bits_succeeded;
  wire        _GEN_828 = _GEN_827 | l_is_forwarding_24;
  wire [31:0] _GEN_829 = ldq_24_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_830 = do_st_search_0 & ldq_24_valid & ldq_24_bits_addr_valid & _GEN_828 & ~ldq_24_bits_addr_is_virtual & _GEN_829[0] & dword_addr_matches_24_0 & (|_mask_overlap_T_96);
  wire        _forwarded_is_older_T_197 = l_forward_stq_idx_24 < ldq_24_bits_youngest_stq_idx;
  wire        _GEN_95048 = ~ldq_24_bits_forward_std_val | l_forward_stq_idx_24 != lcam_stq_idx_0 & (l_forward_stq_idx_24 < lcam_stq_idx_0 ^ _forwarded_is_older_T_197 ^ lcam_stq_idx_0 < ldq_24_bits_youngest_stq_idx);
  wire        _GEN_831 = _do_ld_search_T_2 & ldq_24_valid & ldq_24_bits_addr_valid & ~ldq_24_bits_addr_is_virtual & dword_addr_matches_24_0 & (|_mask_overlap_T_96);
  wire        _searcher_is_older_T_199 = ldq_head > 5'h18;
  wire        searcher_is_older_48 = lcam_ldq_idx_0[4:3] != 2'h3 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_199;
  wire        _GEN_832 = _GEN_828 & ~s1_executing_loads_24;
  wire        _GEN_95050 = _GEN_832 & ldq_24_bits_observed;
  wire        _GEN_833 = lcam_ldq_idx_0 != 5'h18;
  reg         older_nacked_REG_48;
  wire        _GEN_116719 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h18;
  wire        _GEN_834 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h18;
  wire        nacking_loads_24 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_834 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116719;
  wire        _GEN_835 = ~_GEN_827 | nacking_loads_24 | older_nacked_REG_48;
  reg         io_dmem_s1_kill_0_REG_24;
  wire        _GEN_95224 = _GEN_830 ? _GEN_95048 : _GEN_831 & searcher_is_older_48 & _GEN_95050;
  wire        _GEN_836 = _GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835);
  wire        _GEN_837 = fired_release_1 & ldq_24_valid & ldq_24_bits_addr_valid & block_addr_matches_24_1;
  wire [31:0] _GEN_838 = ldq_24_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_839 = do_st_search_1 & ldq_24_valid & ldq_24_bits_addr_valid & _GEN_828 & ~ldq_24_bits_addr_is_virtual & _GEN_838[0] & dword_addr_matches_24_1 & (|_mask_overlap_T_98);
  wire        _GEN_840 = ~ldq_24_bits_forward_std_val | l_forward_stq_idx_24 != lcam_stq_idx_1 & (l_forward_stq_idx_24 < lcam_stq_idx_1 ^ _forwarded_is_older_T_197 ^ lcam_stq_idx_1 < ldq_24_bits_youngest_stq_idx);
  wire        _GEN_841 = do_ld_search_1 & ldq_24_valid & ldq_24_bits_addr_valid & ~ldq_24_bits_addr_is_virtual & dword_addr_matches_24_1 & (|_mask_overlap_T_98);
  wire        searcher_is_older_49 = lcam_ldq_idx_1[4:3] != 2'h3 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_199;
  wire        _GEN_842 = lcam_ldq_idx_1 != 5'h18;
  reg         older_nacked_REG_49;
  wire        _GEN_843 = ~_GEN_827 | nacking_loads_24 | older_nacked_REG_49;
  reg         io_dmem_s1_kill_1_REG_24;
  wire        _GEN_844 = _GEN_841 & searcher_is_older_49 & _GEN_832 & ldq_24_bits_observed;
  wire        failed_loads_24 = _GEN_837 ? _GEN_95224 : _GEN_839 ? _GEN_840 | _GEN_95224 : _GEN_844 | _GEN_95224;
  wire        _GEN_845 = _GEN_837 | _GEN_839;
  wire        _GEN_846 = _GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843);
  wire [14:0] _l_mask_mask_T_377 = 15'h1 << ldq_25_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_381 = 15'h3 << {12'h0, ldq_25_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_25_bits_uop_mem_size)
      2'b00:
        casez_tmp_137 = _l_mask_mask_T_377[7:0];
      2'b01:
        casez_tmp_137 = _l_mask_mask_T_381[7:0];
      2'b10:
        casez_tmp_137 = ldq_25_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_137 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_25_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h19;
  wire        l_forwarders_25_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h19;
  wire        l_is_forwarding_25 = l_forwarders_25_0 | l_forwarders_25_1;
  wire [4:0]  l_forward_stq_idx_25 = l_is_forwarding_25 ? (l_forwarders_25_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_25_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_25_bits_forward_stq_idx;
  wire        block_addr_matches_25_1 = lcam_addr_1[39:6] == ldq_25_bits_addr_bits[39:6];
  wire        dword_addr_matches_25_0 = lcam_addr_0[39:6] == ldq_25_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_25_bits_addr_bits[5:3];
  wire        dword_addr_matches_25_1 = block_addr_matches_25_1 & lcam_addr_1[5:3] == ldq_25_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_100 = casez_tmp_137 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_102 = casez_tmp_137 & casez_tmp_109;
  wire        _GEN_847 = ldq_25_bits_executed | ldq_25_bits_succeeded;
  wire        _GEN_848 = _GEN_847 | l_is_forwarding_25;
  wire [31:0] _GEN_849 = ldq_25_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_850 = do_st_search_0 & ldq_25_valid & ldq_25_bits_addr_valid & _GEN_848 & ~ldq_25_bits_addr_is_virtual & _GEN_849[0] & dword_addr_matches_25_0 & (|_mask_overlap_T_100);
  wire        _forwarded_is_older_T_205 = l_forward_stq_idx_25 < ldq_25_bits_youngest_stq_idx;
  wire        _GEN_95546 = ~ldq_25_bits_forward_std_val | l_forward_stq_idx_25 != lcam_stq_idx_0 & (l_forward_stq_idx_25 < lcam_stq_idx_0 ^ _forwarded_is_older_T_205 ^ lcam_stq_idx_0 < ldq_25_bits_youngest_stq_idx);
  wire        _GEN_851 = _do_ld_search_T_2 & ldq_25_valid & ldq_25_bits_addr_valid & ~ldq_25_bits_addr_is_virtual & dword_addr_matches_25_0 & (|_mask_overlap_T_100);
  wire        _searcher_is_older_T_207 = ldq_head > 5'h19;
  wire        searcher_is_older_50 = lcam_ldq_idx_0 < 5'h19 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_207;
  wire        _GEN_852 = _GEN_848 & ~s1_executing_loads_25;
  wire        _GEN_95548 = _GEN_852 & ldq_25_bits_observed;
  wire        _GEN_853 = lcam_ldq_idx_0 != 5'h19;
  reg         older_nacked_REG_50;
  wire        _GEN_116720 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h19;
  wire        _GEN_854 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h19;
  wire        nacking_loads_25 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_854 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116720;
  wire        _GEN_855 = ~_GEN_847 | nacking_loads_25 | older_nacked_REG_50;
  reg         io_dmem_s1_kill_0_REG_25;
  wire        _GEN_95722 = _GEN_850 ? _GEN_95546 : _GEN_851 & searcher_is_older_50 & _GEN_95548;
  wire        _GEN_856 = _GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855);
  wire        _GEN_857 = fired_release_1 & ldq_25_valid & ldq_25_bits_addr_valid & block_addr_matches_25_1;
  wire [31:0] _GEN_858 = ldq_25_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_859 = do_st_search_1 & ldq_25_valid & ldq_25_bits_addr_valid & _GEN_848 & ~ldq_25_bits_addr_is_virtual & _GEN_858[0] & dword_addr_matches_25_1 & (|_mask_overlap_T_102);
  wire        _GEN_860 = ~ldq_25_bits_forward_std_val | l_forward_stq_idx_25 != lcam_stq_idx_1 & (l_forward_stq_idx_25 < lcam_stq_idx_1 ^ _forwarded_is_older_T_205 ^ lcam_stq_idx_1 < ldq_25_bits_youngest_stq_idx);
  wire        _GEN_861 = do_ld_search_1 & ldq_25_valid & ldq_25_bits_addr_valid & ~ldq_25_bits_addr_is_virtual & dword_addr_matches_25_1 & (|_mask_overlap_T_102);
  wire        searcher_is_older_51 = lcam_ldq_idx_1 < 5'h19 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_207;
  wire        _GEN_862 = lcam_ldq_idx_1 != 5'h19;
  reg         older_nacked_REG_51;
  wire        _GEN_863 = ~_GEN_847 | nacking_loads_25 | older_nacked_REG_51;
  reg         io_dmem_s1_kill_1_REG_25;
  wire        _GEN_864 = _GEN_861 & searcher_is_older_51 & _GEN_852 & ldq_25_bits_observed;
  wire        failed_loads_25 = _GEN_857 ? _GEN_95722 : _GEN_859 ? _GEN_860 | _GEN_95722 : _GEN_864 | _GEN_95722;
  wire        _GEN_865 = _GEN_857 | _GEN_859;
  wire        _GEN_866 = _GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863);
  wire [14:0] _l_mask_mask_T_392 = 15'h1 << ldq_26_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_396 = 15'h3 << {12'h0, ldq_26_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_26_bits_uop_mem_size)
      2'b00:
        casez_tmp_138 = _l_mask_mask_T_392[7:0];
      2'b01:
        casez_tmp_138 = _l_mask_mask_T_396[7:0];
      2'b10:
        casez_tmp_138 = ldq_26_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_138 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_26_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1A;
  wire        l_forwarders_26_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1A;
  wire        l_is_forwarding_26 = l_forwarders_26_0 | l_forwarders_26_1;
  wire [4:0]  l_forward_stq_idx_26 = l_is_forwarding_26 ? (l_forwarders_26_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_26_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_26_bits_forward_stq_idx;
  wire        block_addr_matches_26_1 = lcam_addr_1[39:6] == ldq_26_bits_addr_bits[39:6];
  wire        dword_addr_matches_26_0 = lcam_addr_0[39:6] == ldq_26_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_26_bits_addr_bits[5:3];
  wire        dword_addr_matches_26_1 = block_addr_matches_26_1 & lcam_addr_1[5:3] == ldq_26_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_104 = casez_tmp_138 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_106 = casez_tmp_138 & casez_tmp_109;
  wire        _GEN_867 = ldq_26_bits_executed | ldq_26_bits_succeeded;
  wire        _GEN_868 = _GEN_867 | l_is_forwarding_26;
  wire [31:0] _GEN_869 = ldq_26_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_870 = do_st_search_0 & ldq_26_valid & ldq_26_bits_addr_valid & _GEN_868 & ~ldq_26_bits_addr_is_virtual & _GEN_869[0] & dword_addr_matches_26_0 & (|_mask_overlap_T_104);
  wire        _forwarded_is_older_T_213 = l_forward_stq_idx_26 < ldq_26_bits_youngest_stq_idx;
  wire        _GEN_96044 = ~ldq_26_bits_forward_std_val | l_forward_stq_idx_26 != lcam_stq_idx_0 & (l_forward_stq_idx_26 < lcam_stq_idx_0 ^ _forwarded_is_older_T_213 ^ lcam_stq_idx_0 < ldq_26_bits_youngest_stq_idx);
  wire        _GEN_871 = _do_ld_search_T_2 & ldq_26_valid & ldq_26_bits_addr_valid & ~ldq_26_bits_addr_is_virtual & dword_addr_matches_26_0 & (|_mask_overlap_T_104);
  wire        _searcher_is_older_T_215 = ldq_head > 5'h1A;
  wire        searcher_is_older_52 = lcam_ldq_idx_0 < 5'h1A ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_215;
  wire        _GEN_872 = _GEN_868 & ~s1_executing_loads_26;
  wire        _GEN_96046 = _GEN_872 & ldq_26_bits_observed;
  wire        _GEN_873 = lcam_ldq_idx_0 != 5'h1A;
  reg         older_nacked_REG_52;
  wire        _GEN_116721 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1A;
  wire        _GEN_874 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1A;
  wire        nacking_loads_26 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_874 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116721;
  wire        _GEN_875 = ~_GEN_867 | nacking_loads_26 | older_nacked_REG_52;
  reg         io_dmem_s1_kill_0_REG_26;
  wire        _GEN_96220 = _GEN_870 ? _GEN_96044 : _GEN_871 & searcher_is_older_52 & _GEN_96046;
  wire        _GEN_876 = _GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875);
  wire        _GEN_877 = fired_release_1 & ldq_26_valid & ldq_26_bits_addr_valid & block_addr_matches_26_1;
  wire [31:0] _GEN_878 = ldq_26_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_879 = do_st_search_1 & ldq_26_valid & ldq_26_bits_addr_valid & _GEN_868 & ~ldq_26_bits_addr_is_virtual & _GEN_878[0] & dword_addr_matches_26_1 & (|_mask_overlap_T_106);
  wire        _GEN_880 = ~ldq_26_bits_forward_std_val | l_forward_stq_idx_26 != lcam_stq_idx_1 & (l_forward_stq_idx_26 < lcam_stq_idx_1 ^ _forwarded_is_older_T_213 ^ lcam_stq_idx_1 < ldq_26_bits_youngest_stq_idx);
  wire        _GEN_881 = do_ld_search_1 & ldq_26_valid & ldq_26_bits_addr_valid & ~ldq_26_bits_addr_is_virtual & dword_addr_matches_26_1 & (|_mask_overlap_T_106);
  wire        searcher_is_older_53 = lcam_ldq_idx_1 < 5'h1A ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_215;
  wire        _GEN_882 = lcam_ldq_idx_1 != 5'h1A;
  reg         older_nacked_REG_53;
  wire        _GEN_883 = ~_GEN_867 | nacking_loads_26 | older_nacked_REG_53;
  reg         io_dmem_s1_kill_1_REG_26;
  wire        _GEN_884 = _GEN_881 & searcher_is_older_53 & _GEN_872 & ldq_26_bits_observed;
  wire        failed_loads_26 = _GEN_877 ? _GEN_96220 : _GEN_879 ? _GEN_880 | _GEN_96220 : _GEN_884 | _GEN_96220;
  wire        _GEN_885 = _GEN_877 | _GEN_879;
  wire        _GEN_886 = _GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883);
  wire [14:0] _l_mask_mask_T_407 = 15'h1 << ldq_27_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_411 = 15'h3 << {12'h0, ldq_27_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_27_bits_uop_mem_size)
      2'b00:
        casez_tmp_139 = _l_mask_mask_T_407[7:0];
      2'b01:
        casez_tmp_139 = _l_mask_mask_T_411[7:0];
      2'b10:
        casez_tmp_139 = ldq_27_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_139 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_27_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1B;
  wire        l_forwarders_27_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1B;
  wire        l_is_forwarding_27 = l_forwarders_27_0 | l_forwarders_27_1;
  wire [4:0]  l_forward_stq_idx_27 = l_is_forwarding_27 ? (l_forwarders_27_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_27_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_27_bits_forward_stq_idx;
  wire        block_addr_matches_27_1 = lcam_addr_1[39:6] == ldq_27_bits_addr_bits[39:6];
  wire        dword_addr_matches_27_0 = lcam_addr_0[39:6] == ldq_27_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_27_bits_addr_bits[5:3];
  wire        dword_addr_matches_27_1 = block_addr_matches_27_1 & lcam_addr_1[5:3] == ldq_27_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_108 = casez_tmp_139 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_110 = casez_tmp_139 & casez_tmp_109;
  wire        _GEN_887 = ldq_27_bits_executed | ldq_27_bits_succeeded;
  wire        _GEN_888 = _GEN_887 | l_is_forwarding_27;
  wire [31:0] _GEN_889 = ldq_27_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_890 = do_st_search_0 & ldq_27_valid & ldq_27_bits_addr_valid & _GEN_888 & ~ldq_27_bits_addr_is_virtual & _GEN_889[0] & dword_addr_matches_27_0 & (|_mask_overlap_T_108);
  wire        _forwarded_is_older_T_221 = l_forward_stq_idx_27 < ldq_27_bits_youngest_stq_idx;
  wire        _GEN_96542 = ~ldq_27_bits_forward_std_val | l_forward_stq_idx_27 != lcam_stq_idx_0 & (l_forward_stq_idx_27 < lcam_stq_idx_0 ^ _forwarded_is_older_T_221 ^ lcam_stq_idx_0 < ldq_27_bits_youngest_stq_idx);
  wire        _GEN_891 = _do_ld_search_T_2 & ldq_27_valid & ldq_27_bits_addr_valid & ~ldq_27_bits_addr_is_virtual & dword_addr_matches_27_0 & (|_mask_overlap_T_108);
  wire        _searcher_is_older_T_223 = ldq_head > 5'h1B;
  wire        searcher_is_older_54 = lcam_ldq_idx_0 < 5'h1B ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_223;
  wire        _GEN_892 = _GEN_888 & ~s1_executing_loads_27;
  wire        _GEN_96544 = _GEN_892 & ldq_27_bits_observed;
  wire        _GEN_893 = lcam_ldq_idx_0 != 5'h1B;
  reg         older_nacked_REG_54;
  wire        _GEN_116722 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1B;
  wire        _GEN_894 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1B;
  wire        nacking_loads_27 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_894 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116722;
  wire        _GEN_895 = ~_GEN_887 | nacking_loads_27 | older_nacked_REG_54;
  reg         io_dmem_s1_kill_0_REG_27;
  wire        _GEN_96718 = _GEN_890 ? _GEN_96542 : _GEN_891 & searcher_is_older_54 & _GEN_96544;
  wire        _GEN_896 = _GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895);
  wire        _GEN_897 = fired_release_1 & ldq_27_valid & ldq_27_bits_addr_valid & block_addr_matches_27_1;
  wire [31:0] _GEN_898 = ldq_27_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_899 = do_st_search_1 & ldq_27_valid & ldq_27_bits_addr_valid & _GEN_888 & ~ldq_27_bits_addr_is_virtual & _GEN_898[0] & dword_addr_matches_27_1 & (|_mask_overlap_T_110);
  wire        _GEN_900 = ~ldq_27_bits_forward_std_val | l_forward_stq_idx_27 != lcam_stq_idx_1 & (l_forward_stq_idx_27 < lcam_stq_idx_1 ^ _forwarded_is_older_T_221 ^ lcam_stq_idx_1 < ldq_27_bits_youngest_stq_idx);
  wire        _GEN_901 = do_ld_search_1 & ldq_27_valid & ldq_27_bits_addr_valid & ~ldq_27_bits_addr_is_virtual & dword_addr_matches_27_1 & (|_mask_overlap_T_110);
  wire        searcher_is_older_55 = lcam_ldq_idx_1 < 5'h1B ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_223;
  wire        _GEN_902 = lcam_ldq_idx_1 != 5'h1B;
  reg         older_nacked_REG_55;
  wire        _GEN_903 = ~_GEN_887 | nacking_loads_27 | older_nacked_REG_55;
  reg         io_dmem_s1_kill_1_REG_27;
  wire        _GEN_904 = _GEN_901 & searcher_is_older_55 & _GEN_892 & ldq_27_bits_observed;
  wire        failed_loads_27 = _GEN_897 ? _GEN_96718 : _GEN_899 ? _GEN_900 | _GEN_96718 : _GEN_904 | _GEN_96718;
  wire        _GEN_905 = _GEN_897 | _GEN_899;
  wire        _GEN_906 = _GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903);
  wire [14:0] _l_mask_mask_T_422 = 15'h1 << ldq_28_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_426 = 15'h3 << {12'h0, ldq_28_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_28_bits_uop_mem_size)
      2'b00:
        casez_tmp_140 = _l_mask_mask_T_422[7:0];
      2'b01:
        casez_tmp_140 = _l_mask_mask_T_426[7:0];
      2'b10:
        casez_tmp_140 = ldq_28_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_140 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_28_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1C;
  wire        l_forwarders_28_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1C;
  wire        l_is_forwarding_28 = l_forwarders_28_0 | l_forwarders_28_1;
  wire [4:0]  l_forward_stq_idx_28 = l_is_forwarding_28 ? (l_forwarders_28_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_28_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_28_bits_forward_stq_idx;
  wire        block_addr_matches_28_1 = lcam_addr_1[39:6] == ldq_28_bits_addr_bits[39:6];
  wire        dword_addr_matches_28_0 = lcam_addr_0[39:6] == ldq_28_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_28_bits_addr_bits[5:3];
  wire        dword_addr_matches_28_1 = block_addr_matches_28_1 & lcam_addr_1[5:3] == ldq_28_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_112 = casez_tmp_140 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_114 = casez_tmp_140 & casez_tmp_109;
  wire        _GEN_907 = ldq_28_bits_executed | ldq_28_bits_succeeded;
  wire        _GEN_908 = _GEN_907 | l_is_forwarding_28;
  wire [31:0] _GEN_909 = ldq_28_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_910 = do_st_search_0 & ldq_28_valid & ldq_28_bits_addr_valid & _GEN_908 & ~ldq_28_bits_addr_is_virtual & _GEN_909[0] & dword_addr_matches_28_0 & (|_mask_overlap_T_112);
  wire        _forwarded_is_older_T_229 = l_forward_stq_idx_28 < ldq_28_bits_youngest_stq_idx;
  wire        _GEN_97040 = ~ldq_28_bits_forward_std_val | l_forward_stq_idx_28 != lcam_stq_idx_0 & (l_forward_stq_idx_28 < lcam_stq_idx_0 ^ _forwarded_is_older_T_229 ^ lcam_stq_idx_0 < ldq_28_bits_youngest_stq_idx);
  wire        _GEN_911 = _do_ld_search_T_2 & ldq_28_valid & ldq_28_bits_addr_valid & ~ldq_28_bits_addr_is_virtual & dword_addr_matches_28_0 & (|_mask_overlap_T_112);
  wire        _searcher_is_older_T_231 = ldq_head > 5'h1C;
  wire        searcher_is_older_56 = lcam_ldq_idx_0[4:2] != 3'h7 ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_231;
  wire        _GEN_912 = _GEN_908 & ~s1_executing_loads_28;
  wire        _GEN_97042 = _GEN_912 & ldq_28_bits_observed;
  wire        _GEN_913 = lcam_ldq_idx_0 != 5'h1C;
  reg         older_nacked_REG_56;
  wire        _GEN_116723 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1C;
  wire        _GEN_914 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1C;
  wire        nacking_loads_28 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_914 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116723;
  wire        _GEN_915 = ~_GEN_907 | nacking_loads_28 | older_nacked_REG_56;
  reg         io_dmem_s1_kill_0_REG_28;
  wire        _GEN_97216 = _GEN_910 ? _GEN_97040 : _GEN_911 & searcher_is_older_56 & _GEN_97042;
  wire        _GEN_916 = _GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915);
  wire        _GEN_917 = fired_release_1 & ldq_28_valid & ldq_28_bits_addr_valid & block_addr_matches_28_1;
  wire [31:0] _GEN_918 = ldq_28_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_919 = do_st_search_1 & ldq_28_valid & ldq_28_bits_addr_valid & _GEN_908 & ~ldq_28_bits_addr_is_virtual & _GEN_918[0] & dword_addr_matches_28_1 & (|_mask_overlap_T_114);
  wire        _GEN_920 = ~ldq_28_bits_forward_std_val | l_forward_stq_idx_28 != lcam_stq_idx_1 & (l_forward_stq_idx_28 < lcam_stq_idx_1 ^ _forwarded_is_older_T_229 ^ lcam_stq_idx_1 < ldq_28_bits_youngest_stq_idx);
  wire        _GEN_921 = do_ld_search_1 & ldq_28_valid & ldq_28_bits_addr_valid & ~ldq_28_bits_addr_is_virtual & dword_addr_matches_28_1 & (|_mask_overlap_T_114);
  wire        searcher_is_older_57 = lcam_ldq_idx_1[4:2] != 3'h7 ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_231;
  wire        _GEN_922 = lcam_ldq_idx_1 != 5'h1C;
  reg         older_nacked_REG_57;
  wire        _GEN_923 = ~_GEN_907 | nacking_loads_28 | older_nacked_REG_57;
  reg         io_dmem_s1_kill_1_REG_28;
  wire        _GEN_924 = _GEN_921 & searcher_is_older_57 & _GEN_912 & ldq_28_bits_observed;
  wire        failed_loads_28 = _GEN_917 ? _GEN_97216 : _GEN_919 ? _GEN_920 | _GEN_97216 : _GEN_924 | _GEN_97216;
  wire        _GEN_925 = _GEN_917 | _GEN_919;
  wire        _GEN_926 = _GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923);
  wire [14:0] _l_mask_mask_T_437 = 15'h1 << ldq_29_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_441 = 15'h3 << {12'h0, ldq_29_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_29_bits_uop_mem_size)
      2'b00:
        casez_tmp_141 = _l_mask_mask_T_437[7:0];
      2'b01:
        casez_tmp_141 = _l_mask_mask_T_441[7:0];
      2'b10:
        casez_tmp_141 = ldq_29_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_141 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_29_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1D;
  wire        l_forwarders_29_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1D;
  wire        l_is_forwarding_29 = l_forwarders_29_0 | l_forwarders_29_1;
  wire [4:0]  l_forward_stq_idx_29 = l_is_forwarding_29 ? (l_forwarders_29_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_29_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_29_bits_forward_stq_idx;
  wire        block_addr_matches_29_1 = lcam_addr_1[39:6] == ldq_29_bits_addr_bits[39:6];
  wire        dword_addr_matches_29_0 = lcam_addr_0[39:6] == ldq_29_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_29_bits_addr_bits[5:3];
  wire        dword_addr_matches_29_1 = block_addr_matches_29_1 & lcam_addr_1[5:3] == ldq_29_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_116 = casez_tmp_141 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_118 = casez_tmp_141 & casez_tmp_109;
  wire        _GEN_927 = ldq_29_bits_executed | ldq_29_bits_succeeded;
  wire        _GEN_928 = _GEN_927 | l_is_forwarding_29;
  wire [31:0] _GEN_929 = ldq_29_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_930 = do_st_search_0 & ldq_29_valid & ldq_29_bits_addr_valid & _GEN_928 & ~ldq_29_bits_addr_is_virtual & _GEN_929[0] & dword_addr_matches_29_0 & (|_mask_overlap_T_116);
  wire        _forwarded_is_older_T_237 = l_forward_stq_idx_29 < ldq_29_bits_youngest_stq_idx;
  wire        _GEN_97538 = ~ldq_29_bits_forward_std_val | l_forward_stq_idx_29 != lcam_stq_idx_0 & (l_forward_stq_idx_29 < lcam_stq_idx_0 ^ _forwarded_is_older_T_237 ^ lcam_stq_idx_0 < ldq_29_bits_youngest_stq_idx);
  wire        _GEN_931 = _do_ld_search_T_2 & ldq_29_valid & ldq_29_bits_addr_valid & ~ldq_29_bits_addr_is_virtual & dword_addr_matches_29_0 & (|_mask_overlap_T_116);
  wire        _searcher_is_older_T_239 = ldq_head > 5'h1D;
  wire        searcher_is_older_58 = lcam_ldq_idx_0 < 5'h1D ^ _searcher_is_older_T_249 ^ _searcher_is_older_T_239;
  wire        _GEN_932 = _GEN_928 & ~s1_executing_loads_29;
  wire        _GEN_97540 = _GEN_932 & ldq_29_bits_observed;
  wire        _GEN_933 = lcam_ldq_idx_0 != 5'h1D;
  reg         older_nacked_REG_58;
  wire        _GEN_116724 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1D;
  wire        _GEN_934 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1D;
  wire        nacking_loads_29 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_934 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116724;
  wire        _GEN_935 = ~_GEN_927 | nacking_loads_29 | older_nacked_REG_58;
  reg         io_dmem_s1_kill_0_REG_29;
  wire        _GEN_97714 = _GEN_930 ? _GEN_97538 : _GEN_931 & searcher_is_older_58 & _GEN_97540;
  wire        _GEN_936 = _GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935);
  wire        _GEN_937 = fired_release_1 & ldq_29_valid & ldq_29_bits_addr_valid & block_addr_matches_29_1;
  wire [31:0] _GEN_938 = ldq_29_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_939 = do_st_search_1 & ldq_29_valid & ldq_29_bits_addr_valid & _GEN_928 & ~ldq_29_bits_addr_is_virtual & _GEN_938[0] & dword_addr_matches_29_1 & (|_mask_overlap_T_118);
  wire        _GEN_940 = ~ldq_29_bits_forward_std_val | l_forward_stq_idx_29 != lcam_stq_idx_1 & (l_forward_stq_idx_29 < lcam_stq_idx_1 ^ _forwarded_is_older_T_237 ^ lcam_stq_idx_1 < ldq_29_bits_youngest_stq_idx);
  wire        _GEN_941 = do_ld_search_1 & ldq_29_valid & ldq_29_bits_addr_valid & ~ldq_29_bits_addr_is_virtual & dword_addr_matches_29_1 & (|_mask_overlap_T_118);
  wire        searcher_is_older_59 = lcam_ldq_idx_1 < 5'h1D ^ _searcher_is_older_T_253 ^ _searcher_is_older_T_239;
  wire        _GEN_942 = lcam_ldq_idx_1 != 5'h1D;
  reg         older_nacked_REG_59;
  wire        _GEN_943 = ~_GEN_927 | nacking_loads_29 | older_nacked_REG_59;
  reg         io_dmem_s1_kill_1_REG_29;
  wire        _GEN_944 = _GEN_941 & searcher_is_older_59 & _GEN_932 & ldq_29_bits_observed;
  wire        failed_loads_29 = _GEN_937 ? _GEN_97714 : _GEN_939 ? _GEN_940 | _GEN_97714 : _GEN_944 | _GEN_97714;
  wire        _GEN_945 = _GEN_937 | _GEN_939;
  wire        _GEN_946 = _GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943);
  wire [14:0] _l_mask_mask_T_452 = 15'h1 << ldq_30_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_456 = 15'h3 << {12'h0, ldq_30_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_30_bits_uop_mem_size)
      2'b00:
        casez_tmp_142 = _l_mask_mask_T_452[7:0];
      2'b01:
        casez_tmp_142 = _l_mask_mask_T_456[7:0];
      2'b10:
        casez_tmp_142 = ldq_30_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_142 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_30_0 = wb_forward_valid_0 & wb_forward_ldq_idx_0 == 5'h1E;
  wire        l_forwarders_30_1 = wb_forward_valid_1 & wb_forward_ldq_idx_1 == 5'h1E;
  wire        l_is_forwarding_30 = l_forwarders_30_0 | l_forwarders_30_1;
  wire [4:0]  l_forward_stq_idx_30 = l_is_forwarding_30 ? (l_forwarders_30_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_30_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_30_bits_forward_stq_idx;
  wire        block_addr_matches_30_1 = lcam_addr_1[39:6] == ldq_30_bits_addr_bits[39:6];
  wire        dword_addr_matches_30_0 = lcam_addr_0[39:6] == ldq_30_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_30_bits_addr_bits[5:3];
  wire        dword_addr_matches_30_1 = block_addr_matches_30_1 & lcam_addr_1[5:3] == ldq_30_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_120 = casez_tmp_142 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_122 = casez_tmp_142 & casez_tmp_109;
  wire        _GEN_947 = ldq_30_bits_executed | ldq_30_bits_succeeded;
  wire        _GEN_948 = _GEN_947 | l_is_forwarding_30;
  wire [31:0] _GEN_949 = ldq_30_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_950 = do_st_search_0 & ldq_30_valid & ldq_30_bits_addr_valid & _GEN_948 & ~ldq_30_bits_addr_is_virtual & _GEN_949[0] & dword_addr_matches_30_0 & (|_mask_overlap_T_120);
  wire        _forwarded_is_older_T_245 = l_forward_stq_idx_30 < ldq_30_bits_youngest_stq_idx;
  wire        _GEN_98036 = ~ldq_30_bits_forward_std_val | l_forward_stq_idx_30 != lcam_stq_idx_0 & (l_forward_stq_idx_30 < lcam_stq_idx_0 ^ _forwarded_is_older_T_245 ^ lcam_stq_idx_0 < ldq_30_bits_youngest_stq_idx);
  wire        _GEN_951 = _do_ld_search_T_2 & ldq_30_valid & ldq_30_bits_addr_valid & ~ldq_30_bits_addr_is_virtual & dword_addr_matches_30_0 & (|_mask_overlap_T_120);
  wire        searcher_is_older_60 = lcam_ldq_idx_0[4:1] != 4'hF ^ _searcher_is_older_T_249 ^ (&ldq_head);
  wire        _GEN_952 = _GEN_948 & ~s1_executing_loads_30;
  wire        _GEN_98038 = _GEN_952 & ldq_30_bits_observed;
  wire        _GEN_953 = lcam_ldq_idx_0 != 5'h1E;
  reg         older_nacked_REG_60;
  wire        _GEN_116725 = io_dmem_nack_0_bits_uop_ldq_idx == 5'h1E;
  wire        _GEN_954 = io_dmem_nack_1_bits_uop_uses_ldq & io_dmem_nack_1_bits_uop_ldq_idx == 5'h1E;
  wire        nacking_loads_30 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_954 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116725;
  wire        _GEN_955 = ~_GEN_947 | nacking_loads_30 | older_nacked_REG_60;
  reg         io_dmem_s1_kill_0_REG_30;
  wire        _GEN_98212 = _GEN_950 ? _GEN_98036 : _GEN_951 & searcher_is_older_60 & _GEN_98038;
  wire        _GEN_956 = _GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955);
  wire        _GEN_957 = fired_release_1 & ldq_30_valid & ldq_30_bits_addr_valid & block_addr_matches_30_1;
  wire [31:0] _GEN_958 = ldq_30_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_959 = do_st_search_1 & ldq_30_valid & ldq_30_bits_addr_valid & _GEN_948 & ~ldq_30_bits_addr_is_virtual & _GEN_958[0] & dword_addr_matches_30_1 & (|_mask_overlap_T_122);
  wire        _GEN_960 = ~ldq_30_bits_forward_std_val | l_forward_stq_idx_30 != lcam_stq_idx_1 & (l_forward_stq_idx_30 < lcam_stq_idx_1 ^ _forwarded_is_older_T_245 ^ lcam_stq_idx_1 < ldq_30_bits_youngest_stq_idx);
  wire        _GEN_961 = do_ld_search_1 & ldq_30_valid & ldq_30_bits_addr_valid & ~ldq_30_bits_addr_is_virtual & dword_addr_matches_30_1 & (|_mask_overlap_T_122);
  wire        searcher_is_older_61 = lcam_ldq_idx_1[4:1] != 4'hF ^ _searcher_is_older_T_253 ^ (&ldq_head);
  wire        _GEN_962 = lcam_ldq_idx_1 != 5'h1E;
  reg         older_nacked_REG_61;
  wire        _GEN_963 = ~_GEN_947 | nacking_loads_30 | older_nacked_REG_61;
  reg         io_dmem_s1_kill_1_REG_30;
  wire        _GEN_964 = _GEN_961 & searcher_is_older_61 & _GEN_952 & ldq_30_bits_observed;
  wire        failed_loads_30 = _GEN_957 ? _GEN_98212 : _GEN_959 ? _GEN_960 | _GEN_98212 : _GEN_964 | _GEN_98212;
  wire        _GEN_965 = _GEN_957 | _GEN_959;
  wire        _GEN_966 = _GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963);
  wire [14:0] _l_mask_mask_T_467 = 15'h1 << ldq_31_bits_addr_bits[2:0];
  wire [14:0] _l_mask_mask_T_471 = 15'h3 << {12'h0, ldq_31_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (ldq_31_bits_uop_mem_size)
      2'b00:
        casez_tmp_143 = _l_mask_mask_T_467[7:0];
      2'b01:
        casez_tmp_143 = _l_mask_mask_T_471[7:0];
      2'b10:
        casez_tmp_143 = ldq_31_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_143 = 8'hFF;
    endcase
  end // always @(*)
  wire        l_forwarders_31_0 = wb_forward_valid_0 & (&wb_forward_ldq_idx_0);
  wire        l_forwarders_31_1 = wb_forward_valid_1 & (&wb_forward_ldq_idx_1);
  wire        l_is_forwarding_31 = l_forwarders_31_0 | l_forwarders_31_1;
  wire [4:0]  l_forward_stq_idx_31 = l_is_forwarding_31 ? (l_forwarders_31_0 ? wb_forward_stq_idx_0 : 5'h0) | (l_forwarders_31_1 ? wb_forward_stq_idx_1 : 5'h0) : ldq_31_bits_forward_stq_idx;
  wire        block_addr_matches_31_1 = lcam_addr_1[39:6] == ldq_31_bits_addr_bits[39:6];
  wire        dword_addr_matches_31_0 = lcam_addr_0[39:6] == ldq_31_bits_addr_bits[39:6] & lcam_addr_0[5:3] == ldq_31_bits_addr_bits[5:3];
  wire        dword_addr_matches_31_1 = block_addr_matches_31_1 & lcam_addr_1[5:3] == ldq_31_bits_addr_bits[5:3];
  wire [7:0]  _mask_overlap_T_124 = casez_tmp_143 & casez_tmp_108;
  wire [7:0]  _mask_overlap_T_126 = casez_tmp_143 & casez_tmp_109;
  wire        _GEN_967 = ldq_31_bits_executed | ldq_31_bits_succeeded;
  wire        _GEN_968 = _GEN_967 | l_is_forwarding_31;
  wire [31:0] _GEN_969 = ldq_31_bits_st_dep_mask >> _GEN_349;
  wire        _GEN_970 = do_st_search_0 & ldq_31_valid & ldq_31_bits_addr_valid & _GEN_968 & ~ldq_31_bits_addr_is_virtual & _GEN_969[0] & dword_addr_matches_31_0 & (|_mask_overlap_T_124);
  wire        _forwarded_is_older_T_253 = l_forward_stq_idx_31 < ldq_31_bits_youngest_stq_idx;
  wire        _GEN_98534 = ~ldq_31_bits_forward_std_val | l_forward_stq_idx_31 != lcam_stq_idx_0 & (l_forward_stq_idx_31 < lcam_stq_idx_0 ^ _forwarded_is_older_T_253 ^ lcam_stq_idx_0 < ldq_31_bits_youngest_stq_idx);
  wire        _GEN_971 = _do_ld_search_T_2 & ldq_31_valid & ldq_31_bits_addr_valid & ~ldq_31_bits_addr_is_virtual & dword_addr_matches_31_0 & (|_mask_overlap_T_124);
  wire        searcher_is_older_62 = lcam_ldq_idx_0 != 5'h1F ^ _searcher_is_older_T_249;
  wire        _GEN_972 = _GEN_968 & ~s1_executing_loads_31;
  wire        _GEN_98536 = _GEN_972 & ldq_31_bits_observed;
  reg         older_nacked_REG_62;
  wire        _GEN_973 = io_dmem_nack_1_bits_uop_uses_ldq & (&io_dmem_nack_1_bits_uop_ldq_idx);
  wire        nacking_loads_31 = io_dmem_nack_1_valid & ~io_dmem_nack_1_bits_is_hella & _GEN_973 | io_dmem_nack_0_valid & ~io_dmem_nack_0_bits_is_hella & io_dmem_nack_0_bits_uop_uses_ldq & (&io_dmem_nack_0_bits_uop_ldq_idx);
  wire        _GEN_974 = ~_GEN_967 | nacking_loads_31 | older_nacked_REG_62;
  reg         io_dmem_s1_kill_0_REG_31;
  wire        _GEN_98710 = _GEN_970 ? _GEN_98534 : _GEN_971 & searcher_is_older_62 & _GEN_98536;
  wire        _GEN_975 = _GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974);
  wire        _GEN_98780 = _GEN_975 ? (_GEN_956 ? (_GEN_936 ? (_GEN_916 ? (_GEN_896 ? (_GEN_876 ? (_GEN_856 ? (_GEN_836 ? (_GEN_816 ? (_GEN_796 ? (_GEN_776 ? (_GEN_756 ? (_GEN_736 ? (_GEN_716 ? (_GEN_696 ? (_GEN_676 ? (_GEN_656 ? (_GEN_636 ? (_GEN_616 ? (_GEN_596 ? (_GEN_576 ? (_GEN_556 ? (_GEN_536 ? (_GEN_516 ? (_GEN_496 ? (_GEN_476 ? (_GEN_456 ? (_GEN_436 ? (_GEN_416 ? (_GEN_396 ? (_GEN_376 ? ~_GEN_351 & _GEN_352 & ~searcher_is_older & _GEN_356 & io_dmem_s1_kill_0_REG : io_dmem_s1_kill_0_REG_1) : io_dmem_s1_kill_0_REG_2) : io_dmem_s1_kill_0_REG_3) : io_dmem_s1_kill_0_REG_4) : io_dmem_s1_kill_0_REG_5) : io_dmem_s1_kill_0_REG_6) : io_dmem_s1_kill_0_REG_7) : io_dmem_s1_kill_0_REG_8) : io_dmem_s1_kill_0_REG_9) : io_dmem_s1_kill_0_REG_10) : io_dmem_s1_kill_0_REG_11) : io_dmem_s1_kill_0_REG_12) : io_dmem_s1_kill_0_REG_13) : io_dmem_s1_kill_0_REG_14) : io_dmem_s1_kill_0_REG_15) : io_dmem_s1_kill_0_REG_16) : io_dmem_s1_kill_0_REG_17) : io_dmem_s1_kill_0_REG_18) : io_dmem_s1_kill_0_REG_19) : io_dmem_s1_kill_0_REG_20) : io_dmem_s1_kill_0_REG_21) : io_dmem_s1_kill_0_REG_22) : io_dmem_s1_kill_0_REG_23) : io_dmem_s1_kill_0_REG_24) : io_dmem_s1_kill_0_REG_25) : io_dmem_s1_kill_0_REG_26) : io_dmem_s1_kill_0_REG_27) : io_dmem_s1_kill_0_REG_28) : io_dmem_s1_kill_0_REG_29) : io_dmem_s1_kill_0_REG_30) : io_dmem_s1_kill_0_REG_31;
  wire        can_forward_0 = _GEN_975 & _GEN_956 & _GEN_936 & _GEN_916 & _GEN_896 & _GEN_876 & _GEN_856 & _GEN_836 & _GEN_816 & _GEN_796 & _GEN_776 & _GEN_756 & _GEN_736 & _GEN_716 & _GEN_696 & _GEN_676 & _GEN_656 & _GEN_636 & _GEN_616 & _GEN_596 & _GEN_576 & _GEN_556 & _GEN_536 & _GEN_516 & _GEN_496 & _GEN_476 & _GEN_456 & _GEN_436 & _GEN_416 & _GEN_396 & _GEN_376 & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~_GEN_356) & (fired_load_incoming_0 ? ~mem_tlb_uncacheable_0 : ~casez_tmp_110);
  wire        _GEN_976 = fired_release_1 & ldq_31_valid & ldq_31_bits_addr_valid & block_addr_matches_31_1;
  wire [31:0] _GEN_977 = ldq_31_bits_st_dep_mask >> _GEN_358;
  wire        _GEN_978 = do_st_search_1 & ldq_31_valid & ldq_31_bits_addr_valid & _GEN_968 & ~ldq_31_bits_addr_is_virtual & _GEN_977[0] & dword_addr_matches_31_1 & (|_mask_overlap_T_126);
  wire        _GEN_979 = ~ldq_31_bits_forward_std_val | l_forward_stq_idx_31 != lcam_stq_idx_1 & (l_forward_stq_idx_31 < lcam_stq_idx_1 ^ _forwarded_is_older_T_253 ^ lcam_stq_idx_1 < ldq_31_bits_youngest_stq_idx);
  wire        _GEN_980 = do_ld_search_1 & ldq_31_valid & ldq_31_bits_addr_valid & ~ldq_31_bits_addr_is_virtual & dword_addr_matches_31_1 & (|_mask_overlap_T_126);
  wire        searcher_is_older_63 = lcam_ldq_idx_1 != 5'h1F ^ _searcher_is_older_T_253;
  reg         older_nacked_REG_63;
  wire        _GEN_981 = ~_GEN_967 | nacking_loads_31 | older_nacked_REG_63;
  reg         io_dmem_s1_kill_1_REG_31;
  wire        _GEN_982 = _GEN_980 & searcher_is_older_63 & _GEN_972 & ldq_31_bits_observed;
  wire        failed_loads_31 = _GEN_976 ? _GEN_98710 : _GEN_978 ? _GEN_979 | _GEN_98710 : _GEN_982 | _GEN_98710;
  wire        _GEN_983 = _GEN_976 | _GEN_978;
  wire        _GEN_984 = _GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981);
  wire        _GEN_99029 = _GEN_984 ? (_GEN_966 ? (_GEN_946 ? (_GEN_926 ? (_GEN_906 ? (_GEN_886 ? (_GEN_866 ? (_GEN_846 ? (_GEN_826 ? (_GEN_806 ? (_GEN_786 ? (_GEN_766 ? (_GEN_746 ? (_GEN_726 ? (_GEN_706 ? (_GEN_686 ? (_GEN_666 ? (_GEN_646 ? (_GEN_626 ? (_GEN_606 ? (_GEN_586 ? (_GEN_566 ? (_GEN_546 ? (_GEN_526 ? (_GEN_506 ? (_GEN_486 ? (_GEN_466 ? (_GEN_446 ? (_GEN_426 ? (_GEN_406 ? (_GEN_386 ? ~_GEN_366 & _GEN_362 & ~searcher_is_older_1 & _GEN_364 & io_dmem_s1_kill_1_REG : io_dmem_s1_kill_1_REG_1) : io_dmem_s1_kill_1_REG_2) : io_dmem_s1_kill_1_REG_3) : io_dmem_s1_kill_1_REG_4) : io_dmem_s1_kill_1_REG_5) : io_dmem_s1_kill_1_REG_6) : io_dmem_s1_kill_1_REG_7) : io_dmem_s1_kill_1_REG_8) : io_dmem_s1_kill_1_REG_9) : io_dmem_s1_kill_1_REG_10) : io_dmem_s1_kill_1_REG_11) : io_dmem_s1_kill_1_REG_12) : io_dmem_s1_kill_1_REG_13) : io_dmem_s1_kill_1_REG_14) : io_dmem_s1_kill_1_REG_15) : io_dmem_s1_kill_1_REG_16) : io_dmem_s1_kill_1_REG_17) : io_dmem_s1_kill_1_REG_18) : io_dmem_s1_kill_1_REG_19) : io_dmem_s1_kill_1_REG_20) : io_dmem_s1_kill_1_REG_21) : io_dmem_s1_kill_1_REG_22) : io_dmem_s1_kill_1_REG_23) : io_dmem_s1_kill_1_REG_24) : io_dmem_s1_kill_1_REG_25) : io_dmem_s1_kill_1_REG_26) : io_dmem_s1_kill_1_REG_27) : io_dmem_s1_kill_1_REG_28) : io_dmem_s1_kill_1_REG_29) : io_dmem_s1_kill_1_REG_30) : io_dmem_s1_kill_1_REG_31;
  wire        can_forward_1 = _GEN_984 & _GEN_966 & _GEN_946 & _GEN_926 & _GEN_906 & _GEN_886 & _GEN_866 & _GEN_846 & _GEN_826 & _GEN_806 & _GEN_786 & _GEN_766 & _GEN_746 & _GEN_726 & _GEN_706 & _GEN_686 & _GEN_666 & _GEN_646 & _GEN_626 & _GEN_606 & _GEN_586 & _GEN_566 & _GEN_546 & _GEN_526 & _GEN_506 & _GEN_486 & _GEN_466 & _GEN_446 & _GEN_426 & _GEN_406 & _GEN_386 & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~_GEN_364) & (_can_forward_T_6 ? ~mem_tlb_uncacheable_1 : ~casez_tmp_111);
  wire        dword_addr_matches_32_0 = stq_0_bits_addr_valid & ~stq_0_bits_addr_is_virtual & stq_0_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_32_1 = stq_0_bits_addr_valid & ~stq_0_bits_addr_is_virtual & stq_0_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_2 = 15'h1 << stq_0_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_6 = 15'h3 << {12'h0, stq_0_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_0_bits_uop_mem_size)
      2'b00:
        casez_tmp_144 = _write_mask_mask_T_2[7:0];
      2'b01:
        casez_tmp_144 = _write_mask_mask_T_6[7:0];
      2'b10:
        casez_tmp_144 = stq_0_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_144 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_985 = _do_ld_search_T_2 & stq_0_valid & lcam_st_dep_mask_0[0];
  wire [7:0]  _GEN_986 = casez_tmp_108 & casez_tmp_144;
  wire        _GEN_99196 = _GEN_986 == casez_tmp_108 & ~stq_0_bits_uop_is_fence & ~stq_0_bits_uop_is_amo & dword_addr_matches_32_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_32;
  wire        _GEN_987 = (|_GEN_986) & dword_addr_matches_32_0;
  reg         io_dmem_s1_kill_0_REG_33;
  wire        _GEN_99361 = stq_0_bits_uop_is_fence | stq_0_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_34;
  wire        _GEN_99232 = _GEN_985 ? (_GEN_99196 ? io_dmem_s1_kill_0_REG_32 : _GEN_987 ? io_dmem_s1_kill_0_REG_33 : _GEN_99361 ? io_dmem_s1_kill_0_REG_34 : _GEN_98780) : _GEN_98780;
  wire        _GEN_988 = do_ld_search_1 & stq_0_valid & lcam_st_dep_mask_1[0];
  wire [7:0]  _GEN_989 = casez_tmp_109 & casez_tmp_144;
  wire        _GEN_99430 = _GEN_989 == casez_tmp_109 & ~stq_0_bits_uop_is_fence & ~stq_0_bits_uop_is_amo & dword_addr_matches_32_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_32;
  wire        _GEN_990 = (|_GEN_989) & dword_addr_matches_32_1;
  reg         io_dmem_s1_kill_1_REG_33;
  reg         io_dmem_s1_kill_1_REG_34;
  wire        _GEN_99466 = _GEN_988 ? (_GEN_99430 ? io_dmem_s1_kill_1_REG_32 : _GEN_990 ? io_dmem_s1_kill_1_REG_33 : _GEN_99361 ? io_dmem_s1_kill_1_REG_34 : _GEN_99029) : _GEN_99029;
  wire        dword_addr_matches_33_0 = stq_1_bits_addr_valid & ~stq_1_bits_addr_is_virtual & stq_1_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_33_1 = stq_1_bits_addr_valid & ~stq_1_bits_addr_is_virtual & stq_1_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_17 = 15'h1 << stq_1_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_21 = 15'h3 << {12'h0, stq_1_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_1_bits_uop_mem_size)
      2'b00:
        casez_tmp_145 = _write_mask_mask_T_17[7:0];
      2'b01:
        casez_tmp_145 = _write_mask_mask_T_21[7:0];
      2'b10:
        casez_tmp_145 = stq_1_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_145 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_991 = _do_ld_search_T_2 & stq_1_valid & lcam_st_dep_mask_0[1];
  wire [7:0]  _GEN_992 = casez_tmp_108 & casez_tmp_145;
  wire        _GEN_99664 = _GEN_992 == casez_tmp_108 & ~stq_1_bits_uop_is_fence & ~stq_1_bits_uop_is_amo & dword_addr_matches_33_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_35;
  wire        _GEN_993 = (|_GEN_992) & dword_addr_matches_33_0;
  reg         io_dmem_s1_kill_0_REG_36;
  wire        _GEN_99829 = stq_1_bits_uop_is_fence | stq_1_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_37;
  wire        _GEN_99700 = _GEN_991 ? (_GEN_99664 ? io_dmem_s1_kill_0_REG_35 : _GEN_993 ? io_dmem_s1_kill_0_REG_36 : _GEN_99829 ? io_dmem_s1_kill_0_REG_37 : _GEN_99232) : _GEN_99232;
  wire        _GEN_994 = do_ld_search_1 & stq_1_valid & lcam_st_dep_mask_1[1];
  wire [7:0]  _GEN_995 = casez_tmp_109 & casez_tmp_145;
  wire        _GEN_99898 = _GEN_995 == casez_tmp_109 & ~stq_1_bits_uop_is_fence & ~stq_1_bits_uop_is_amo & dword_addr_matches_33_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_35;
  wire        _GEN_996 = (|_GEN_995) & dword_addr_matches_33_1;
  reg         io_dmem_s1_kill_1_REG_36;
  reg         io_dmem_s1_kill_1_REG_37;
  wire        _GEN_99934 = _GEN_994 ? (_GEN_99898 ? io_dmem_s1_kill_1_REG_35 : _GEN_996 ? io_dmem_s1_kill_1_REG_36 : _GEN_99829 ? io_dmem_s1_kill_1_REG_37 : _GEN_99466) : _GEN_99466;
  wire        dword_addr_matches_34_0 = stq_2_bits_addr_valid & ~stq_2_bits_addr_is_virtual & stq_2_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_34_1 = stq_2_bits_addr_valid & ~stq_2_bits_addr_is_virtual & stq_2_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_32 = 15'h1 << stq_2_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_36 = 15'h3 << {12'h0, stq_2_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_2_bits_uop_mem_size)
      2'b00:
        casez_tmp_146 = _write_mask_mask_T_32[7:0];
      2'b01:
        casez_tmp_146 = _write_mask_mask_T_36[7:0];
      2'b10:
        casez_tmp_146 = stq_2_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_146 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_997 = _do_ld_search_T_2 & stq_2_valid & lcam_st_dep_mask_0[2];
  wire [7:0]  _GEN_998 = casez_tmp_108 & casez_tmp_146;
  wire        _GEN_100132 = _GEN_998 == casez_tmp_108 & ~stq_2_bits_uop_is_fence & ~stq_2_bits_uop_is_amo & dword_addr_matches_34_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_38;
  wire        _GEN_999 = (|_GEN_998) & dword_addr_matches_34_0;
  reg         io_dmem_s1_kill_0_REG_39;
  wire        _GEN_100297 = stq_2_bits_uop_is_fence | stq_2_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_40;
  wire        _GEN_100168 = _GEN_997 ? (_GEN_100132 ? io_dmem_s1_kill_0_REG_38 : _GEN_999 ? io_dmem_s1_kill_0_REG_39 : _GEN_100297 ? io_dmem_s1_kill_0_REG_40 : _GEN_99700) : _GEN_99700;
  wire        _GEN_1000 = do_ld_search_1 & stq_2_valid & lcam_st_dep_mask_1[2];
  wire [7:0]  _GEN_1001 = casez_tmp_109 & casez_tmp_146;
  wire        _GEN_100366 = _GEN_1001 == casez_tmp_109 & ~stq_2_bits_uop_is_fence & ~stq_2_bits_uop_is_amo & dword_addr_matches_34_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_38;
  wire        _GEN_1002 = (|_GEN_1001) & dword_addr_matches_34_1;
  reg         io_dmem_s1_kill_1_REG_39;
  reg         io_dmem_s1_kill_1_REG_40;
  wire        _GEN_100402 = _GEN_1000 ? (_GEN_100366 ? io_dmem_s1_kill_1_REG_38 : _GEN_1002 ? io_dmem_s1_kill_1_REG_39 : _GEN_100297 ? io_dmem_s1_kill_1_REG_40 : _GEN_99934) : _GEN_99934;
  wire        dword_addr_matches_35_0 = stq_3_bits_addr_valid & ~stq_3_bits_addr_is_virtual & stq_3_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_35_1 = stq_3_bits_addr_valid & ~stq_3_bits_addr_is_virtual & stq_3_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_47 = 15'h1 << stq_3_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_51 = 15'h3 << {12'h0, stq_3_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_3_bits_uop_mem_size)
      2'b00:
        casez_tmp_147 = _write_mask_mask_T_47[7:0];
      2'b01:
        casez_tmp_147 = _write_mask_mask_T_51[7:0];
      2'b10:
        casez_tmp_147 = stq_3_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_147 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1003 = _do_ld_search_T_2 & stq_3_valid & lcam_st_dep_mask_0[3];
  wire [7:0]  _GEN_1004 = casez_tmp_108 & casez_tmp_147;
  wire        _GEN_100600 = _GEN_1004 == casez_tmp_108 & ~stq_3_bits_uop_is_fence & ~stq_3_bits_uop_is_amo & dword_addr_matches_35_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_41;
  wire        _GEN_1005 = (|_GEN_1004) & dword_addr_matches_35_0;
  reg         io_dmem_s1_kill_0_REG_42;
  wire        _GEN_100765 = stq_3_bits_uop_is_fence | stq_3_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_43;
  wire        _GEN_100636 = _GEN_1003 ? (_GEN_100600 ? io_dmem_s1_kill_0_REG_41 : _GEN_1005 ? io_dmem_s1_kill_0_REG_42 : _GEN_100765 ? io_dmem_s1_kill_0_REG_43 : _GEN_100168) : _GEN_100168;
  wire        _GEN_1006 = do_ld_search_1 & stq_3_valid & lcam_st_dep_mask_1[3];
  wire [7:0]  _GEN_1007 = casez_tmp_109 & casez_tmp_147;
  wire        _GEN_100834 = _GEN_1007 == casez_tmp_109 & ~stq_3_bits_uop_is_fence & ~stq_3_bits_uop_is_amo & dword_addr_matches_35_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_41;
  wire        _GEN_1008 = (|_GEN_1007) & dword_addr_matches_35_1;
  reg         io_dmem_s1_kill_1_REG_42;
  reg         io_dmem_s1_kill_1_REG_43;
  wire        _GEN_100870 = _GEN_1006 ? (_GEN_100834 ? io_dmem_s1_kill_1_REG_41 : _GEN_1008 ? io_dmem_s1_kill_1_REG_42 : _GEN_100765 ? io_dmem_s1_kill_1_REG_43 : _GEN_100402) : _GEN_100402;
  wire        dword_addr_matches_36_0 = stq_4_bits_addr_valid & ~stq_4_bits_addr_is_virtual & stq_4_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_36_1 = stq_4_bits_addr_valid & ~stq_4_bits_addr_is_virtual & stq_4_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_62 = 15'h1 << stq_4_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_66 = 15'h3 << {12'h0, stq_4_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_4_bits_uop_mem_size)
      2'b00:
        casez_tmp_148 = _write_mask_mask_T_62[7:0];
      2'b01:
        casez_tmp_148 = _write_mask_mask_T_66[7:0];
      2'b10:
        casez_tmp_148 = stq_4_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_148 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1009 = _do_ld_search_T_2 & stq_4_valid & lcam_st_dep_mask_0[4];
  wire [7:0]  _GEN_1010 = casez_tmp_108 & casez_tmp_148;
  wire        _GEN_101068 = _GEN_1010 == casez_tmp_108 & ~stq_4_bits_uop_is_fence & ~stq_4_bits_uop_is_amo & dword_addr_matches_36_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_44;
  wire        _GEN_1011 = (|_GEN_1010) & dword_addr_matches_36_0;
  reg         io_dmem_s1_kill_0_REG_45;
  wire        _GEN_101233 = stq_4_bits_uop_is_fence | stq_4_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_46;
  wire        _GEN_101104 = _GEN_1009 ? (_GEN_101068 ? io_dmem_s1_kill_0_REG_44 : _GEN_1011 ? io_dmem_s1_kill_0_REG_45 : _GEN_101233 ? io_dmem_s1_kill_0_REG_46 : _GEN_100636) : _GEN_100636;
  wire        _GEN_1012 = do_ld_search_1 & stq_4_valid & lcam_st_dep_mask_1[4];
  wire [7:0]  _GEN_1013 = casez_tmp_109 & casez_tmp_148;
  wire        _GEN_101302 = _GEN_1013 == casez_tmp_109 & ~stq_4_bits_uop_is_fence & ~stq_4_bits_uop_is_amo & dword_addr_matches_36_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_44;
  wire        _GEN_1014 = (|_GEN_1013) & dword_addr_matches_36_1;
  reg         io_dmem_s1_kill_1_REG_45;
  reg         io_dmem_s1_kill_1_REG_46;
  wire        _GEN_101338 = _GEN_1012 ? (_GEN_101302 ? io_dmem_s1_kill_1_REG_44 : _GEN_1014 ? io_dmem_s1_kill_1_REG_45 : _GEN_101233 ? io_dmem_s1_kill_1_REG_46 : _GEN_100870) : _GEN_100870;
  wire        dword_addr_matches_37_0 = stq_5_bits_addr_valid & ~stq_5_bits_addr_is_virtual & stq_5_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_37_1 = stq_5_bits_addr_valid & ~stq_5_bits_addr_is_virtual & stq_5_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_77 = 15'h1 << stq_5_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_81 = 15'h3 << {12'h0, stq_5_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_5_bits_uop_mem_size)
      2'b00:
        casez_tmp_149 = _write_mask_mask_T_77[7:0];
      2'b01:
        casez_tmp_149 = _write_mask_mask_T_81[7:0];
      2'b10:
        casez_tmp_149 = stq_5_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_149 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1015 = _do_ld_search_T_2 & stq_5_valid & lcam_st_dep_mask_0[5];
  wire [7:0]  _GEN_1016 = casez_tmp_108 & casez_tmp_149;
  wire        _GEN_101536 = _GEN_1016 == casez_tmp_108 & ~stq_5_bits_uop_is_fence & ~stq_5_bits_uop_is_amo & dword_addr_matches_37_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_47;
  wire        _GEN_1017 = (|_GEN_1016) & dword_addr_matches_37_0;
  reg         io_dmem_s1_kill_0_REG_48;
  wire        _GEN_101701 = stq_5_bits_uop_is_fence | stq_5_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_49;
  wire        _GEN_101572 = _GEN_1015 ? (_GEN_101536 ? io_dmem_s1_kill_0_REG_47 : _GEN_1017 ? io_dmem_s1_kill_0_REG_48 : _GEN_101701 ? io_dmem_s1_kill_0_REG_49 : _GEN_101104) : _GEN_101104;
  wire        _GEN_1018 = do_ld_search_1 & stq_5_valid & lcam_st_dep_mask_1[5];
  wire [7:0]  _GEN_1019 = casez_tmp_109 & casez_tmp_149;
  wire        _GEN_101770 = _GEN_1019 == casez_tmp_109 & ~stq_5_bits_uop_is_fence & ~stq_5_bits_uop_is_amo & dword_addr_matches_37_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_47;
  wire        _GEN_1020 = (|_GEN_1019) & dword_addr_matches_37_1;
  reg         io_dmem_s1_kill_1_REG_48;
  reg         io_dmem_s1_kill_1_REG_49;
  wire        _GEN_101806 = _GEN_1018 ? (_GEN_101770 ? io_dmem_s1_kill_1_REG_47 : _GEN_1020 ? io_dmem_s1_kill_1_REG_48 : _GEN_101701 ? io_dmem_s1_kill_1_REG_49 : _GEN_101338) : _GEN_101338;
  wire        dword_addr_matches_38_0 = stq_6_bits_addr_valid & ~stq_6_bits_addr_is_virtual & stq_6_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_38_1 = stq_6_bits_addr_valid & ~stq_6_bits_addr_is_virtual & stq_6_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_92 = 15'h1 << stq_6_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_96 = 15'h3 << {12'h0, stq_6_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_6_bits_uop_mem_size)
      2'b00:
        casez_tmp_150 = _write_mask_mask_T_92[7:0];
      2'b01:
        casez_tmp_150 = _write_mask_mask_T_96[7:0];
      2'b10:
        casez_tmp_150 = stq_6_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_150 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1021 = _do_ld_search_T_2 & stq_6_valid & lcam_st_dep_mask_0[6];
  wire [7:0]  _GEN_1022 = casez_tmp_108 & casez_tmp_150;
  wire        _GEN_102004 = _GEN_1022 == casez_tmp_108 & ~stq_6_bits_uop_is_fence & ~stq_6_bits_uop_is_amo & dword_addr_matches_38_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_50;
  wire        _GEN_1023 = (|_GEN_1022) & dword_addr_matches_38_0;
  reg         io_dmem_s1_kill_0_REG_51;
  wire        _GEN_102169 = stq_6_bits_uop_is_fence | stq_6_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_52;
  wire        _GEN_102040 = _GEN_1021 ? (_GEN_102004 ? io_dmem_s1_kill_0_REG_50 : _GEN_1023 ? io_dmem_s1_kill_0_REG_51 : _GEN_102169 ? io_dmem_s1_kill_0_REG_52 : _GEN_101572) : _GEN_101572;
  wire        _GEN_1024 = do_ld_search_1 & stq_6_valid & lcam_st_dep_mask_1[6];
  wire [7:0]  _GEN_1025 = casez_tmp_109 & casez_tmp_150;
  wire        _GEN_102238 = _GEN_1025 == casez_tmp_109 & ~stq_6_bits_uop_is_fence & ~stq_6_bits_uop_is_amo & dword_addr_matches_38_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_50;
  wire        _GEN_1026 = (|_GEN_1025) & dword_addr_matches_38_1;
  reg         io_dmem_s1_kill_1_REG_51;
  reg         io_dmem_s1_kill_1_REG_52;
  wire        _GEN_102274 = _GEN_1024 ? (_GEN_102238 ? io_dmem_s1_kill_1_REG_50 : _GEN_1026 ? io_dmem_s1_kill_1_REG_51 : _GEN_102169 ? io_dmem_s1_kill_1_REG_52 : _GEN_101806) : _GEN_101806;
  wire        dword_addr_matches_39_0 = stq_7_bits_addr_valid & ~stq_7_bits_addr_is_virtual & stq_7_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_39_1 = stq_7_bits_addr_valid & ~stq_7_bits_addr_is_virtual & stq_7_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_107 = 15'h1 << stq_7_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_111 = 15'h3 << {12'h0, stq_7_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_7_bits_uop_mem_size)
      2'b00:
        casez_tmp_151 = _write_mask_mask_T_107[7:0];
      2'b01:
        casez_tmp_151 = _write_mask_mask_T_111[7:0];
      2'b10:
        casez_tmp_151 = stq_7_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_151 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1027 = _do_ld_search_T_2 & stq_7_valid & lcam_st_dep_mask_0[7];
  wire [7:0]  _GEN_1028 = casez_tmp_108 & casez_tmp_151;
  wire        _GEN_102472 = _GEN_1028 == casez_tmp_108 & ~stq_7_bits_uop_is_fence & ~stq_7_bits_uop_is_amo & dword_addr_matches_39_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_53;
  wire        _GEN_1029 = (|_GEN_1028) & dword_addr_matches_39_0;
  reg         io_dmem_s1_kill_0_REG_54;
  wire        _GEN_102637 = stq_7_bits_uop_is_fence | stq_7_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_55;
  wire        _GEN_102508 = _GEN_1027 ? (_GEN_102472 ? io_dmem_s1_kill_0_REG_53 : _GEN_1029 ? io_dmem_s1_kill_0_REG_54 : _GEN_102637 ? io_dmem_s1_kill_0_REG_55 : _GEN_102040) : _GEN_102040;
  wire        _GEN_1030 = do_ld_search_1 & stq_7_valid & lcam_st_dep_mask_1[7];
  wire [7:0]  _GEN_1031 = casez_tmp_109 & casez_tmp_151;
  wire        _GEN_102706 = _GEN_1031 == casez_tmp_109 & ~stq_7_bits_uop_is_fence & ~stq_7_bits_uop_is_amo & dword_addr_matches_39_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_53;
  wire        _GEN_1032 = (|_GEN_1031) & dword_addr_matches_39_1;
  reg         io_dmem_s1_kill_1_REG_54;
  reg         io_dmem_s1_kill_1_REG_55;
  wire        _GEN_102742 = _GEN_1030 ? (_GEN_102706 ? io_dmem_s1_kill_1_REG_53 : _GEN_1032 ? io_dmem_s1_kill_1_REG_54 : _GEN_102637 ? io_dmem_s1_kill_1_REG_55 : _GEN_102274) : _GEN_102274;
  wire        dword_addr_matches_40_0 = stq_8_bits_addr_valid & ~stq_8_bits_addr_is_virtual & stq_8_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_40_1 = stq_8_bits_addr_valid & ~stq_8_bits_addr_is_virtual & stq_8_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_122 = 15'h1 << stq_8_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_126 = 15'h3 << {12'h0, stq_8_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_8_bits_uop_mem_size)
      2'b00:
        casez_tmp_152 = _write_mask_mask_T_122[7:0];
      2'b01:
        casez_tmp_152 = _write_mask_mask_T_126[7:0];
      2'b10:
        casez_tmp_152 = stq_8_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_152 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1033 = _do_ld_search_T_2 & stq_8_valid & lcam_st_dep_mask_0[8];
  wire [7:0]  _GEN_1034 = casez_tmp_108 & casez_tmp_152;
  wire        _GEN_102940 = _GEN_1034 == casez_tmp_108 & ~stq_8_bits_uop_is_fence & ~stq_8_bits_uop_is_amo & dword_addr_matches_40_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_56;
  wire        _GEN_1035 = (|_GEN_1034) & dword_addr_matches_40_0;
  reg         io_dmem_s1_kill_0_REG_57;
  wire        _GEN_103105 = stq_8_bits_uop_is_fence | stq_8_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_58;
  wire        _GEN_102976 = _GEN_1033 ? (_GEN_102940 ? io_dmem_s1_kill_0_REG_56 : _GEN_1035 ? io_dmem_s1_kill_0_REG_57 : _GEN_103105 ? io_dmem_s1_kill_0_REG_58 : _GEN_102508) : _GEN_102508;
  wire        _GEN_1036 = do_ld_search_1 & stq_8_valid & lcam_st_dep_mask_1[8];
  wire [7:0]  _GEN_1037 = casez_tmp_109 & casez_tmp_152;
  wire        _GEN_103174 = _GEN_1037 == casez_tmp_109 & ~stq_8_bits_uop_is_fence & ~stq_8_bits_uop_is_amo & dword_addr_matches_40_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_56;
  wire        _GEN_1038 = (|_GEN_1037) & dword_addr_matches_40_1;
  reg         io_dmem_s1_kill_1_REG_57;
  reg         io_dmem_s1_kill_1_REG_58;
  wire        _GEN_103210 = _GEN_1036 ? (_GEN_103174 ? io_dmem_s1_kill_1_REG_56 : _GEN_1038 ? io_dmem_s1_kill_1_REG_57 : _GEN_103105 ? io_dmem_s1_kill_1_REG_58 : _GEN_102742) : _GEN_102742;
  wire        dword_addr_matches_41_0 = stq_9_bits_addr_valid & ~stq_9_bits_addr_is_virtual & stq_9_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_41_1 = stq_9_bits_addr_valid & ~stq_9_bits_addr_is_virtual & stq_9_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_137 = 15'h1 << stq_9_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_141 = 15'h3 << {12'h0, stq_9_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_9_bits_uop_mem_size)
      2'b00:
        casez_tmp_153 = _write_mask_mask_T_137[7:0];
      2'b01:
        casez_tmp_153 = _write_mask_mask_T_141[7:0];
      2'b10:
        casez_tmp_153 = stq_9_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_153 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1039 = _do_ld_search_T_2 & stq_9_valid & lcam_st_dep_mask_0[9];
  wire [7:0]  _GEN_1040 = casez_tmp_108 & casez_tmp_153;
  wire        _GEN_103408 = _GEN_1040 == casez_tmp_108 & ~stq_9_bits_uop_is_fence & ~stq_9_bits_uop_is_amo & dword_addr_matches_41_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_59;
  wire        _GEN_1041 = (|_GEN_1040) & dword_addr_matches_41_0;
  reg         io_dmem_s1_kill_0_REG_60;
  wire        _GEN_103573 = stq_9_bits_uop_is_fence | stq_9_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_61;
  wire        _GEN_103444 = _GEN_1039 ? (_GEN_103408 ? io_dmem_s1_kill_0_REG_59 : _GEN_1041 ? io_dmem_s1_kill_0_REG_60 : _GEN_103573 ? io_dmem_s1_kill_0_REG_61 : _GEN_102976) : _GEN_102976;
  wire        _GEN_1042 = do_ld_search_1 & stq_9_valid & lcam_st_dep_mask_1[9];
  wire [7:0]  _GEN_1043 = casez_tmp_109 & casez_tmp_153;
  wire        _GEN_103642 = _GEN_1043 == casez_tmp_109 & ~stq_9_bits_uop_is_fence & ~stq_9_bits_uop_is_amo & dword_addr_matches_41_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_59;
  wire        _GEN_1044 = (|_GEN_1043) & dword_addr_matches_41_1;
  reg         io_dmem_s1_kill_1_REG_60;
  reg         io_dmem_s1_kill_1_REG_61;
  wire        _GEN_103678 = _GEN_1042 ? (_GEN_103642 ? io_dmem_s1_kill_1_REG_59 : _GEN_1044 ? io_dmem_s1_kill_1_REG_60 : _GEN_103573 ? io_dmem_s1_kill_1_REG_61 : _GEN_103210) : _GEN_103210;
  wire        dword_addr_matches_42_0 = stq_10_bits_addr_valid & ~stq_10_bits_addr_is_virtual & stq_10_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_42_1 = stq_10_bits_addr_valid & ~stq_10_bits_addr_is_virtual & stq_10_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_152 = 15'h1 << stq_10_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_156 = 15'h3 << {12'h0, stq_10_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_10_bits_uop_mem_size)
      2'b00:
        casez_tmp_154 = _write_mask_mask_T_152[7:0];
      2'b01:
        casez_tmp_154 = _write_mask_mask_T_156[7:0];
      2'b10:
        casez_tmp_154 = stq_10_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_154 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1045 = _do_ld_search_T_2 & stq_10_valid & lcam_st_dep_mask_0[10];
  wire [7:0]  _GEN_1046 = casez_tmp_108 & casez_tmp_154;
  wire        _GEN_103876 = _GEN_1046 == casez_tmp_108 & ~stq_10_bits_uop_is_fence & ~stq_10_bits_uop_is_amo & dword_addr_matches_42_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_62;
  wire        _GEN_1047 = (|_GEN_1046) & dword_addr_matches_42_0;
  reg         io_dmem_s1_kill_0_REG_63;
  wire        _GEN_104041 = stq_10_bits_uop_is_fence | stq_10_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_64;
  wire        _GEN_103912 = _GEN_1045 ? (_GEN_103876 ? io_dmem_s1_kill_0_REG_62 : _GEN_1047 ? io_dmem_s1_kill_0_REG_63 : _GEN_104041 ? io_dmem_s1_kill_0_REG_64 : _GEN_103444) : _GEN_103444;
  wire        _GEN_1048 = do_ld_search_1 & stq_10_valid & lcam_st_dep_mask_1[10];
  wire [7:0]  _GEN_1049 = casez_tmp_109 & casez_tmp_154;
  wire        _GEN_104110 = _GEN_1049 == casez_tmp_109 & ~stq_10_bits_uop_is_fence & ~stq_10_bits_uop_is_amo & dword_addr_matches_42_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_62;
  wire        _GEN_1050 = (|_GEN_1049) & dword_addr_matches_42_1;
  reg         io_dmem_s1_kill_1_REG_63;
  reg         io_dmem_s1_kill_1_REG_64;
  wire        _GEN_104146 = _GEN_1048 ? (_GEN_104110 ? io_dmem_s1_kill_1_REG_62 : _GEN_1050 ? io_dmem_s1_kill_1_REG_63 : _GEN_104041 ? io_dmem_s1_kill_1_REG_64 : _GEN_103678) : _GEN_103678;
  wire        dword_addr_matches_43_0 = stq_11_bits_addr_valid & ~stq_11_bits_addr_is_virtual & stq_11_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_43_1 = stq_11_bits_addr_valid & ~stq_11_bits_addr_is_virtual & stq_11_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_167 = 15'h1 << stq_11_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_171 = 15'h3 << {12'h0, stq_11_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_11_bits_uop_mem_size)
      2'b00:
        casez_tmp_155 = _write_mask_mask_T_167[7:0];
      2'b01:
        casez_tmp_155 = _write_mask_mask_T_171[7:0];
      2'b10:
        casez_tmp_155 = stq_11_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_155 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1051 = _do_ld_search_T_2 & stq_11_valid & lcam_st_dep_mask_0[11];
  wire [7:0]  _GEN_1052 = casez_tmp_108 & casez_tmp_155;
  wire        _GEN_104344 = _GEN_1052 == casez_tmp_108 & ~stq_11_bits_uop_is_fence & ~stq_11_bits_uop_is_amo & dword_addr_matches_43_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_65;
  wire        _GEN_1053 = (|_GEN_1052) & dword_addr_matches_43_0;
  reg         io_dmem_s1_kill_0_REG_66;
  wire        _GEN_104509 = stq_11_bits_uop_is_fence | stq_11_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_67;
  wire        _GEN_104380 = _GEN_1051 ? (_GEN_104344 ? io_dmem_s1_kill_0_REG_65 : _GEN_1053 ? io_dmem_s1_kill_0_REG_66 : _GEN_104509 ? io_dmem_s1_kill_0_REG_67 : _GEN_103912) : _GEN_103912;
  wire        _GEN_1054 = do_ld_search_1 & stq_11_valid & lcam_st_dep_mask_1[11];
  wire [7:0]  _GEN_1055 = casez_tmp_109 & casez_tmp_155;
  wire        _GEN_104578 = _GEN_1055 == casez_tmp_109 & ~stq_11_bits_uop_is_fence & ~stq_11_bits_uop_is_amo & dword_addr_matches_43_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_65;
  wire        _GEN_1056 = (|_GEN_1055) & dword_addr_matches_43_1;
  reg         io_dmem_s1_kill_1_REG_66;
  reg         io_dmem_s1_kill_1_REG_67;
  wire        _GEN_104614 = _GEN_1054 ? (_GEN_104578 ? io_dmem_s1_kill_1_REG_65 : _GEN_1056 ? io_dmem_s1_kill_1_REG_66 : _GEN_104509 ? io_dmem_s1_kill_1_REG_67 : _GEN_104146) : _GEN_104146;
  wire        dword_addr_matches_44_0 = stq_12_bits_addr_valid & ~stq_12_bits_addr_is_virtual & stq_12_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_44_1 = stq_12_bits_addr_valid & ~stq_12_bits_addr_is_virtual & stq_12_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_182 = 15'h1 << stq_12_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_186 = 15'h3 << {12'h0, stq_12_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_12_bits_uop_mem_size)
      2'b00:
        casez_tmp_156 = _write_mask_mask_T_182[7:0];
      2'b01:
        casez_tmp_156 = _write_mask_mask_T_186[7:0];
      2'b10:
        casez_tmp_156 = stq_12_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_156 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1057 = _do_ld_search_T_2 & stq_12_valid & lcam_st_dep_mask_0[12];
  wire [7:0]  _GEN_1058 = casez_tmp_108 & casez_tmp_156;
  wire        _GEN_104812 = _GEN_1058 == casez_tmp_108 & ~stq_12_bits_uop_is_fence & ~stq_12_bits_uop_is_amo & dword_addr_matches_44_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_68;
  wire        _GEN_1059 = (|_GEN_1058) & dword_addr_matches_44_0;
  reg         io_dmem_s1_kill_0_REG_69;
  wire        _GEN_104977 = stq_12_bits_uop_is_fence | stq_12_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_70;
  wire        _GEN_104848 = _GEN_1057 ? (_GEN_104812 ? io_dmem_s1_kill_0_REG_68 : _GEN_1059 ? io_dmem_s1_kill_0_REG_69 : _GEN_104977 ? io_dmem_s1_kill_0_REG_70 : _GEN_104380) : _GEN_104380;
  wire        _GEN_1060 = do_ld_search_1 & stq_12_valid & lcam_st_dep_mask_1[12];
  wire [7:0]  _GEN_1061 = casez_tmp_109 & casez_tmp_156;
  wire        _GEN_105046 = _GEN_1061 == casez_tmp_109 & ~stq_12_bits_uop_is_fence & ~stq_12_bits_uop_is_amo & dword_addr_matches_44_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_68;
  wire        _GEN_1062 = (|_GEN_1061) & dword_addr_matches_44_1;
  reg         io_dmem_s1_kill_1_REG_69;
  reg         io_dmem_s1_kill_1_REG_70;
  wire        _GEN_105082 = _GEN_1060 ? (_GEN_105046 ? io_dmem_s1_kill_1_REG_68 : _GEN_1062 ? io_dmem_s1_kill_1_REG_69 : _GEN_104977 ? io_dmem_s1_kill_1_REG_70 : _GEN_104614) : _GEN_104614;
  wire        dword_addr_matches_45_0 = stq_13_bits_addr_valid & ~stq_13_bits_addr_is_virtual & stq_13_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_45_1 = stq_13_bits_addr_valid & ~stq_13_bits_addr_is_virtual & stq_13_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_197 = 15'h1 << stq_13_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_201 = 15'h3 << {12'h0, stq_13_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_13_bits_uop_mem_size)
      2'b00:
        casez_tmp_157 = _write_mask_mask_T_197[7:0];
      2'b01:
        casez_tmp_157 = _write_mask_mask_T_201[7:0];
      2'b10:
        casez_tmp_157 = stq_13_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_157 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1063 = _do_ld_search_T_2 & stq_13_valid & lcam_st_dep_mask_0[13];
  wire [7:0]  _GEN_1064 = casez_tmp_108 & casez_tmp_157;
  wire        _GEN_105280 = _GEN_1064 == casez_tmp_108 & ~stq_13_bits_uop_is_fence & ~stq_13_bits_uop_is_amo & dword_addr_matches_45_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_71;
  wire        _GEN_1065 = (|_GEN_1064) & dword_addr_matches_45_0;
  reg         io_dmem_s1_kill_0_REG_72;
  wire        _GEN_105445 = stq_13_bits_uop_is_fence | stq_13_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_73;
  wire        _GEN_105316 = _GEN_1063 ? (_GEN_105280 ? io_dmem_s1_kill_0_REG_71 : _GEN_1065 ? io_dmem_s1_kill_0_REG_72 : _GEN_105445 ? io_dmem_s1_kill_0_REG_73 : _GEN_104848) : _GEN_104848;
  wire        _GEN_1066 = do_ld_search_1 & stq_13_valid & lcam_st_dep_mask_1[13];
  wire [7:0]  _GEN_1067 = casez_tmp_109 & casez_tmp_157;
  wire        _GEN_105514 = _GEN_1067 == casez_tmp_109 & ~stq_13_bits_uop_is_fence & ~stq_13_bits_uop_is_amo & dword_addr_matches_45_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_71;
  wire        _GEN_1068 = (|_GEN_1067) & dword_addr_matches_45_1;
  reg         io_dmem_s1_kill_1_REG_72;
  reg         io_dmem_s1_kill_1_REG_73;
  wire        _GEN_105550 = _GEN_1066 ? (_GEN_105514 ? io_dmem_s1_kill_1_REG_71 : _GEN_1068 ? io_dmem_s1_kill_1_REG_72 : _GEN_105445 ? io_dmem_s1_kill_1_REG_73 : _GEN_105082) : _GEN_105082;
  wire        dword_addr_matches_46_0 = stq_14_bits_addr_valid & ~stq_14_bits_addr_is_virtual & stq_14_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_46_1 = stq_14_bits_addr_valid & ~stq_14_bits_addr_is_virtual & stq_14_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_212 = 15'h1 << stq_14_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_216 = 15'h3 << {12'h0, stq_14_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_14_bits_uop_mem_size)
      2'b00:
        casez_tmp_158 = _write_mask_mask_T_212[7:0];
      2'b01:
        casez_tmp_158 = _write_mask_mask_T_216[7:0];
      2'b10:
        casez_tmp_158 = stq_14_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_158 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1069 = _do_ld_search_T_2 & stq_14_valid & lcam_st_dep_mask_0[14];
  wire [7:0]  _GEN_1070 = casez_tmp_108 & casez_tmp_158;
  wire        _GEN_105748 = _GEN_1070 == casez_tmp_108 & ~stq_14_bits_uop_is_fence & ~stq_14_bits_uop_is_amo & dword_addr_matches_46_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_74;
  wire        _GEN_1071 = (|_GEN_1070) & dword_addr_matches_46_0;
  reg         io_dmem_s1_kill_0_REG_75;
  wire        _GEN_105913 = stq_14_bits_uop_is_fence | stq_14_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_76;
  wire        _GEN_105784 = _GEN_1069 ? (_GEN_105748 ? io_dmem_s1_kill_0_REG_74 : _GEN_1071 ? io_dmem_s1_kill_0_REG_75 : _GEN_105913 ? io_dmem_s1_kill_0_REG_76 : _GEN_105316) : _GEN_105316;
  wire        _GEN_1072 = do_ld_search_1 & stq_14_valid & lcam_st_dep_mask_1[14];
  wire [7:0]  _GEN_1073 = casez_tmp_109 & casez_tmp_158;
  wire        _GEN_105982 = _GEN_1073 == casez_tmp_109 & ~stq_14_bits_uop_is_fence & ~stq_14_bits_uop_is_amo & dword_addr_matches_46_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_74;
  wire        _GEN_1074 = (|_GEN_1073) & dword_addr_matches_46_1;
  reg         io_dmem_s1_kill_1_REG_75;
  reg         io_dmem_s1_kill_1_REG_76;
  wire        _GEN_106018 = _GEN_1072 ? (_GEN_105982 ? io_dmem_s1_kill_1_REG_74 : _GEN_1074 ? io_dmem_s1_kill_1_REG_75 : _GEN_105913 ? io_dmem_s1_kill_1_REG_76 : _GEN_105550) : _GEN_105550;
  wire        dword_addr_matches_47_0 = stq_15_bits_addr_valid & ~stq_15_bits_addr_is_virtual & stq_15_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_47_1 = stq_15_bits_addr_valid & ~stq_15_bits_addr_is_virtual & stq_15_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_227 = 15'h1 << stq_15_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_231 = 15'h3 << {12'h0, stq_15_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_15_bits_uop_mem_size)
      2'b00:
        casez_tmp_159 = _write_mask_mask_T_227[7:0];
      2'b01:
        casez_tmp_159 = _write_mask_mask_T_231[7:0];
      2'b10:
        casez_tmp_159 = stq_15_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_159 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1075 = _do_ld_search_T_2 & stq_15_valid & lcam_st_dep_mask_0[15];
  wire [7:0]  _GEN_1076 = casez_tmp_108 & casez_tmp_159;
  wire        _GEN_106216 = _GEN_1076 == casez_tmp_108 & ~stq_15_bits_uop_is_fence & ~stq_15_bits_uop_is_amo & dword_addr_matches_47_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_77;
  wire        _GEN_1077 = (|_GEN_1076) & dword_addr_matches_47_0;
  reg         io_dmem_s1_kill_0_REG_78;
  wire        _GEN_106381 = stq_15_bits_uop_is_fence | stq_15_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_79;
  wire        _GEN_106252 = _GEN_1075 ? (_GEN_106216 ? io_dmem_s1_kill_0_REG_77 : _GEN_1077 ? io_dmem_s1_kill_0_REG_78 : _GEN_106381 ? io_dmem_s1_kill_0_REG_79 : _GEN_105784) : _GEN_105784;
  wire        _GEN_1078 = do_ld_search_1 & stq_15_valid & lcam_st_dep_mask_1[15];
  wire [7:0]  _GEN_1079 = casez_tmp_109 & casez_tmp_159;
  wire        _GEN_106450 = _GEN_1079 == casez_tmp_109 & ~stq_15_bits_uop_is_fence & ~stq_15_bits_uop_is_amo & dword_addr_matches_47_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_77;
  wire        _GEN_1080 = (|_GEN_1079) & dword_addr_matches_47_1;
  reg         io_dmem_s1_kill_1_REG_78;
  reg         io_dmem_s1_kill_1_REG_79;
  wire        _GEN_106486 = _GEN_1078 ? (_GEN_106450 ? io_dmem_s1_kill_1_REG_77 : _GEN_1080 ? io_dmem_s1_kill_1_REG_78 : _GEN_106381 ? io_dmem_s1_kill_1_REG_79 : _GEN_106018) : _GEN_106018;
  wire        dword_addr_matches_48_0 = stq_16_bits_addr_valid & ~stq_16_bits_addr_is_virtual & stq_16_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_48_1 = stq_16_bits_addr_valid & ~stq_16_bits_addr_is_virtual & stq_16_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_242 = 15'h1 << stq_16_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_246 = 15'h3 << {12'h0, stq_16_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_16_bits_uop_mem_size)
      2'b00:
        casez_tmp_160 = _write_mask_mask_T_242[7:0];
      2'b01:
        casez_tmp_160 = _write_mask_mask_T_246[7:0];
      2'b10:
        casez_tmp_160 = stq_16_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_160 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1081 = _do_ld_search_T_2 & stq_16_valid & lcam_st_dep_mask_0[16];
  wire [7:0]  _GEN_1082 = casez_tmp_108 & casez_tmp_160;
  wire        _GEN_106684 = _GEN_1082 == casez_tmp_108 & ~stq_16_bits_uop_is_fence & ~stq_16_bits_uop_is_amo & dword_addr_matches_48_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_80;
  wire        _GEN_1083 = (|_GEN_1082) & dword_addr_matches_48_0;
  reg         io_dmem_s1_kill_0_REG_81;
  wire        _GEN_106849 = stq_16_bits_uop_is_fence | stq_16_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_82;
  wire        _GEN_106720 = _GEN_1081 ? (_GEN_106684 ? io_dmem_s1_kill_0_REG_80 : _GEN_1083 ? io_dmem_s1_kill_0_REG_81 : _GEN_106849 ? io_dmem_s1_kill_0_REG_82 : _GEN_106252) : _GEN_106252;
  wire        _GEN_1084 = do_ld_search_1 & stq_16_valid & lcam_st_dep_mask_1[16];
  wire [7:0]  _GEN_1085 = casez_tmp_109 & casez_tmp_160;
  wire        _GEN_106918 = _GEN_1085 == casez_tmp_109 & ~stq_16_bits_uop_is_fence & ~stq_16_bits_uop_is_amo & dword_addr_matches_48_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_80;
  wire        _GEN_1086 = (|_GEN_1085) & dword_addr_matches_48_1;
  reg         io_dmem_s1_kill_1_REG_81;
  reg         io_dmem_s1_kill_1_REG_82;
  wire        _GEN_106954 = _GEN_1084 ? (_GEN_106918 ? io_dmem_s1_kill_1_REG_80 : _GEN_1086 ? io_dmem_s1_kill_1_REG_81 : _GEN_106849 ? io_dmem_s1_kill_1_REG_82 : _GEN_106486) : _GEN_106486;
  wire        dword_addr_matches_49_0 = stq_17_bits_addr_valid & ~stq_17_bits_addr_is_virtual & stq_17_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_49_1 = stq_17_bits_addr_valid & ~stq_17_bits_addr_is_virtual & stq_17_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_257 = 15'h1 << stq_17_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_261 = 15'h3 << {12'h0, stq_17_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_17_bits_uop_mem_size)
      2'b00:
        casez_tmp_161 = _write_mask_mask_T_257[7:0];
      2'b01:
        casez_tmp_161 = _write_mask_mask_T_261[7:0];
      2'b10:
        casez_tmp_161 = stq_17_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_161 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1087 = _do_ld_search_T_2 & stq_17_valid & lcam_st_dep_mask_0[17];
  wire [7:0]  _GEN_1088 = casez_tmp_108 & casez_tmp_161;
  wire        _GEN_107152 = _GEN_1088 == casez_tmp_108 & ~stq_17_bits_uop_is_fence & ~stq_17_bits_uop_is_amo & dword_addr_matches_49_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_83;
  wire        _GEN_1089 = (|_GEN_1088) & dword_addr_matches_49_0;
  reg         io_dmem_s1_kill_0_REG_84;
  wire        _GEN_107317 = stq_17_bits_uop_is_fence | stq_17_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_85;
  wire        _GEN_107188 = _GEN_1087 ? (_GEN_107152 ? io_dmem_s1_kill_0_REG_83 : _GEN_1089 ? io_dmem_s1_kill_0_REG_84 : _GEN_107317 ? io_dmem_s1_kill_0_REG_85 : _GEN_106720) : _GEN_106720;
  wire        _GEN_1090 = do_ld_search_1 & stq_17_valid & lcam_st_dep_mask_1[17];
  wire [7:0]  _GEN_1091 = casez_tmp_109 & casez_tmp_161;
  wire        _GEN_107386 = _GEN_1091 == casez_tmp_109 & ~stq_17_bits_uop_is_fence & ~stq_17_bits_uop_is_amo & dword_addr_matches_49_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_83;
  wire        _GEN_1092 = (|_GEN_1091) & dword_addr_matches_49_1;
  reg         io_dmem_s1_kill_1_REG_84;
  reg         io_dmem_s1_kill_1_REG_85;
  wire        _GEN_107422 = _GEN_1090 ? (_GEN_107386 ? io_dmem_s1_kill_1_REG_83 : _GEN_1092 ? io_dmem_s1_kill_1_REG_84 : _GEN_107317 ? io_dmem_s1_kill_1_REG_85 : _GEN_106954) : _GEN_106954;
  wire        dword_addr_matches_50_0 = stq_18_bits_addr_valid & ~stq_18_bits_addr_is_virtual & stq_18_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_50_1 = stq_18_bits_addr_valid & ~stq_18_bits_addr_is_virtual & stq_18_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_272 = 15'h1 << stq_18_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_276 = 15'h3 << {12'h0, stq_18_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_18_bits_uop_mem_size)
      2'b00:
        casez_tmp_162 = _write_mask_mask_T_272[7:0];
      2'b01:
        casez_tmp_162 = _write_mask_mask_T_276[7:0];
      2'b10:
        casez_tmp_162 = stq_18_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_162 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1093 = _do_ld_search_T_2 & stq_18_valid & lcam_st_dep_mask_0[18];
  wire [7:0]  _GEN_1094 = casez_tmp_108 & casez_tmp_162;
  wire        _GEN_107620 = _GEN_1094 == casez_tmp_108 & ~stq_18_bits_uop_is_fence & ~stq_18_bits_uop_is_amo & dword_addr_matches_50_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_86;
  wire        _GEN_1095 = (|_GEN_1094) & dword_addr_matches_50_0;
  reg         io_dmem_s1_kill_0_REG_87;
  wire        _GEN_107785 = stq_18_bits_uop_is_fence | stq_18_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_88;
  wire        _GEN_107656 = _GEN_1093 ? (_GEN_107620 ? io_dmem_s1_kill_0_REG_86 : _GEN_1095 ? io_dmem_s1_kill_0_REG_87 : _GEN_107785 ? io_dmem_s1_kill_0_REG_88 : _GEN_107188) : _GEN_107188;
  wire        _GEN_1096 = do_ld_search_1 & stq_18_valid & lcam_st_dep_mask_1[18];
  wire [7:0]  _GEN_1097 = casez_tmp_109 & casez_tmp_162;
  wire        _GEN_107854 = _GEN_1097 == casez_tmp_109 & ~stq_18_bits_uop_is_fence & ~stq_18_bits_uop_is_amo & dword_addr_matches_50_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_86;
  wire        _GEN_1098 = (|_GEN_1097) & dword_addr_matches_50_1;
  reg         io_dmem_s1_kill_1_REG_87;
  reg         io_dmem_s1_kill_1_REG_88;
  wire        _GEN_107890 = _GEN_1096 ? (_GEN_107854 ? io_dmem_s1_kill_1_REG_86 : _GEN_1098 ? io_dmem_s1_kill_1_REG_87 : _GEN_107785 ? io_dmem_s1_kill_1_REG_88 : _GEN_107422) : _GEN_107422;
  wire        dword_addr_matches_51_0 = stq_19_bits_addr_valid & ~stq_19_bits_addr_is_virtual & stq_19_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_51_1 = stq_19_bits_addr_valid & ~stq_19_bits_addr_is_virtual & stq_19_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_287 = 15'h1 << stq_19_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_291 = 15'h3 << {12'h0, stq_19_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_19_bits_uop_mem_size)
      2'b00:
        casez_tmp_163 = _write_mask_mask_T_287[7:0];
      2'b01:
        casez_tmp_163 = _write_mask_mask_T_291[7:0];
      2'b10:
        casez_tmp_163 = stq_19_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_163 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1099 = _do_ld_search_T_2 & stq_19_valid & lcam_st_dep_mask_0[19];
  wire [7:0]  _GEN_1100 = casez_tmp_108 & casez_tmp_163;
  wire        _GEN_108088 = _GEN_1100 == casez_tmp_108 & ~stq_19_bits_uop_is_fence & ~stq_19_bits_uop_is_amo & dword_addr_matches_51_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_89;
  wire        _GEN_1101 = (|_GEN_1100) & dword_addr_matches_51_0;
  reg         io_dmem_s1_kill_0_REG_90;
  wire        _GEN_108253 = stq_19_bits_uop_is_fence | stq_19_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_91;
  wire        _GEN_108124 = _GEN_1099 ? (_GEN_108088 ? io_dmem_s1_kill_0_REG_89 : _GEN_1101 ? io_dmem_s1_kill_0_REG_90 : _GEN_108253 ? io_dmem_s1_kill_0_REG_91 : _GEN_107656) : _GEN_107656;
  wire        _GEN_1102 = do_ld_search_1 & stq_19_valid & lcam_st_dep_mask_1[19];
  wire [7:0]  _GEN_1103 = casez_tmp_109 & casez_tmp_163;
  wire        _GEN_108322 = _GEN_1103 == casez_tmp_109 & ~stq_19_bits_uop_is_fence & ~stq_19_bits_uop_is_amo & dword_addr_matches_51_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_89;
  wire        _GEN_1104 = (|_GEN_1103) & dword_addr_matches_51_1;
  reg         io_dmem_s1_kill_1_REG_90;
  reg         io_dmem_s1_kill_1_REG_91;
  wire        _GEN_108358 = _GEN_1102 ? (_GEN_108322 ? io_dmem_s1_kill_1_REG_89 : _GEN_1104 ? io_dmem_s1_kill_1_REG_90 : _GEN_108253 ? io_dmem_s1_kill_1_REG_91 : _GEN_107890) : _GEN_107890;
  wire        dword_addr_matches_52_0 = stq_20_bits_addr_valid & ~stq_20_bits_addr_is_virtual & stq_20_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_52_1 = stq_20_bits_addr_valid & ~stq_20_bits_addr_is_virtual & stq_20_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_302 = 15'h1 << stq_20_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_306 = 15'h3 << {12'h0, stq_20_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_20_bits_uop_mem_size)
      2'b00:
        casez_tmp_164 = _write_mask_mask_T_302[7:0];
      2'b01:
        casez_tmp_164 = _write_mask_mask_T_306[7:0];
      2'b10:
        casez_tmp_164 = stq_20_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_164 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1105 = _do_ld_search_T_2 & stq_20_valid & lcam_st_dep_mask_0[20];
  wire [7:0]  _GEN_1106 = casez_tmp_108 & casez_tmp_164;
  wire        _GEN_108556 = _GEN_1106 == casez_tmp_108 & ~stq_20_bits_uop_is_fence & ~stq_20_bits_uop_is_amo & dword_addr_matches_52_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_92;
  wire        _GEN_1107 = (|_GEN_1106) & dword_addr_matches_52_0;
  reg         io_dmem_s1_kill_0_REG_93;
  wire        _GEN_108721 = stq_20_bits_uop_is_fence | stq_20_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_94;
  wire        _GEN_108592 = _GEN_1105 ? (_GEN_108556 ? io_dmem_s1_kill_0_REG_92 : _GEN_1107 ? io_dmem_s1_kill_0_REG_93 : _GEN_108721 ? io_dmem_s1_kill_0_REG_94 : _GEN_108124) : _GEN_108124;
  wire        _GEN_1108 = do_ld_search_1 & stq_20_valid & lcam_st_dep_mask_1[20];
  wire [7:0]  _GEN_1109 = casez_tmp_109 & casez_tmp_164;
  wire        _GEN_108790 = _GEN_1109 == casez_tmp_109 & ~stq_20_bits_uop_is_fence & ~stq_20_bits_uop_is_amo & dword_addr_matches_52_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_92;
  wire        _GEN_1110 = (|_GEN_1109) & dword_addr_matches_52_1;
  reg         io_dmem_s1_kill_1_REG_93;
  reg         io_dmem_s1_kill_1_REG_94;
  wire        _GEN_108826 = _GEN_1108 ? (_GEN_108790 ? io_dmem_s1_kill_1_REG_92 : _GEN_1110 ? io_dmem_s1_kill_1_REG_93 : _GEN_108721 ? io_dmem_s1_kill_1_REG_94 : _GEN_108358) : _GEN_108358;
  wire        dword_addr_matches_53_0 = stq_21_bits_addr_valid & ~stq_21_bits_addr_is_virtual & stq_21_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_53_1 = stq_21_bits_addr_valid & ~stq_21_bits_addr_is_virtual & stq_21_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_317 = 15'h1 << stq_21_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_321 = 15'h3 << {12'h0, stq_21_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_21_bits_uop_mem_size)
      2'b00:
        casez_tmp_165 = _write_mask_mask_T_317[7:0];
      2'b01:
        casez_tmp_165 = _write_mask_mask_T_321[7:0];
      2'b10:
        casez_tmp_165 = stq_21_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_165 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1111 = _do_ld_search_T_2 & stq_21_valid & lcam_st_dep_mask_0[21];
  wire [7:0]  _GEN_1112 = casez_tmp_108 & casez_tmp_165;
  wire        _GEN_109024 = _GEN_1112 == casez_tmp_108 & ~stq_21_bits_uop_is_fence & ~stq_21_bits_uop_is_amo & dword_addr_matches_53_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_95;
  wire        _GEN_1113 = (|_GEN_1112) & dword_addr_matches_53_0;
  reg         io_dmem_s1_kill_0_REG_96;
  wire        _GEN_109189 = stq_21_bits_uop_is_fence | stq_21_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_97;
  wire        _GEN_109060 = _GEN_1111 ? (_GEN_109024 ? io_dmem_s1_kill_0_REG_95 : _GEN_1113 ? io_dmem_s1_kill_0_REG_96 : _GEN_109189 ? io_dmem_s1_kill_0_REG_97 : _GEN_108592) : _GEN_108592;
  wire        _GEN_1114 = do_ld_search_1 & stq_21_valid & lcam_st_dep_mask_1[21];
  wire [7:0]  _GEN_1115 = casez_tmp_109 & casez_tmp_165;
  wire        _GEN_109258 = _GEN_1115 == casez_tmp_109 & ~stq_21_bits_uop_is_fence & ~stq_21_bits_uop_is_amo & dword_addr_matches_53_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_95;
  wire        _GEN_1116 = (|_GEN_1115) & dword_addr_matches_53_1;
  reg         io_dmem_s1_kill_1_REG_96;
  reg         io_dmem_s1_kill_1_REG_97;
  wire        _GEN_109294 = _GEN_1114 ? (_GEN_109258 ? io_dmem_s1_kill_1_REG_95 : _GEN_1116 ? io_dmem_s1_kill_1_REG_96 : _GEN_109189 ? io_dmem_s1_kill_1_REG_97 : _GEN_108826) : _GEN_108826;
  wire        dword_addr_matches_54_0 = stq_22_bits_addr_valid & ~stq_22_bits_addr_is_virtual & stq_22_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_54_1 = stq_22_bits_addr_valid & ~stq_22_bits_addr_is_virtual & stq_22_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_332 = 15'h1 << stq_22_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_336 = 15'h3 << {12'h0, stq_22_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_22_bits_uop_mem_size)
      2'b00:
        casez_tmp_166 = _write_mask_mask_T_332[7:0];
      2'b01:
        casez_tmp_166 = _write_mask_mask_T_336[7:0];
      2'b10:
        casez_tmp_166 = stq_22_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_166 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1117 = _do_ld_search_T_2 & stq_22_valid & lcam_st_dep_mask_0[22];
  wire [7:0]  _GEN_1118 = casez_tmp_108 & casez_tmp_166;
  wire        _GEN_109492 = _GEN_1118 == casez_tmp_108 & ~stq_22_bits_uop_is_fence & ~stq_22_bits_uop_is_amo & dword_addr_matches_54_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_98;
  wire        _GEN_1119 = (|_GEN_1118) & dword_addr_matches_54_0;
  reg         io_dmem_s1_kill_0_REG_99;
  wire        _GEN_109657 = stq_22_bits_uop_is_fence | stq_22_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_100;
  wire        _GEN_109528 = _GEN_1117 ? (_GEN_109492 ? io_dmem_s1_kill_0_REG_98 : _GEN_1119 ? io_dmem_s1_kill_0_REG_99 : _GEN_109657 ? io_dmem_s1_kill_0_REG_100 : _GEN_109060) : _GEN_109060;
  wire        _GEN_1120 = do_ld_search_1 & stq_22_valid & lcam_st_dep_mask_1[22];
  wire [7:0]  _GEN_1121 = casez_tmp_109 & casez_tmp_166;
  wire        _GEN_109726 = _GEN_1121 == casez_tmp_109 & ~stq_22_bits_uop_is_fence & ~stq_22_bits_uop_is_amo & dword_addr_matches_54_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_98;
  wire        _GEN_1122 = (|_GEN_1121) & dword_addr_matches_54_1;
  reg         io_dmem_s1_kill_1_REG_99;
  reg         io_dmem_s1_kill_1_REG_100;
  wire        _GEN_109762 = _GEN_1120 ? (_GEN_109726 ? io_dmem_s1_kill_1_REG_98 : _GEN_1122 ? io_dmem_s1_kill_1_REG_99 : _GEN_109657 ? io_dmem_s1_kill_1_REG_100 : _GEN_109294) : _GEN_109294;
  wire        dword_addr_matches_55_0 = stq_23_bits_addr_valid & ~stq_23_bits_addr_is_virtual & stq_23_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_55_1 = stq_23_bits_addr_valid & ~stq_23_bits_addr_is_virtual & stq_23_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_347 = 15'h1 << stq_23_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_351 = 15'h3 << {12'h0, stq_23_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_23_bits_uop_mem_size)
      2'b00:
        casez_tmp_167 = _write_mask_mask_T_347[7:0];
      2'b01:
        casez_tmp_167 = _write_mask_mask_T_351[7:0];
      2'b10:
        casez_tmp_167 = stq_23_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_167 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1123 = _do_ld_search_T_2 & stq_23_valid & lcam_st_dep_mask_0[23];
  wire [7:0]  _GEN_1124 = casez_tmp_108 & casez_tmp_167;
  wire        _GEN_109960 = _GEN_1124 == casez_tmp_108 & ~stq_23_bits_uop_is_fence & ~stq_23_bits_uop_is_amo & dword_addr_matches_55_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_101;
  wire        _GEN_1125 = (|_GEN_1124) & dword_addr_matches_55_0;
  reg         io_dmem_s1_kill_0_REG_102;
  wire        _GEN_110125 = stq_23_bits_uop_is_fence | stq_23_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_103;
  wire        _GEN_109996 = _GEN_1123 ? (_GEN_109960 ? io_dmem_s1_kill_0_REG_101 : _GEN_1125 ? io_dmem_s1_kill_0_REG_102 : _GEN_110125 ? io_dmem_s1_kill_0_REG_103 : _GEN_109528) : _GEN_109528;
  wire        _GEN_1126 = do_ld_search_1 & stq_23_valid & lcam_st_dep_mask_1[23];
  wire [7:0]  _GEN_1127 = casez_tmp_109 & casez_tmp_167;
  wire        _GEN_110194 = _GEN_1127 == casez_tmp_109 & ~stq_23_bits_uop_is_fence & ~stq_23_bits_uop_is_amo & dword_addr_matches_55_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_101;
  wire        _GEN_1128 = (|_GEN_1127) & dword_addr_matches_55_1;
  reg         io_dmem_s1_kill_1_REG_102;
  reg         io_dmem_s1_kill_1_REG_103;
  wire        _GEN_110230 = _GEN_1126 ? (_GEN_110194 ? io_dmem_s1_kill_1_REG_101 : _GEN_1128 ? io_dmem_s1_kill_1_REG_102 : _GEN_110125 ? io_dmem_s1_kill_1_REG_103 : _GEN_109762) : _GEN_109762;
  wire        dword_addr_matches_56_0 = stq_24_bits_addr_valid & ~stq_24_bits_addr_is_virtual & stq_24_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_56_1 = stq_24_bits_addr_valid & ~stq_24_bits_addr_is_virtual & stq_24_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_362 = 15'h1 << stq_24_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_366 = 15'h3 << {12'h0, stq_24_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_24_bits_uop_mem_size)
      2'b00:
        casez_tmp_168 = _write_mask_mask_T_362[7:0];
      2'b01:
        casez_tmp_168 = _write_mask_mask_T_366[7:0];
      2'b10:
        casez_tmp_168 = stq_24_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_168 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1129 = _do_ld_search_T_2 & stq_24_valid & lcam_st_dep_mask_0[24];
  wire [7:0]  _GEN_1130 = casez_tmp_108 & casez_tmp_168;
  wire        _GEN_110428 = _GEN_1130 == casez_tmp_108 & ~stq_24_bits_uop_is_fence & ~stq_24_bits_uop_is_amo & dword_addr_matches_56_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_104;
  wire        _GEN_1131 = (|_GEN_1130) & dword_addr_matches_56_0;
  reg         io_dmem_s1_kill_0_REG_105;
  wire        _GEN_110593 = stq_24_bits_uop_is_fence | stq_24_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_106;
  wire        _GEN_110464 = _GEN_1129 ? (_GEN_110428 ? io_dmem_s1_kill_0_REG_104 : _GEN_1131 ? io_dmem_s1_kill_0_REG_105 : _GEN_110593 ? io_dmem_s1_kill_0_REG_106 : _GEN_109996) : _GEN_109996;
  wire        _GEN_1132 = do_ld_search_1 & stq_24_valid & lcam_st_dep_mask_1[24];
  wire [7:0]  _GEN_1133 = casez_tmp_109 & casez_tmp_168;
  wire        _GEN_110662 = _GEN_1133 == casez_tmp_109 & ~stq_24_bits_uop_is_fence & ~stq_24_bits_uop_is_amo & dword_addr_matches_56_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_104;
  wire        _GEN_1134 = (|_GEN_1133) & dword_addr_matches_56_1;
  reg         io_dmem_s1_kill_1_REG_105;
  reg         io_dmem_s1_kill_1_REG_106;
  wire        _GEN_110698 = _GEN_1132 ? (_GEN_110662 ? io_dmem_s1_kill_1_REG_104 : _GEN_1134 ? io_dmem_s1_kill_1_REG_105 : _GEN_110593 ? io_dmem_s1_kill_1_REG_106 : _GEN_110230) : _GEN_110230;
  wire        dword_addr_matches_57_0 = stq_25_bits_addr_valid & ~stq_25_bits_addr_is_virtual & stq_25_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_57_1 = stq_25_bits_addr_valid & ~stq_25_bits_addr_is_virtual & stq_25_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_377 = 15'h1 << stq_25_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_381 = 15'h3 << {12'h0, stq_25_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_25_bits_uop_mem_size)
      2'b00:
        casez_tmp_169 = _write_mask_mask_T_377[7:0];
      2'b01:
        casez_tmp_169 = _write_mask_mask_T_381[7:0];
      2'b10:
        casez_tmp_169 = stq_25_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_169 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1135 = _do_ld_search_T_2 & stq_25_valid & lcam_st_dep_mask_0[25];
  wire [7:0]  _GEN_1136 = casez_tmp_108 & casez_tmp_169;
  wire        _GEN_110896 = _GEN_1136 == casez_tmp_108 & ~stq_25_bits_uop_is_fence & ~stq_25_bits_uop_is_amo & dword_addr_matches_57_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_107;
  wire        _GEN_1137 = (|_GEN_1136) & dword_addr_matches_57_0;
  reg         io_dmem_s1_kill_0_REG_108;
  wire        _GEN_111061 = stq_25_bits_uop_is_fence | stq_25_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_109;
  wire        _GEN_110932 = _GEN_1135 ? (_GEN_110896 ? io_dmem_s1_kill_0_REG_107 : _GEN_1137 ? io_dmem_s1_kill_0_REG_108 : _GEN_111061 ? io_dmem_s1_kill_0_REG_109 : _GEN_110464) : _GEN_110464;
  wire        _GEN_1138 = do_ld_search_1 & stq_25_valid & lcam_st_dep_mask_1[25];
  wire [7:0]  _GEN_1139 = casez_tmp_109 & casez_tmp_169;
  wire        _GEN_111130 = _GEN_1139 == casez_tmp_109 & ~stq_25_bits_uop_is_fence & ~stq_25_bits_uop_is_amo & dword_addr_matches_57_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_107;
  wire        _GEN_1140 = (|_GEN_1139) & dword_addr_matches_57_1;
  reg         io_dmem_s1_kill_1_REG_108;
  reg         io_dmem_s1_kill_1_REG_109;
  wire        _GEN_111166 = _GEN_1138 ? (_GEN_111130 ? io_dmem_s1_kill_1_REG_107 : _GEN_1140 ? io_dmem_s1_kill_1_REG_108 : _GEN_111061 ? io_dmem_s1_kill_1_REG_109 : _GEN_110698) : _GEN_110698;
  wire        dword_addr_matches_58_0 = stq_26_bits_addr_valid & ~stq_26_bits_addr_is_virtual & stq_26_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_58_1 = stq_26_bits_addr_valid & ~stq_26_bits_addr_is_virtual & stq_26_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_392 = 15'h1 << stq_26_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_396 = 15'h3 << {12'h0, stq_26_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_26_bits_uop_mem_size)
      2'b00:
        casez_tmp_170 = _write_mask_mask_T_392[7:0];
      2'b01:
        casez_tmp_170 = _write_mask_mask_T_396[7:0];
      2'b10:
        casez_tmp_170 = stq_26_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_170 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1141 = _do_ld_search_T_2 & stq_26_valid & lcam_st_dep_mask_0[26];
  wire [7:0]  _GEN_1142 = casez_tmp_108 & casez_tmp_170;
  wire        _GEN_111364 = _GEN_1142 == casez_tmp_108 & ~stq_26_bits_uop_is_fence & ~stq_26_bits_uop_is_amo & dword_addr_matches_58_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_110;
  wire        _GEN_1143 = (|_GEN_1142) & dword_addr_matches_58_0;
  reg         io_dmem_s1_kill_0_REG_111;
  wire        _GEN_111529 = stq_26_bits_uop_is_fence | stq_26_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_112;
  wire        _GEN_111400 = _GEN_1141 ? (_GEN_111364 ? io_dmem_s1_kill_0_REG_110 : _GEN_1143 ? io_dmem_s1_kill_0_REG_111 : _GEN_111529 ? io_dmem_s1_kill_0_REG_112 : _GEN_110932) : _GEN_110932;
  wire        _GEN_1144 = do_ld_search_1 & stq_26_valid & lcam_st_dep_mask_1[26];
  wire [7:0]  _GEN_1145 = casez_tmp_109 & casez_tmp_170;
  wire        _GEN_111598 = _GEN_1145 == casez_tmp_109 & ~stq_26_bits_uop_is_fence & ~stq_26_bits_uop_is_amo & dword_addr_matches_58_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_110;
  wire        _GEN_1146 = (|_GEN_1145) & dword_addr_matches_58_1;
  reg         io_dmem_s1_kill_1_REG_111;
  reg         io_dmem_s1_kill_1_REG_112;
  wire        _GEN_111634 = _GEN_1144 ? (_GEN_111598 ? io_dmem_s1_kill_1_REG_110 : _GEN_1146 ? io_dmem_s1_kill_1_REG_111 : _GEN_111529 ? io_dmem_s1_kill_1_REG_112 : _GEN_111166) : _GEN_111166;
  wire        dword_addr_matches_59_0 = stq_27_bits_addr_valid & ~stq_27_bits_addr_is_virtual & stq_27_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_59_1 = stq_27_bits_addr_valid & ~stq_27_bits_addr_is_virtual & stq_27_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_407 = 15'h1 << stq_27_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_411 = 15'h3 << {12'h0, stq_27_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_27_bits_uop_mem_size)
      2'b00:
        casez_tmp_171 = _write_mask_mask_T_407[7:0];
      2'b01:
        casez_tmp_171 = _write_mask_mask_T_411[7:0];
      2'b10:
        casez_tmp_171 = stq_27_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_171 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1147 = _do_ld_search_T_2 & stq_27_valid & lcam_st_dep_mask_0[27];
  wire [7:0]  _GEN_1148 = casez_tmp_108 & casez_tmp_171;
  wire        _GEN_111832 = _GEN_1148 == casez_tmp_108 & ~stq_27_bits_uop_is_fence & ~stq_27_bits_uop_is_amo & dword_addr_matches_59_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_113;
  wire        _GEN_1149 = (|_GEN_1148) & dword_addr_matches_59_0;
  reg         io_dmem_s1_kill_0_REG_114;
  wire        _GEN_111997 = stq_27_bits_uop_is_fence | stq_27_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_115;
  wire        _GEN_111868 = _GEN_1147 ? (_GEN_111832 ? io_dmem_s1_kill_0_REG_113 : _GEN_1149 ? io_dmem_s1_kill_0_REG_114 : _GEN_111997 ? io_dmem_s1_kill_0_REG_115 : _GEN_111400) : _GEN_111400;
  wire        _GEN_1150 = do_ld_search_1 & stq_27_valid & lcam_st_dep_mask_1[27];
  wire [7:0]  _GEN_1151 = casez_tmp_109 & casez_tmp_171;
  wire        _GEN_112066 = _GEN_1151 == casez_tmp_109 & ~stq_27_bits_uop_is_fence & ~stq_27_bits_uop_is_amo & dword_addr_matches_59_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_113;
  wire        _GEN_1152 = (|_GEN_1151) & dword_addr_matches_59_1;
  reg         io_dmem_s1_kill_1_REG_114;
  reg         io_dmem_s1_kill_1_REG_115;
  wire        _GEN_112102 = _GEN_1150 ? (_GEN_112066 ? io_dmem_s1_kill_1_REG_113 : _GEN_1152 ? io_dmem_s1_kill_1_REG_114 : _GEN_111997 ? io_dmem_s1_kill_1_REG_115 : _GEN_111634) : _GEN_111634;
  wire        dword_addr_matches_60_0 = stq_28_bits_addr_valid & ~stq_28_bits_addr_is_virtual & stq_28_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_60_1 = stq_28_bits_addr_valid & ~stq_28_bits_addr_is_virtual & stq_28_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_422 = 15'h1 << stq_28_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_426 = 15'h3 << {12'h0, stq_28_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_28_bits_uop_mem_size)
      2'b00:
        casez_tmp_172 = _write_mask_mask_T_422[7:0];
      2'b01:
        casez_tmp_172 = _write_mask_mask_T_426[7:0];
      2'b10:
        casez_tmp_172 = stq_28_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_172 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1153 = _do_ld_search_T_2 & stq_28_valid & lcam_st_dep_mask_0[28];
  wire [7:0]  _GEN_1154 = casez_tmp_108 & casez_tmp_172;
  wire        _GEN_112300 = _GEN_1154 == casez_tmp_108 & ~stq_28_bits_uop_is_fence & ~stq_28_bits_uop_is_amo & dword_addr_matches_60_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_116;
  wire        _GEN_1155 = (|_GEN_1154) & dword_addr_matches_60_0;
  reg         io_dmem_s1_kill_0_REG_117;
  wire        _GEN_112465 = stq_28_bits_uop_is_fence | stq_28_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_118;
  wire        _GEN_112336 = _GEN_1153 ? (_GEN_112300 ? io_dmem_s1_kill_0_REG_116 : _GEN_1155 ? io_dmem_s1_kill_0_REG_117 : _GEN_112465 ? io_dmem_s1_kill_0_REG_118 : _GEN_111868) : _GEN_111868;
  wire        _GEN_1156 = do_ld_search_1 & stq_28_valid & lcam_st_dep_mask_1[28];
  wire [7:0]  _GEN_1157 = casez_tmp_109 & casez_tmp_172;
  wire        _GEN_112534 = _GEN_1157 == casez_tmp_109 & ~stq_28_bits_uop_is_fence & ~stq_28_bits_uop_is_amo & dword_addr_matches_60_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_116;
  wire        _GEN_1158 = (|_GEN_1157) & dword_addr_matches_60_1;
  reg         io_dmem_s1_kill_1_REG_117;
  reg         io_dmem_s1_kill_1_REG_118;
  wire        _GEN_112570 = _GEN_1156 ? (_GEN_112534 ? io_dmem_s1_kill_1_REG_116 : _GEN_1158 ? io_dmem_s1_kill_1_REG_117 : _GEN_112465 ? io_dmem_s1_kill_1_REG_118 : _GEN_112102) : _GEN_112102;
  wire        dword_addr_matches_61_0 = stq_29_bits_addr_valid & ~stq_29_bits_addr_is_virtual & stq_29_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_61_1 = stq_29_bits_addr_valid & ~stq_29_bits_addr_is_virtual & stq_29_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_437 = 15'h1 << stq_29_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_441 = 15'h3 << {12'h0, stq_29_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_29_bits_uop_mem_size)
      2'b00:
        casez_tmp_173 = _write_mask_mask_T_437[7:0];
      2'b01:
        casez_tmp_173 = _write_mask_mask_T_441[7:0];
      2'b10:
        casez_tmp_173 = stq_29_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_173 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1159 = _do_ld_search_T_2 & stq_29_valid & lcam_st_dep_mask_0[29];
  wire [7:0]  _GEN_1160 = casez_tmp_108 & casez_tmp_173;
  wire        _GEN_112768 = _GEN_1160 == casez_tmp_108 & ~stq_29_bits_uop_is_fence & ~stq_29_bits_uop_is_amo & dword_addr_matches_61_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_119;
  wire        _GEN_1161 = (|_GEN_1160) & dword_addr_matches_61_0;
  reg         io_dmem_s1_kill_0_REG_120;
  wire        _GEN_112933 = stq_29_bits_uop_is_fence | stq_29_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_121;
  wire        _GEN_112804 = _GEN_1159 ? (_GEN_112768 ? io_dmem_s1_kill_0_REG_119 : _GEN_1161 ? io_dmem_s1_kill_0_REG_120 : _GEN_112933 ? io_dmem_s1_kill_0_REG_121 : _GEN_112336) : _GEN_112336;
  wire        _GEN_1162 = do_ld_search_1 & stq_29_valid & lcam_st_dep_mask_1[29];
  wire [7:0]  _GEN_1163 = casez_tmp_109 & casez_tmp_173;
  wire        _GEN_113002 = _GEN_1163 == casez_tmp_109 & ~stq_29_bits_uop_is_fence & ~stq_29_bits_uop_is_amo & dword_addr_matches_61_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_119;
  wire        _GEN_1164 = (|_GEN_1163) & dword_addr_matches_61_1;
  reg         io_dmem_s1_kill_1_REG_120;
  reg         io_dmem_s1_kill_1_REG_121;
  wire        _GEN_113038 = _GEN_1162 ? (_GEN_113002 ? io_dmem_s1_kill_1_REG_119 : _GEN_1164 ? io_dmem_s1_kill_1_REG_120 : _GEN_112933 ? io_dmem_s1_kill_1_REG_121 : _GEN_112570) : _GEN_112570;
  wire        dword_addr_matches_62_0 = stq_30_bits_addr_valid & ~stq_30_bits_addr_is_virtual & stq_30_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_62_1 = stq_30_bits_addr_valid & ~stq_30_bits_addr_is_virtual & stq_30_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_452 = 15'h1 << stq_30_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_456 = 15'h3 << {12'h0, stq_30_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_30_bits_uop_mem_size)
      2'b00:
        casez_tmp_174 = _write_mask_mask_T_452[7:0];
      2'b01:
        casez_tmp_174 = _write_mask_mask_T_456[7:0];
      2'b10:
        casez_tmp_174 = stq_30_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_174 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1165 = _do_ld_search_T_2 & stq_30_valid & lcam_st_dep_mask_0[30];
  wire [7:0]  _GEN_1166 = casez_tmp_108 & casez_tmp_174;
  wire        _GEN_113236 = _GEN_1166 == casez_tmp_108 & ~stq_30_bits_uop_is_fence & ~stq_30_bits_uop_is_amo & dword_addr_matches_62_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_122;
  wire        _GEN_1167 = (|_GEN_1166) & dword_addr_matches_62_0;
  reg         io_dmem_s1_kill_0_REG_123;
  wire        _GEN_113401 = stq_30_bits_uop_is_fence | stq_30_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_124;
  wire        _GEN_113272 = _GEN_1165 ? (_GEN_113236 ? io_dmem_s1_kill_0_REG_122 : _GEN_1167 ? io_dmem_s1_kill_0_REG_123 : _GEN_113401 ? io_dmem_s1_kill_0_REG_124 : _GEN_112804) : _GEN_112804;
  wire        _GEN_1168 = do_ld_search_1 & stq_30_valid & lcam_st_dep_mask_1[30];
  wire [7:0]  _GEN_1169 = casez_tmp_109 & casez_tmp_174;
  wire        _GEN_113470 = _GEN_1169 == casez_tmp_109 & ~stq_30_bits_uop_is_fence & ~stq_30_bits_uop_is_amo & dword_addr_matches_62_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_122;
  wire        _GEN_1170 = (|_GEN_1169) & dword_addr_matches_62_1;
  reg         io_dmem_s1_kill_1_REG_123;
  reg         io_dmem_s1_kill_1_REG_124;
  wire        _GEN_113506 = _GEN_1168 ? (_GEN_113470 ? io_dmem_s1_kill_1_REG_122 : _GEN_1170 ? io_dmem_s1_kill_1_REG_123 : _GEN_113401 ? io_dmem_s1_kill_1_REG_124 : _GEN_113038) : _GEN_113038;
  wire        dword_addr_matches_63_0 = stq_31_bits_addr_valid & ~stq_31_bits_addr_is_virtual & stq_31_bits_addr_bits[31:3] == lcam_addr_0[31:3];
  wire        dword_addr_matches_63_1 = stq_31_bits_addr_valid & ~stq_31_bits_addr_is_virtual & stq_31_bits_addr_bits[31:3] == lcam_addr_1[31:3];
  wire [14:0] _write_mask_mask_T_467 = 15'h1 << stq_31_bits_addr_bits[2:0];
  wire [14:0] _write_mask_mask_T_471 = 15'h3 << {12'h0, stq_31_bits_addr_bits[2:1], 1'h0};
  always @(*) begin
    casez (stq_31_bits_uop_mem_size)
      2'b00:
        casez_tmp_175 = _write_mask_mask_T_467[7:0];
      2'b01:
        casez_tmp_175 = _write_mask_mask_T_471[7:0];
      2'b10:
        casez_tmp_175 = stq_31_bits_addr_bits[2] ? 8'hF0 : 8'hF;
      default:
        casez_tmp_175 = 8'hFF;
    endcase
  end // always @(*)
  wire        _GEN_1171 = _do_ld_search_T_2 & stq_31_valid & lcam_st_dep_mask_0[31];
  wire [7:0]  _GEN_1172 = casez_tmp_108 & casez_tmp_175;
  wire        _GEN_113704 = _GEN_1172 == casez_tmp_108 & ~stq_31_bits_uop_is_fence & ~stq_31_bits_uop_is_amo & dword_addr_matches_63_0 & can_forward_0;
  reg         io_dmem_s1_kill_0_REG_125;
  wire        _GEN_1173 = (|_GEN_1172) & dword_addr_matches_63_0;
  reg         io_dmem_s1_kill_0_REG_126;
  wire        _GEN_113869 = stq_31_bits_uop_is_fence | stq_31_bits_uop_is_amo;
  reg         io_dmem_s1_kill_0_REG_127;
  wire        _GEN_1174 = do_ld_search_1 & stq_31_valid & lcam_st_dep_mask_1[31];
  wire [7:0]  _GEN_1175 = casez_tmp_109 & casez_tmp_175;
  wire        _GEN_113938 = _GEN_1175 == casez_tmp_109 & ~stq_31_bits_uop_is_fence & ~stq_31_bits_uop_is_amo & dword_addr_matches_63_1 & can_forward_1;
  reg         io_dmem_s1_kill_1_REG_125;
  wire        _GEN_1176 = (|_GEN_1175) & dword_addr_matches_63_1;
  reg         io_dmem_s1_kill_1_REG_126;
  reg         io_dmem_s1_kill_1_REG_127;
  always @(*) begin
    casez (_forwarding_age_logic_0_io_forwarding_idx)
      5'b00000:
        casez_tmp_176 = _GEN_985 & _GEN_99196;
      5'b00001:
        casez_tmp_176 = _GEN_991 & _GEN_99664;
      5'b00010:
        casez_tmp_176 = _GEN_997 & _GEN_100132;
      5'b00011:
        casez_tmp_176 = _GEN_1003 & _GEN_100600;
      5'b00100:
        casez_tmp_176 = _GEN_1009 & _GEN_101068;
      5'b00101:
        casez_tmp_176 = _GEN_1015 & _GEN_101536;
      5'b00110:
        casez_tmp_176 = _GEN_1021 & _GEN_102004;
      5'b00111:
        casez_tmp_176 = _GEN_1027 & _GEN_102472;
      5'b01000:
        casez_tmp_176 = _GEN_1033 & _GEN_102940;
      5'b01001:
        casez_tmp_176 = _GEN_1039 & _GEN_103408;
      5'b01010:
        casez_tmp_176 = _GEN_1045 & _GEN_103876;
      5'b01011:
        casez_tmp_176 = _GEN_1051 & _GEN_104344;
      5'b01100:
        casez_tmp_176 = _GEN_1057 & _GEN_104812;
      5'b01101:
        casez_tmp_176 = _GEN_1063 & _GEN_105280;
      5'b01110:
        casez_tmp_176 = _GEN_1069 & _GEN_105748;
      5'b01111:
        casez_tmp_176 = _GEN_1075 & _GEN_106216;
      5'b10000:
        casez_tmp_176 = _GEN_1081 & _GEN_106684;
      5'b10001:
        casez_tmp_176 = _GEN_1087 & _GEN_107152;
      5'b10010:
        casez_tmp_176 = _GEN_1093 & _GEN_107620;
      5'b10011:
        casez_tmp_176 = _GEN_1099 & _GEN_108088;
      5'b10100:
        casez_tmp_176 = _GEN_1105 & _GEN_108556;
      5'b10101:
        casez_tmp_176 = _GEN_1111 & _GEN_109024;
      5'b10110:
        casez_tmp_176 = _GEN_1117 & _GEN_109492;
      5'b10111:
        casez_tmp_176 = _GEN_1123 & _GEN_109960;
      5'b11000:
        casez_tmp_176 = _GEN_1129 & _GEN_110428;
      5'b11001:
        casez_tmp_176 = _GEN_1135 & _GEN_110896;
      5'b11010:
        casez_tmp_176 = _GEN_1141 & _GEN_111364;
      5'b11011:
        casez_tmp_176 = _GEN_1147 & _GEN_111832;
      5'b11100:
        casez_tmp_176 = _GEN_1153 & _GEN_112300;
      5'b11101:
        casez_tmp_176 = _GEN_1159 & _GEN_112768;
      5'b11110:
        casez_tmp_176 = _GEN_1165 & _GEN_113236;
      default:
        casez_tmp_176 = _GEN_1171 & _GEN_113704;
    endcase
  end // always @(*)
  reg         REG_2;
  always @(*) begin
    casez (_forwarding_age_logic_1_io_forwarding_idx)
      5'b00000:
        casez_tmp_177 = _GEN_988 & _GEN_99430;
      5'b00001:
        casez_tmp_177 = _GEN_994 & _GEN_99898;
      5'b00010:
        casez_tmp_177 = _GEN_1000 & _GEN_100366;
      5'b00011:
        casez_tmp_177 = _GEN_1006 & _GEN_100834;
      5'b00100:
        casez_tmp_177 = _GEN_1012 & _GEN_101302;
      5'b00101:
        casez_tmp_177 = _GEN_1018 & _GEN_101770;
      5'b00110:
        casez_tmp_177 = _GEN_1024 & _GEN_102238;
      5'b00111:
        casez_tmp_177 = _GEN_1030 & _GEN_102706;
      5'b01000:
        casez_tmp_177 = _GEN_1036 & _GEN_103174;
      5'b01001:
        casez_tmp_177 = _GEN_1042 & _GEN_103642;
      5'b01010:
        casez_tmp_177 = _GEN_1048 & _GEN_104110;
      5'b01011:
        casez_tmp_177 = _GEN_1054 & _GEN_104578;
      5'b01100:
        casez_tmp_177 = _GEN_1060 & _GEN_105046;
      5'b01101:
        casez_tmp_177 = _GEN_1066 & _GEN_105514;
      5'b01110:
        casez_tmp_177 = _GEN_1072 & _GEN_105982;
      5'b01111:
        casez_tmp_177 = _GEN_1078 & _GEN_106450;
      5'b10000:
        casez_tmp_177 = _GEN_1084 & _GEN_106918;
      5'b10001:
        casez_tmp_177 = _GEN_1090 & _GEN_107386;
      5'b10010:
        casez_tmp_177 = _GEN_1096 & _GEN_107854;
      5'b10011:
        casez_tmp_177 = _GEN_1102 & _GEN_108322;
      5'b10100:
        casez_tmp_177 = _GEN_1108 & _GEN_108790;
      5'b10101:
        casez_tmp_177 = _GEN_1114 & _GEN_109258;
      5'b10110:
        casez_tmp_177 = _GEN_1120 & _GEN_109726;
      5'b10111:
        casez_tmp_177 = _GEN_1126 & _GEN_110194;
      5'b11000:
        casez_tmp_177 = _GEN_1132 & _GEN_110662;
      5'b11001:
        casez_tmp_177 = _GEN_1138 & _GEN_111130;
      5'b11010:
        casez_tmp_177 = _GEN_1144 & _GEN_111598;
      5'b11011:
        casez_tmp_177 = _GEN_1150 & _GEN_112066;
      5'b11100:
        casez_tmp_177 = _GEN_1156 & _GEN_112534;
      5'b11101:
        casez_tmp_177 = _GEN_1162 & _GEN_113002;
      5'b11110:
        casez_tmp_177 = _GEN_1168 & _GEN_113470;
      default:
        casez_tmp_177 = _GEN_1174 & _GEN_113938;
    endcase
  end // always @(*)
  reg         REG_3;
  wire [5:0]  _l_idx_T_117 = failed_loads_9 & _temp_bits_T_18 ? 6'h9 : failed_loads_10 & _temp_bits_T_20 ? 6'hA : failed_loads_11 & _temp_bits_T_22 ? 6'hB : failed_loads_12 & _temp_bits_T_24 ? 6'hC : failed_loads_13 & _temp_bits_T_26 ? 6'hD : failed_loads_14 & _temp_bits_T_28 ? 6'hE : failed_loads_15 & ~(ldq_head[4]) ? 6'hF : failed_loads_16 & _temp_bits_T_32 ? 6'h10 : failed_loads_17 & _temp_bits_T_34 ? 6'h11 : failed_loads_18 & _temp_bits_T_36 ? 6'h12 : failed_loads_19 & _temp_bits_T_38 ? 6'h13 : failed_loads_20 & _temp_bits_T_40 ? 6'h14 : failed_loads_21 & _temp_bits_T_42 ? 6'h15 : failed_loads_22 & _temp_bits_T_44 ? 6'h16 : failed_loads_23 & _temp_bits_T_46 ? 6'h17 : failed_loads_24 & _temp_bits_T_48 ? 6'h18 : failed_loads_25 & _temp_bits_T_50 ? 6'h19 : failed_loads_26 & _temp_bits_T_52 ? 6'h1A : failed_loads_27 & _temp_bits_T_54 ? 6'h1B : failed_loads_28 & _temp_bits_T_56 ? 6'h1C : failed_loads_29 & _temp_bits_T_58 ? 6'h1D : failed_loads_30 & _temp_bits_T_60 ? 6'h1E : failed_loads_31 ? 6'h1F : failed_loads_0 ? 6'h20 : failed_loads_1 ? 6'h21 : failed_loads_2 ? 6'h22 : failed_loads_3 ? 6'h23 : failed_loads_4 ? 6'h24 : failed_loads_5 ? 6'h25 : failed_loads_6 ? 6'h26 : failed_loads_7 ? 6'h27 : failed_loads_8 ? 6'h28 : failed_loads_9 ? 6'h29 : failed_loads_10 ? 6'h2A : failed_loads_11 ? 6'h2B : failed_loads_12 ? 6'h2C : failed_loads_13 ? 6'h2D : failed_loads_14 ? 6'h2E : failed_loads_15 ? 6'h2F : failed_loads_16 ? 6'h30 : failed_loads_17 ? 6'h31 : failed_loads_18 ? 6'h32 : failed_loads_19 ? 6'h33 : failed_loads_20 ? 6'h34 : failed_loads_21 ? 6'h35 : failed_loads_22 ? 6'h36 : failed_loads_23 ? 6'h37 : failed_loads_24 ? 6'h38 : failed_loads_25 ? 6'h39 : failed_loads_26 ? 6'h3A : failed_loads_27 ? 6'h3B : failed_loads_28 ? 6'h3C : failed_loads_29 ? 6'h3D : {5'h1F, ~failed_loads_30};
  wire [4:0]  l_idx = failed_loads_0 & _temp_bits_T ? 5'h0 : failed_loads_1 & _temp_bits_T_2 ? 5'h1 : failed_loads_2 & _temp_bits_T_4 ? 5'h2 : failed_loads_3 & _temp_bits_T_6 ? 5'h3 : failed_loads_4 & _temp_bits_T_8 ? 5'h4 : failed_loads_5 & _temp_bits_T_10 ? 5'h5 : failed_loads_6 & _temp_bits_T_12 ? 5'h6 : failed_loads_7 & _temp_bits_T_14 ? 5'h7 : failed_loads_8 & _temp_bits_T_16 ? 5'h8 : _l_idx_T_117[4:0];
  reg         r_xcpt_valid;
  reg  [19:0] r_xcpt_uop_br_mask;
  reg  [6:0]  r_xcpt_uop_rob_idx;
  reg  [4:0]  r_xcpt_cause;
  reg  [39:0] r_xcpt_badvaddr;
  always @(*) begin
    casez (l_idx)
      5'b00000:
        casez_tmp_178 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_178 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_178 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_178 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_178 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_178 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_178 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_178 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_178 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_178 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_178 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_178 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_178 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_178 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_178 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_178 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_178 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_178 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_178 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_178 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_178 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_178 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_178 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_178 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_178 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_178 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_178 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_178 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_178 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_178 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_178 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_178 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (l_idx)
      5'b00000:
        casez_tmp_179 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_179 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_179 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_179 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_179 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_179 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_179 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_179 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_179 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_179 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_179 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_179 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_179 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_179 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_179 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_179 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_179 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_179 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_179 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_179 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_179 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_179 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_179 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_179 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_179 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_179 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_179 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_179 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_179 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_179 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_179 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_179 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  wire        _io_core_spec_ld_wakeup_0_valid_output = fired_load_incoming_0 & ~mem_incoming_uop_0_fp_val & (|mem_incoming_uop_0_pdst);
  wire        _io_core_spec_ld_wakeup_1_valid_output = fired_load_incoming_1 & ~mem_incoming_uop_1_fp_val & (|mem_incoming_uop_1_pdst);
  wire        _GEN_1177 = hella_state == 3'h6;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_180 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_180 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_180 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_180 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_180 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_180 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_180 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_180 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_180 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_180 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_180 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_180 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_180 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_180 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_180 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_180 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_180 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_180 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_180 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_180 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_180 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_180 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_180 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_180 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_180 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_180 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_180 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_180 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_180 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_180 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_180 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_180 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  wire        send_iresp = casez_tmp_180 == 2'h0;
  wire        send_fresp = casez_tmp_180 == 2'h1;
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_181 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_181 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_181 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_181 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_181 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_181 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_181 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_181 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_181 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_181 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_181 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_181 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_181 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_181 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_181 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_181 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_181 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_181 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_181 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_181 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_181 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_181 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_181 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_181 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_181 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_181 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_181 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_181 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_181 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_181 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_181 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_181 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_182 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_182 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_182 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_182 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_182 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_182 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_182 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_182 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_182 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_182 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_182 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_182 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_182 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_182 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_182 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_182 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_182 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_182 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_182 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_182 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_182 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_182 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_182 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_182 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_182 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_182 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_182 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_182 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_182 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_182 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_182 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_182 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_183 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_183 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_183 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_183 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_183 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_183 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_183 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_183 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_183 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_183 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_183 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_183 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_183 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_183 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_183 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_183 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_183 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_183 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_183 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_183 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_183 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_183 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_183 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_183 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_183 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_183 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_183 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_183 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_183 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_183 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_183 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_183 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_184 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_184 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_184 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_184 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_184 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_184 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_184 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_184 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_184 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_184 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_184 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_184 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_184 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_184 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_184 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_184 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_184 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_184 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_184 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_184 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_184 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_184 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_184 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_184 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_184 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_184 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_184 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_184 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_184 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_184 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_184 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_184 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_185 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_185 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_185 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_185 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_185 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_185 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_185 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_185 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_185 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_185 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_185 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_185 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_185 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_185 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_185 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_185 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_185 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_185 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_185 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_185 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_185 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_185 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_185 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_185 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_185 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_185 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_185 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_185 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_185 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_185 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_185 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_185 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_186 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_186 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_186 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_186 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_186 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_186 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_186 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_186 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_186 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_186 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_186 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_186 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_186 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_186 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_186 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_186 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_186 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_186 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_186 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_186 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_186 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_186 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_186 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_186 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_186 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_186 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_186 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_186 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_186 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_186 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_186 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_186 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_187 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_187 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_187 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_187 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_187 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_187 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_187 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_187 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_187 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_187 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_187 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_187 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_187 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_187 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_187 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_187 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_187 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_187 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_187 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_187 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_187 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_187 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_187 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_187 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_187 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_187 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_187 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_187 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_187 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_187 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_187 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_187 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_188 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_188 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_188 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_188 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_188 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_188 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_188 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_188 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_188 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_188 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_188 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_188 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_188 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_188 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_188 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_188 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_188 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_188 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_188 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_188 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_188 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_188 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_188 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_188 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_188 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_188 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_188 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_188 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_188 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_188 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_188 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_188 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_189 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_189 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_189 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_189 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_189 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_189 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_189 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_189 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_189 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_189 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_189 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_189 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_189 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_189 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_189 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_189 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_189 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_189 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_189 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_189 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_189 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_189 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_189 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_189 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_189 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_189 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_189 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_189 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_189 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_189 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_189 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_189 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_190 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_190 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_190 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_190 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_190 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_190 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_190 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_190 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_190 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_190 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_190 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_190 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_190 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_190 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_190 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_190 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_190 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_190 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_190 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_190 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_190 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_190 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_190 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_190 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_190 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_190 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_190 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_190 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_190 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_190 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_190 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_190 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_191 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_191 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_191 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_191 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_191 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_191 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_191 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_191 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_191 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_191 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_191 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_191 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_191 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_191 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_191 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_191 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_191 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_191 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_191 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_191 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_191 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_191 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_191 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_191 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_191 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_191 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_191 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_191 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_191 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_191 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_191 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_191 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_192 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_192 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_192 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_192 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_192 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_192 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_192 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_192 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_192 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_192 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_192 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_192 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_192 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_192 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_192 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_192 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_192 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_192 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_192 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_192 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_192 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_192 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_192 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_192 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_192 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_192 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_192 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_192 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_192 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_192 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_192 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_192 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_193 = stq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_193 = stq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_193 = stq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_193 = stq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_193 = stq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_193 = stq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_193 = stq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_193 = stq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_193 = stq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_193 = stq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_193 = stq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_193 = stq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_193 = stq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_193 = stq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_193 = stq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_193 = stq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_193 = stq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_193 = stq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_193 = stq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_193 = stq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_193 = stq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_193 = stq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_193 = stq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_193 = stq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_193 = stq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_193 = stq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_193 = stq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_193 = stq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_193 = stq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_193 = stq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_193 = stq_30_bits_uop_pdst;
      default:
        casez_tmp_193 = stq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_194 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_194 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_194 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_194 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_194 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_194 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_194 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_194 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_194 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_194 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_194 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_194 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_194 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_194 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_194 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_194 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_194 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_194 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_194 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_194 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_194 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_194 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_194 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_194 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_194 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_194 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_194 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_194 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_194 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_194 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_194 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_194 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_195 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_195 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_195 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_195 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_195 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_195 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_195 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_195 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_195 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_195 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_195 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_195 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_195 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_195 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_195 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_195 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_195 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_195 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_195 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_195 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_195 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_195 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_195 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_195 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_195 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_195 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_195 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_195 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_195 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_195 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_195 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_195 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_0_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_196 = stq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_196 = stq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_196 = stq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_196 = stq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_196 = stq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_196 = stq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_196 = stq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_196 = stq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_196 = stq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_196 = stq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_196 = stq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_196 = stq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_196 = stq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_196 = stq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_196 = stq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_196 = stq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_196 = stq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_196 = stq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_196 = stq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_196 = stq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_196 = stq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_196 = stq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_196 = stq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_196 = stq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_196 = stq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_196 = stq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_196 = stq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_196 = stq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_196 = stq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_196 = stq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_196 = stq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_196 = stq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  wire        _GEN_1178 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq;
  wire        dmem_resp_fired_0 = io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq | io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_is_amo);
  wire        _GEN_1179 = dmem_resp_fired_0 & wb_forward_valid_0;
  wire        _GEN_1180 = ~dmem_resp_fired_0 & wb_forward_valid_0;
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_197 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_197 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_197 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_197 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_197 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_197 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_197 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_197 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_197 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_197 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_197 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_197 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_197 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_197 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_197 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_197 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_197 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_197 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_197 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_197 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_197 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_197 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_197 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_197 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_197 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_197 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_197 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_197 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_197 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_197 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_197 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_197 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  wire        live = (io_core_brupdate_b1_mispredict_mask & casez_tmp_197) == 20'h0;
  always @(*) begin
    casez (wb_forward_stq_idx_0)
      5'b00000:
        casez_tmp_198 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_198 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_198 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_198 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_198 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_198 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_198 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_198 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_198 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_198 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_198 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_198 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_198 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_198 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_198 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_198 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_198 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_198 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_198 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_198 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_198 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_198 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_198 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_198 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_198 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_198 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_198 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_198 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_198 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_198 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_198 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_198 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_stq_idx_0)
      5'b00000:
        casez_tmp_199 = stq_0_bits_data_bits;
      5'b00001:
        casez_tmp_199 = stq_1_bits_data_bits;
      5'b00010:
        casez_tmp_199 = stq_2_bits_data_bits;
      5'b00011:
        casez_tmp_199 = stq_3_bits_data_bits;
      5'b00100:
        casez_tmp_199 = stq_4_bits_data_bits;
      5'b00101:
        casez_tmp_199 = stq_5_bits_data_bits;
      5'b00110:
        casez_tmp_199 = stq_6_bits_data_bits;
      5'b00111:
        casez_tmp_199 = stq_7_bits_data_bits;
      5'b01000:
        casez_tmp_199 = stq_8_bits_data_bits;
      5'b01001:
        casez_tmp_199 = stq_9_bits_data_bits;
      5'b01010:
        casez_tmp_199 = stq_10_bits_data_bits;
      5'b01011:
        casez_tmp_199 = stq_11_bits_data_bits;
      5'b01100:
        casez_tmp_199 = stq_12_bits_data_bits;
      5'b01101:
        casez_tmp_199 = stq_13_bits_data_bits;
      5'b01110:
        casez_tmp_199 = stq_14_bits_data_bits;
      5'b01111:
        casez_tmp_199 = stq_15_bits_data_bits;
      5'b10000:
        casez_tmp_199 = stq_16_bits_data_bits;
      5'b10001:
        casez_tmp_199 = stq_17_bits_data_bits;
      5'b10010:
        casez_tmp_199 = stq_18_bits_data_bits;
      5'b10011:
        casez_tmp_199 = stq_19_bits_data_bits;
      5'b10100:
        casez_tmp_199 = stq_20_bits_data_bits;
      5'b10101:
        casez_tmp_199 = stq_21_bits_data_bits;
      5'b10110:
        casez_tmp_199 = stq_22_bits_data_bits;
      5'b10111:
        casez_tmp_199 = stq_23_bits_data_bits;
      5'b11000:
        casez_tmp_199 = stq_24_bits_data_bits;
      5'b11001:
        casez_tmp_199 = stq_25_bits_data_bits;
      5'b11010:
        casez_tmp_199 = stq_26_bits_data_bits;
      5'b11011:
        casez_tmp_199 = stq_27_bits_data_bits;
      5'b11100:
        casez_tmp_199 = stq_28_bits_data_bits;
      5'b11101:
        casez_tmp_199 = stq_29_bits_data_bits;
      5'b11110:
        casez_tmp_199 = stq_30_bits_data_bits;
      default:
        casez_tmp_199 = stq_31_bits_data_bits;
    endcase
  end // always @(*)
  always @(*) begin
    casez (casez_tmp_198)
      2'b00:
        casez_tmp_200 = {2{{2{{2{casez_tmp_199[7:0]}}}}}};
      2'b01:
        casez_tmp_200 = {2{{2{casez_tmp_199[15:0]}}}};
      2'b10:
        casez_tmp_200 = {2{casez_tmp_199[31:0]}};
      default:
        casez_tmp_200 = casez_tmp_199;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_201 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_201 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_201 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_201 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_201 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_201 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_201 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_201 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_201 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_201 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_201 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_201 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_201 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_201 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_201 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_201 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_201 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_201 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_201 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_201 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_201 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_201 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_201 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_201 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_201 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_201 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_201 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_201 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_201 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_201 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_201 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_201 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_202 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_202 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_202 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_202 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_202 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_202 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_202 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_202 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_202 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_202 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_202 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_202 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_202 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_202 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_202 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_202 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_202 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_202 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_202 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_202 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_202 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_202 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_202 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_202 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_202 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_202 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_202 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_202 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_202 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_202 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_202 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_202 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_stq_idx_0)
      5'b00000:
        casez_tmp_203 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_203 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_203 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_203 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_203 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_203 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_203 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_203 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_203 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_203 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_203 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_203 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_203 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_203 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_203 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_203 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_203 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_203 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_203 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_203 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_203 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_203 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_203 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_203 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_203 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_203 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_203 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_203 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_203 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_203 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_203 = stq_30_bits_data_valid;
      default:
        casez_tmp_203 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_204 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_204 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_204 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_204 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_204 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_204 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_204 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_204 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_204 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_204 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_204 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_204 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_204 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_204 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_204 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_204 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_204 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_204 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_204 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_204 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_204 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_204 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_204 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_204 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_204 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_204 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_204 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_204 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_204 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_204 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_204 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_204 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_205 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_205 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_205 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_205 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_205 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_205 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_205 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_205 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_205 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_205 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_205 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_205 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_205 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_205 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_205 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_205 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_205 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_205 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_205 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_205 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_205 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_205 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_205 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_205 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_205 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_205 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_205 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_205 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_205 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_205 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_205 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_205 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_206 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_206 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_206 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_206 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_206 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_206 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_206 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_206 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_206 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_206 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_206 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_206 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_206 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_206 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_206 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_206 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_206 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_206 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_206 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_206 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_206 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_206 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_206 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_206 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_206 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_206 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_206 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_206 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_206 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_206 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_206 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_206 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_207 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_207 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_207 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_207 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_207 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_207 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_207 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_207 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_207 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_207 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_207 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_207 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_207 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_207 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_207 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_207 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_207 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_207 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_207 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_207 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_207 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_207 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_207 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_207 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_207 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_207 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_207 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_207 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_207 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_207 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_207 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_207 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_208 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_208 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_208 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_208 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_208 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_208 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_208 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_208 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_208 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_208 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_208 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_208 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_208 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_208 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_208 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_208 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_208 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_208 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_208 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_208 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_208 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_208 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_208 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_208 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_208 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_208 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_208 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_208 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_208 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_208 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_208 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_208 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_209 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_209 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_209 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_209 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_209 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_209 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_209 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_209 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_209 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_209 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_209 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_209 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_209 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_209 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_209 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_209 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_209 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_209 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_209 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_209 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_209 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_209 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_209 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_209 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_209 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_209 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_209 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_209 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_209 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_209 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_209 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_209 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_210 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_210 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_210 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_210 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_210 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_210 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_210 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_210 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_210 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_210 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_210 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_210 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_210 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_210 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_210 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_210 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_210 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_210 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_210 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_210 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_210 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_210 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_210 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_210 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_210 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_210 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_210 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_210 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_210 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_210 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_210 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_210 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_211 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_211 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_211 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_211 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_211 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_211 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_211 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_211 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_211 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_211 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_211 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_211 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_211 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_211 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_211 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_211 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_211 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_211 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_211 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_211 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_211 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_211 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_211 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_211 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_211 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_211 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_211 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_211 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_211 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_211 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_211 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_211 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_0)
      5'b00000:
        casez_tmp_212 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_212 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_212 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_212 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_212 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_212 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_212 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_212 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_212 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_212 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_212 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_212 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_212 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_212 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_212 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_212 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_212 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_212 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_212 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_212 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_212 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_212 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_212 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_212 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_212 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_212 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_212 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_212 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_212 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_212 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_212 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_212 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  wire [31:0] io_core_exe_0_iresp_bits_data_zeroed = wb_forward_ld_addr_0[2] ? casez_tmp_200[63:32] : casez_tmp_200[31:0];
  wire        _ldq_bits_debug_wb_data_T_1 = casez_tmp_201 == 2'h2;
  wire [15:0] io_core_exe_0_iresp_bits_data_zeroed_1 = wb_forward_ld_addr_0[1] ? io_core_exe_0_iresp_bits_data_zeroed[31:16] : io_core_exe_0_iresp_bits_data_zeroed[15:0];
  wire        _ldq_bits_debug_wb_data_T_10 = casez_tmp_201 == 2'h1;
  wire [7:0]  io_core_exe_0_iresp_bits_data_zeroed_2 = wb_forward_ld_addr_0[0] ? io_core_exe_0_iresp_bits_data_zeroed_1[15:8] : io_core_exe_0_iresp_bits_data_zeroed_1[7:0];
  wire        _ldq_bits_debug_wb_data_T_19 = casez_tmp_201 == 2'h0;
  wire [31:0] io_core_exe_0_fresp_bits_data_zeroed = wb_forward_ld_addr_0[2] ? casez_tmp_200[63:32] : casez_tmp_200[31:0];
  wire [15:0] io_core_exe_0_fresp_bits_data_zeroed_1 = wb_forward_ld_addr_0[1] ? io_core_exe_0_fresp_bits_data_zeroed[31:16] : io_core_exe_0_fresp_bits_data_zeroed[15:0];
  wire [7:0]  io_core_exe_0_fresp_bits_data_zeroed_2 = wb_forward_ld_addr_0[0] ? io_core_exe_0_fresp_bits_data_zeroed_1[15:8] : io_core_exe_0_fresp_bits_data_zeroed_1[7:0];
  wire        _GEN_1181 = _GEN_1179 | ~_GEN_1180;
  wire        _io_core_exe_0_iresp_valid_output = _GEN_1181 ? io_dmem_resp_0_valid & (io_dmem_resp_0_bits_uop_uses_ldq ? send_iresp : io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_is_amo) : casez_tmp_202 == 2'h0 & casez_tmp_203 & live;
  wire        _io_core_exe_0_fresp_valid_output = _GEN_1181 ? _GEN_1178 & send_fresp : casez_tmp_202 == 2'h1 & casez_tmp_203 & live;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_213 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_213 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_213 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_213 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_213 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_213 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_213 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_213 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_213 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_213 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_213 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_213 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_213 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_213 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_213 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_213 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_213 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_213 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_213 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_213 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_213 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_213 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_213 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_213 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_213 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_213 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_213 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_213 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_213 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_213 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_213 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_213 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  wire        send_iresp_1 = casez_tmp_213 == 2'h0;
  wire        send_fresp_1 = casez_tmp_213 == 2'h1;
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_214 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_214 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_214 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_214 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_214 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_214 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_214 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_214 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_214 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_214 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_214 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_214 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_214 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_214 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_214 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_214 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_214 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_214 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_214 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_214 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_214 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_214 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_214 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_214 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_214 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_214 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_214 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_214 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_214 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_214 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_214 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_214 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_215 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_215 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_215 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_215 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_215 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_215 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_215 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_215 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_215 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_215 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_215 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_215 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_215 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_215 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_215 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_215 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_215 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_215 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_215 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_215 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_215 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_215 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_215 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_215 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_215 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_215 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_215 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_215 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_215 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_215 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_215 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_215 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_216 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_216 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_216 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_216 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_216 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_216 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_216 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_216 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_216 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_216 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_216 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_216 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_216 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_216 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_216 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_216 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_216 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_216 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_216 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_216 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_216 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_216 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_216 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_216 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_216 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_216 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_216 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_216 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_216 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_216 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_216 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_216 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_217 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_217 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_217 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_217 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_217 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_217 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_217 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_217 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_217 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_217 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_217 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_217 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_217 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_217 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_217 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_217 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_217 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_217 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_217 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_217 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_217 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_217 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_217 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_217 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_217 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_217 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_217 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_217 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_217 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_217 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_217 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_217 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_218 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_218 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_218 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_218 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_218 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_218 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_218 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_218 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_218 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_218 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_218 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_218 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_218 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_218 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_218 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_218 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_218 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_218 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_218 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_218 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_218 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_218 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_218 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_218 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_218 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_218 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_218 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_218 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_218 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_218 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_218 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_218 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_219 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_219 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_219 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_219 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_219 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_219 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_219 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_219 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_219 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_219 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_219 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_219 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_219 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_219 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_219 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_219 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_219 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_219 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_219 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_219 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_219 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_219 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_219 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_219 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_219 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_219 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_219 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_219 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_219 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_219 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_219 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_219 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_220 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_220 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_220 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_220 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_220 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_220 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_220 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_220 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_220 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_220 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_220 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_220 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_220 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_220 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_220 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_220 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_220 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_220 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_220 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_220 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_220 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_220 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_220 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_220 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_220 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_220 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_220 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_220 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_220 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_220 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_220 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_220 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_221 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_221 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_221 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_221 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_221 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_221 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_221 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_221 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_221 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_221 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_221 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_221 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_221 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_221 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_221 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_221 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_221 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_221 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_221 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_221 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_221 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_221 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_221 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_221 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_221 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_221 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_221 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_221 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_221 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_221 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_221 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_221 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_222 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_222 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_222 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_222 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_222 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_222 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_222 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_222 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_222 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_222 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_222 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_222 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_222 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_222 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_222 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_222 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_222 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_222 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_222 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_222 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_222 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_222 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_222 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_222 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_222 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_222 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_222 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_222 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_222 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_222 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_222 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_222 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_ldq_idx)
      5'b00000:
        casez_tmp_223 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_223 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_223 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_223 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_223 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_223 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_223 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_223 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_223 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_223 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_223 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_223 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_223 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_223 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_223 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_223 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_223 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_223 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_223 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_223 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_223 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_223 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_223 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_223 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_223 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_223 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_223 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_223 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_223 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_223 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_223 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_223 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_224 = stq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_224 = stq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_224 = stq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_224 = stq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_224 = stq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_224 = stq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_224 = stq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_224 = stq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_224 = stq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_224 = stq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_224 = stq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_224 = stq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_224 = stq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_224 = stq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_224 = stq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_224 = stq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_224 = stq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_224 = stq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_224 = stq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_224 = stq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_224 = stq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_224 = stq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_224 = stq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_224 = stq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_224 = stq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_224 = stq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_224 = stq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_224 = stq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_224 = stq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_224 = stq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_224 = stq_30_bits_uop_rob_idx;
      default:
        casez_tmp_224 = stq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_225 = stq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_225 = stq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_225 = stq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_225 = stq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_225 = stq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_225 = stq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_225 = stq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_225 = stq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_225 = stq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_225 = stq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_225 = stq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_225 = stq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_225 = stq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_225 = stq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_225 = stq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_225 = stq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_225 = stq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_225 = stq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_225 = stq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_225 = stq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_225 = stq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_225 = stq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_225 = stq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_225 = stq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_225 = stq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_225 = stq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_225 = stq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_225 = stq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_225 = stq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_225 = stq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_225 = stq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_225 = stq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_226 = stq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_226 = stq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_226 = stq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_226 = stq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_226 = stq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_226 = stq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_226 = stq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_226 = stq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_226 = stq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_226 = stq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_226 = stq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_226 = stq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_226 = stq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_226 = stq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_226 = stq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_226 = stq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_226 = stq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_226 = stq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_226 = stq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_226 = stq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_226 = stq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_226 = stq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_226 = stq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_226 = stq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_226 = stq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_226 = stq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_226 = stq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_226 = stq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_226 = stq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_226 = stq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_226 = stq_30_bits_uop_pdst;
      default:
        casez_tmp_226 = stq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_227 = stq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_227 = stq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_227 = stq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_227 = stq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_227 = stq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_227 = stq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_227 = stq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_227 = stq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_227 = stq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_227 = stq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_227 = stq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_227 = stq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_227 = stq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_227 = stq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_227 = stq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_227 = stq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_227 = stq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_227 = stq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_227 = stq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_227 = stq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_227 = stq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_227 = stq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_227 = stq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_227 = stq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_227 = stq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_227 = stq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_227 = stq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_227 = stq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_227 = stq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_227 = stq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_227 = stq_30_bits_uop_is_amo;
      default:
        casez_tmp_227 = stq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_228 = stq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_228 = stq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_228 = stq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_228 = stq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_228 = stq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_228 = stq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_228 = stq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_228 = stq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_228 = stq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_228 = stq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_228 = stq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_228 = stq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_228 = stq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_228 = stq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_228 = stq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_228 = stq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_228 = stq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_228 = stq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_228 = stq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_228 = stq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_228 = stq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_228 = stq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_228 = stq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_228 = stq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_228 = stq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_228 = stq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_228 = stq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_228 = stq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_228 = stq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_228 = stq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_228 = stq_30_bits_uop_uses_stq;
      default:
        casez_tmp_228 = stq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (io_dmem_resp_1_bits_uop_stq_idx)
      5'b00000:
        casez_tmp_229 = stq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_229 = stq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_229 = stq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_229 = stq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_229 = stq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_229 = stq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_229 = stq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_229 = stq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_229 = stq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_229 = stq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_229 = stq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_229 = stq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_229 = stq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_229 = stq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_229 = stq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_229 = stq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_229 = stq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_229 = stq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_229 = stq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_229 = stq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_229 = stq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_229 = stq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_229 = stq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_229 = stq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_229 = stq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_229 = stq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_229 = stq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_229 = stq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_229 = stq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_229 = stq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_229 = stq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_229 = stq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  wire        _GEN_1182 = io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq;
  wire        dmem_resp_fired_1 = io_dmem_resp_1_valid & (io_dmem_resp_1_bits_uop_uses_ldq | io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_is_amo);
  wire        _GEN_1183 = dmem_resp_fired_1 & wb_forward_valid_1;
  wire        _GEN_1184 = ~dmem_resp_fired_1 & wb_forward_valid_1;
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_230 = ldq_0_bits_uop_br_mask;
      5'b00001:
        casez_tmp_230 = ldq_1_bits_uop_br_mask;
      5'b00010:
        casez_tmp_230 = ldq_2_bits_uop_br_mask;
      5'b00011:
        casez_tmp_230 = ldq_3_bits_uop_br_mask;
      5'b00100:
        casez_tmp_230 = ldq_4_bits_uop_br_mask;
      5'b00101:
        casez_tmp_230 = ldq_5_bits_uop_br_mask;
      5'b00110:
        casez_tmp_230 = ldq_6_bits_uop_br_mask;
      5'b00111:
        casez_tmp_230 = ldq_7_bits_uop_br_mask;
      5'b01000:
        casez_tmp_230 = ldq_8_bits_uop_br_mask;
      5'b01001:
        casez_tmp_230 = ldq_9_bits_uop_br_mask;
      5'b01010:
        casez_tmp_230 = ldq_10_bits_uop_br_mask;
      5'b01011:
        casez_tmp_230 = ldq_11_bits_uop_br_mask;
      5'b01100:
        casez_tmp_230 = ldq_12_bits_uop_br_mask;
      5'b01101:
        casez_tmp_230 = ldq_13_bits_uop_br_mask;
      5'b01110:
        casez_tmp_230 = ldq_14_bits_uop_br_mask;
      5'b01111:
        casez_tmp_230 = ldq_15_bits_uop_br_mask;
      5'b10000:
        casez_tmp_230 = ldq_16_bits_uop_br_mask;
      5'b10001:
        casez_tmp_230 = ldq_17_bits_uop_br_mask;
      5'b10010:
        casez_tmp_230 = ldq_18_bits_uop_br_mask;
      5'b10011:
        casez_tmp_230 = ldq_19_bits_uop_br_mask;
      5'b10100:
        casez_tmp_230 = ldq_20_bits_uop_br_mask;
      5'b10101:
        casez_tmp_230 = ldq_21_bits_uop_br_mask;
      5'b10110:
        casez_tmp_230 = ldq_22_bits_uop_br_mask;
      5'b10111:
        casez_tmp_230 = ldq_23_bits_uop_br_mask;
      5'b11000:
        casez_tmp_230 = ldq_24_bits_uop_br_mask;
      5'b11001:
        casez_tmp_230 = ldq_25_bits_uop_br_mask;
      5'b11010:
        casez_tmp_230 = ldq_26_bits_uop_br_mask;
      5'b11011:
        casez_tmp_230 = ldq_27_bits_uop_br_mask;
      5'b11100:
        casez_tmp_230 = ldq_28_bits_uop_br_mask;
      5'b11101:
        casez_tmp_230 = ldq_29_bits_uop_br_mask;
      5'b11110:
        casez_tmp_230 = ldq_30_bits_uop_br_mask;
      default:
        casez_tmp_230 = ldq_31_bits_uop_br_mask;
    endcase
  end // always @(*)
  wire        live_1 = (io_core_brupdate_b1_mispredict_mask & casez_tmp_230) == 20'h0;
  always @(*) begin
    casez (wb_forward_stq_idx_1)
      5'b00000:
        casez_tmp_231 = stq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_231 = stq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_231 = stq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_231 = stq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_231 = stq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_231 = stq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_231 = stq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_231 = stq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_231 = stq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_231 = stq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_231 = stq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_231 = stq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_231 = stq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_231 = stq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_231 = stq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_231 = stq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_231 = stq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_231 = stq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_231 = stq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_231 = stq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_231 = stq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_231 = stq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_231 = stq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_231 = stq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_231 = stq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_231 = stq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_231 = stq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_231 = stq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_231 = stq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_231 = stq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_231 = stq_30_bits_uop_mem_size;
      default:
        casez_tmp_231 = stq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_stq_idx_1)
      5'b00000:
        casez_tmp_232 = stq_0_bits_data_bits;
      5'b00001:
        casez_tmp_232 = stq_1_bits_data_bits;
      5'b00010:
        casez_tmp_232 = stq_2_bits_data_bits;
      5'b00011:
        casez_tmp_232 = stq_3_bits_data_bits;
      5'b00100:
        casez_tmp_232 = stq_4_bits_data_bits;
      5'b00101:
        casez_tmp_232 = stq_5_bits_data_bits;
      5'b00110:
        casez_tmp_232 = stq_6_bits_data_bits;
      5'b00111:
        casez_tmp_232 = stq_7_bits_data_bits;
      5'b01000:
        casez_tmp_232 = stq_8_bits_data_bits;
      5'b01001:
        casez_tmp_232 = stq_9_bits_data_bits;
      5'b01010:
        casez_tmp_232 = stq_10_bits_data_bits;
      5'b01011:
        casez_tmp_232 = stq_11_bits_data_bits;
      5'b01100:
        casez_tmp_232 = stq_12_bits_data_bits;
      5'b01101:
        casez_tmp_232 = stq_13_bits_data_bits;
      5'b01110:
        casez_tmp_232 = stq_14_bits_data_bits;
      5'b01111:
        casez_tmp_232 = stq_15_bits_data_bits;
      5'b10000:
        casez_tmp_232 = stq_16_bits_data_bits;
      5'b10001:
        casez_tmp_232 = stq_17_bits_data_bits;
      5'b10010:
        casez_tmp_232 = stq_18_bits_data_bits;
      5'b10011:
        casez_tmp_232 = stq_19_bits_data_bits;
      5'b10100:
        casez_tmp_232 = stq_20_bits_data_bits;
      5'b10101:
        casez_tmp_232 = stq_21_bits_data_bits;
      5'b10110:
        casez_tmp_232 = stq_22_bits_data_bits;
      5'b10111:
        casez_tmp_232 = stq_23_bits_data_bits;
      5'b11000:
        casez_tmp_232 = stq_24_bits_data_bits;
      5'b11001:
        casez_tmp_232 = stq_25_bits_data_bits;
      5'b11010:
        casez_tmp_232 = stq_26_bits_data_bits;
      5'b11011:
        casez_tmp_232 = stq_27_bits_data_bits;
      5'b11100:
        casez_tmp_232 = stq_28_bits_data_bits;
      5'b11101:
        casez_tmp_232 = stq_29_bits_data_bits;
      5'b11110:
        casez_tmp_232 = stq_30_bits_data_bits;
      default:
        casez_tmp_232 = stq_31_bits_data_bits;
    endcase
  end // always @(*)
  always @(*) begin
    casez (casez_tmp_231)
      2'b00:
        casez_tmp_233 = {2{{2{{2{casez_tmp_232[7:0]}}}}}};
      2'b01:
        casez_tmp_233 = {2{{2{casez_tmp_232[15:0]}}}};
      2'b10:
        casez_tmp_233 = {2{casez_tmp_232[31:0]}};
      default:
        casez_tmp_233 = casez_tmp_232;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_234 = ldq_0_bits_uop_mem_size;
      5'b00001:
        casez_tmp_234 = ldq_1_bits_uop_mem_size;
      5'b00010:
        casez_tmp_234 = ldq_2_bits_uop_mem_size;
      5'b00011:
        casez_tmp_234 = ldq_3_bits_uop_mem_size;
      5'b00100:
        casez_tmp_234 = ldq_4_bits_uop_mem_size;
      5'b00101:
        casez_tmp_234 = ldq_5_bits_uop_mem_size;
      5'b00110:
        casez_tmp_234 = ldq_6_bits_uop_mem_size;
      5'b00111:
        casez_tmp_234 = ldq_7_bits_uop_mem_size;
      5'b01000:
        casez_tmp_234 = ldq_8_bits_uop_mem_size;
      5'b01001:
        casez_tmp_234 = ldq_9_bits_uop_mem_size;
      5'b01010:
        casez_tmp_234 = ldq_10_bits_uop_mem_size;
      5'b01011:
        casez_tmp_234 = ldq_11_bits_uop_mem_size;
      5'b01100:
        casez_tmp_234 = ldq_12_bits_uop_mem_size;
      5'b01101:
        casez_tmp_234 = ldq_13_bits_uop_mem_size;
      5'b01110:
        casez_tmp_234 = ldq_14_bits_uop_mem_size;
      5'b01111:
        casez_tmp_234 = ldq_15_bits_uop_mem_size;
      5'b10000:
        casez_tmp_234 = ldq_16_bits_uop_mem_size;
      5'b10001:
        casez_tmp_234 = ldq_17_bits_uop_mem_size;
      5'b10010:
        casez_tmp_234 = ldq_18_bits_uop_mem_size;
      5'b10011:
        casez_tmp_234 = ldq_19_bits_uop_mem_size;
      5'b10100:
        casez_tmp_234 = ldq_20_bits_uop_mem_size;
      5'b10101:
        casez_tmp_234 = ldq_21_bits_uop_mem_size;
      5'b10110:
        casez_tmp_234 = ldq_22_bits_uop_mem_size;
      5'b10111:
        casez_tmp_234 = ldq_23_bits_uop_mem_size;
      5'b11000:
        casez_tmp_234 = ldq_24_bits_uop_mem_size;
      5'b11001:
        casez_tmp_234 = ldq_25_bits_uop_mem_size;
      5'b11010:
        casez_tmp_234 = ldq_26_bits_uop_mem_size;
      5'b11011:
        casez_tmp_234 = ldq_27_bits_uop_mem_size;
      5'b11100:
        casez_tmp_234 = ldq_28_bits_uop_mem_size;
      5'b11101:
        casez_tmp_234 = ldq_29_bits_uop_mem_size;
      5'b11110:
        casez_tmp_234 = ldq_30_bits_uop_mem_size;
      default:
        casez_tmp_234 = ldq_31_bits_uop_mem_size;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_235 = ldq_0_bits_uop_dst_rtype;
      5'b00001:
        casez_tmp_235 = ldq_1_bits_uop_dst_rtype;
      5'b00010:
        casez_tmp_235 = ldq_2_bits_uop_dst_rtype;
      5'b00011:
        casez_tmp_235 = ldq_3_bits_uop_dst_rtype;
      5'b00100:
        casez_tmp_235 = ldq_4_bits_uop_dst_rtype;
      5'b00101:
        casez_tmp_235 = ldq_5_bits_uop_dst_rtype;
      5'b00110:
        casez_tmp_235 = ldq_6_bits_uop_dst_rtype;
      5'b00111:
        casez_tmp_235 = ldq_7_bits_uop_dst_rtype;
      5'b01000:
        casez_tmp_235 = ldq_8_bits_uop_dst_rtype;
      5'b01001:
        casez_tmp_235 = ldq_9_bits_uop_dst_rtype;
      5'b01010:
        casez_tmp_235 = ldq_10_bits_uop_dst_rtype;
      5'b01011:
        casez_tmp_235 = ldq_11_bits_uop_dst_rtype;
      5'b01100:
        casez_tmp_235 = ldq_12_bits_uop_dst_rtype;
      5'b01101:
        casez_tmp_235 = ldq_13_bits_uop_dst_rtype;
      5'b01110:
        casez_tmp_235 = ldq_14_bits_uop_dst_rtype;
      5'b01111:
        casez_tmp_235 = ldq_15_bits_uop_dst_rtype;
      5'b10000:
        casez_tmp_235 = ldq_16_bits_uop_dst_rtype;
      5'b10001:
        casez_tmp_235 = ldq_17_bits_uop_dst_rtype;
      5'b10010:
        casez_tmp_235 = ldq_18_bits_uop_dst_rtype;
      5'b10011:
        casez_tmp_235 = ldq_19_bits_uop_dst_rtype;
      5'b10100:
        casez_tmp_235 = ldq_20_bits_uop_dst_rtype;
      5'b10101:
        casez_tmp_235 = ldq_21_bits_uop_dst_rtype;
      5'b10110:
        casez_tmp_235 = ldq_22_bits_uop_dst_rtype;
      5'b10111:
        casez_tmp_235 = ldq_23_bits_uop_dst_rtype;
      5'b11000:
        casez_tmp_235 = ldq_24_bits_uop_dst_rtype;
      5'b11001:
        casez_tmp_235 = ldq_25_bits_uop_dst_rtype;
      5'b11010:
        casez_tmp_235 = ldq_26_bits_uop_dst_rtype;
      5'b11011:
        casez_tmp_235 = ldq_27_bits_uop_dst_rtype;
      5'b11100:
        casez_tmp_235 = ldq_28_bits_uop_dst_rtype;
      5'b11101:
        casez_tmp_235 = ldq_29_bits_uop_dst_rtype;
      5'b11110:
        casez_tmp_235 = ldq_30_bits_uop_dst_rtype;
      default:
        casez_tmp_235 = ldq_31_bits_uop_dst_rtype;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_stq_idx_1)
      5'b00000:
        casez_tmp_236 = stq_0_bits_data_valid;
      5'b00001:
        casez_tmp_236 = stq_1_bits_data_valid;
      5'b00010:
        casez_tmp_236 = stq_2_bits_data_valid;
      5'b00011:
        casez_tmp_236 = stq_3_bits_data_valid;
      5'b00100:
        casez_tmp_236 = stq_4_bits_data_valid;
      5'b00101:
        casez_tmp_236 = stq_5_bits_data_valid;
      5'b00110:
        casez_tmp_236 = stq_6_bits_data_valid;
      5'b00111:
        casez_tmp_236 = stq_7_bits_data_valid;
      5'b01000:
        casez_tmp_236 = stq_8_bits_data_valid;
      5'b01001:
        casez_tmp_236 = stq_9_bits_data_valid;
      5'b01010:
        casez_tmp_236 = stq_10_bits_data_valid;
      5'b01011:
        casez_tmp_236 = stq_11_bits_data_valid;
      5'b01100:
        casez_tmp_236 = stq_12_bits_data_valid;
      5'b01101:
        casez_tmp_236 = stq_13_bits_data_valid;
      5'b01110:
        casez_tmp_236 = stq_14_bits_data_valid;
      5'b01111:
        casez_tmp_236 = stq_15_bits_data_valid;
      5'b10000:
        casez_tmp_236 = stq_16_bits_data_valid;
      5'b10001:
        casez_tmp_236 = stq_17_bits_data_valid;
      5'b10010:
        casez_tmp_236 = stq_18_bits_data_valid;
      5'b10011:
        casez_tmp_236 = stq_19_bits_data_valid;
      5'b10100:
        casez_tmp_236 = stq_20_bits_data_valid;
      5'b10101:
        casez_tmp_236 = stq_21_bits_data_valid;
      5'b10110:
        casez_tmp_236 = stq_22_bits_data_valid;
      5'b10111:
        casez_tmp_236 = stq_23_bits_data_valid;
      5'b11000:
        casez_tmp_236 = stq_24_bits_data_valid;
      5'b11001:
        casez_tmp_236 = stq_25_bits_data_valid;
      5'b11010:
        casez_tmp_236 = stq_26_bits_data_valid;
      5'b11011:
        casez_tmp_236 = stq_27_bits_data_valid;
      5'b11100:
        casez_tmp_236 = stq_28_bits_data_valid;
      5'b11101:
        casez_tmp_236 = stq_29_bits_data_valid;
      5'b11110:
        casez_tmp_236 = stq_30_bits_data_valid;
      default:
        casez_tmp_236 = stq_31_bits_data_valid;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_237 = ldq_0_bits_uop_uopc;
      5'b00001:
        casez_tmp_237 = ldq_1_bits_uop_uopc;
      5'b00010:
        casez_tmp_237 = ldq_2_bits_uop_uopc;
      5'b00011:
        casez_tmp_237 = ldq_3_bits_uop_uopc;
      5'b00100:
        casez_tmp_237 = ldq_4_bits_uop_uopc;
      5'b00101:
        casez_tmp_237 = ldq_5_bits_uop_uopc;
      5'b00110:
        casez_tmp_237 = ldq_6_bits_uop_uopc;
      5'b00111:
        casez_tmp_237 = ldq_7_bits_uop_uopc;
      5'b01000:
        casez_tmp_237 = ldq_8_bits_uop_uopc;
      5'b01001:
        casez_tmp_237 = ldq_9_bits_uop_uopc;
      5'b01010:
        casez_tmp_237 = ldq_10_bits_uop_uopc;
      5'b01011:
        casez_tmp_237 = ldq_11_bits_uop_uopc;
      5'b01100:
        casez_tmp_237 = ldq_12_bits_uop_uopc;
      5'b01101:
        casez_tmp_237 = ldq_13_bits_uop_uopc;
      5'b01110:
        casez_tmp_237 = ldq_14_bits_uop_uopc;
      5'b01111:
        casez_tmp_237 = ldq_15_bits_uop_uopc;
      5'b10000:
        casez_tmp_237 = ldq_16_bits_uop_uopc;
      5'b10001:
        casez_tmp_237 = ldq_17_bits_uop_uopc;
      5'b10010:
        casez_tmp_237 = ldq_18_bits_uop_uopc;
      5'b10011:
        casez_tmp_237 = ldq_19_bits_uop_uopc;
      5'b10100:
        casez_tmp_237 = ldq_20_bits_uop_uopc;
      5'b10101:
        casez_tmp_237 = ldq_21_bits_uop_uopc;
      5'b10110:
        casez_tmp_237 = ldq_22_bits_uop_uopc;
      5'b10111:
        casez_tmp_237 = ldq_23_bits_uop_uopc;
      5'b11000:
        casez_tmp_237 = ldq_24_bits_uop_uopc;
      5'b11001:
        casez_tmp_237 = ldq_25_bits_uop_uopc;
      5'b11010:
        casez_tmp_237 = ldq_26_bits_uop_uopc;
      5'b11011:
        casez_tmp_237 = ldq_27_bits_uop_uopc;
      5'b11100:
        casez_tmp_237 = ldq_28_bits_uop_uopc;
      5'b11101:
        casez_tmp_237 = ldq_29_bits_uop_uopc;
      5'b11110:
        casez_tmp_237 = ldq_30_bits_uop_uopc;
      default:
        casez_tmp_237 = ldq_31_bits_uop_uopc;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_238 = ldq_0_bits_uop_rob_idx;
      5'b00001:
        casez_tmp_238 = ldq_1_bits_uop_rob_idx;
      5'b00010:
        casez_tmp_238 = ldq_2_bits_uop_rob_idx;
      5'b00011:
        casez_tmp_238 = ldq_3_bits_uop_rob_idx;
      5'b00100:
        casez_tmp_238 = ldq_4_bits_uop_rob_idx;
      5'b00101:
        casez_tmp_238 = ldq_5_bits_uop_rob_idx;
      5'b00110:
        casez_tmp_238 = ldq_6_bits_uop_rob_idx;
      5'b00111:
        casez_tmp_238 = ldq_7_bits_uop_rob_idx;
      5'b01000:
        casez_tmp_238 = ldq_8_bits_uop_rob_idx;
      5'b01001:
        casez_tmp_238 = ldq_9_bits_uop_rob_idx;
      5'b01010:
        casez_tmp_238 = ldq_10_bits_uop_rob_idx;
      5'b01011:
        casez_tmp_238 = ldq_11_bits_uop_rob_idx;
      5'b01100:
        casez_tmp_238 = ldq_12_bits_uop_rob_idx;
      5'b01101:
        casez_tmp_238 = ldq_13_bits_uop_rob_idx;
      5'b01110:
        casez_tmp_238 = ldq_14_bits_uop_rob_idx;
      5'b01111:
        casez_tmp_238 = ldq_15_bits_uop_rob_idx;
      5'b10000:
        casez_tmp_238 = ldq_16_bits_uop_rob_idx;
      5'b10001:
        casez_tmp_238 = ldq_17_bits_uop_rob_idx;
      5'b10010:
        casez_tmp_238 = ldq_18_bits_uop_rob_idx;
      5'b10011:
        casez_tmp_238 = ldq_19_bits_uop_rob_idx;
      5'b10100:
        casez_tmp_238 = ldq_20_bits_uop_rob_idx;
      5'b10101:
        casez_tmp_238 = ldq_21_bits_uop_rob_idx;
      5'b10110:
        casez_tmp_238 = ldq_22_bits_uop_rob_idx;
      5'b10111:
        casez_tmp_238 = ldq_23_bits_uop_rob_idx;
      5'b11000:
        casez_tmp_238 = ldq_24_bits_uop_rob_idx;
      5'b11001:
        casez_tmp_238 = ldq_25_bits_uop_rob_idx;
      5'b11010:
        casez_tmp_238 = ldq_26_bits_uop_rob_idx;
      5'b11011:
        casez_tmp_238 = ldq_27_bits_uop_rob_idx;
      5'b11100:
        casez_tmp_238 = ldq_28_bits_uop_rob_idx;
      5'b11101:
        casez_tmp_238 = ldq_29_bits_uop_rob_idx;
      5'b11110:
        casez_tmp_238 = ldq_30_bits_uop_rob_idx;
      default:
        casez_tmp_238 = ldq_31_bits_uop_rob_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_239 = ldq_0_bits_uop_ldq_idx;
      5'b00001:
        casez_tmp_239 = ldq_1_bits_uop_ldq_idx;
      5'b00010:
        casez_tmp_239 = ldq_2_bits_uop_ldq_idx;
      5'b00011:
        casez_tmp_239 = ldq_3_bits_uop_ldq_idx;
      5'b00100:
        casez_tmp_239 = ldq_4_bits_uop_ldq_idx;
      5'b00101:
        casez_tmp_239 = ldq_5_bits_uop_ldq_idx;
      5'b00110:
        casez_tmp_239 = ldq_6_bits_uop_ldq_idx;
      5'b00111:
        casez_tmp_239 = ldq_7_bits_uop_ldq_idx;
      5'b01000:
        casez_tmp_239 = ldq_8_bits_uop_ldq_idx;
      5'b01001:
        casez_tmp_239 = ldq_9_bits_uop_ldq_idx;
      5'b01010:
        casez_tmp_239 = ldq_10_bits_uop_ldq_idx;
      5'b01011:
        casez_tmp_239 = ldq_11_bits_uop_ldq_idx;
      5'b01100:
        casez_tmp_239 = ldq_12_bits_uop_ldq_idx;
      5'b01101:
        casez_tmp_239 = ldq_13_bits_uop_ldq_idx;
      5'b01110:
        casez_tmp_239 = ldq_14_bits_uop_ldq_idx;
      5'b01111:
        casez_tmp_239 = ldq_15_bits_uop_ldq_idx;
      5'b10000:
        casez_tmp_239 = ldq_16_bits_uop_ldq_idx;
      5'b10001:
        casez_tmp_239 = ldq_17_bits_uop_ldq_idx;
      5'b10010:
        casez_tmp_239 = ldq_18_bits_uop_ldq_idx;
      5'b10011:
        casez_tmp_239 = ldq_19_bits_uop_ldq_idx;
      5'b10100:
        casez_tmp_239 = ldq_20_bits_uop_ldq_idx;
      5'b10101:
        casez_tmp_239 = ldq_21_bits_uop_ldq_idx;
      5'b10110:
        casez_tmp_239 = ldq_22_bits_uop_ldq_idx;
      5'b10111:
        casez_tmp_239 = ldq_23_bits_uop_ldq_idx;
      5'b11000:
        casez_tmp_239 = ldq_24_bits_uop_ldq_idx;
      5'b11001:
        casez_tmp_239 = ldq_25_bits_uop_ldq_idx;
      5'b11010:
        casez_tmp_239 = ldq_26_bits_uop_ldq_idx;
      5'b11011:
        casez_tmp_239 = ldq_27_bits_uop_ldq_idx;
      5'b11100:
        casez_tmp_239 = ldq_28_bits_uop_ldq_idx;
      5'b11101:
        casez_tmp_239 = ldq_29_bits_uop_ldq_idx;
      5'b11110:
        casez_tmp_239 = ldq_30_bits_uop_ldq_idx;
      default:
        casez_tmp_239 = ldq_31_bits_uop_ldq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_240 = ldq_0_bits_uop_stq_idx;
      5'b00001:
        casez_tmp_240 = ldq_1_bits_uop_stq_idx;
      5'b00010:
        casez_tmp_240 = ldq_2_bits_uop_stq_idx;
      5'b00011:
        casez_tmp_240 = ldq_3_bits_uop_stq_idx;
      5'b00100:
        casez_tmp_240 = ldq_4_bits_uop_stq_idx;
      5'b00101:
        casez_tmp_240 = ldq_5_bits_uop_stq_idx;
      5'b00110:
        casez_tmp_240 = ldq_6_bits_uop_stq_idx;
      5'b00111:
        casez_tmp_240 = ldq_7_bits_uop_stq_idx;
      5'b01000:
        casez_tmp_240 = ldq_8_bits_uop_stq_idx;
      5'b01001:
        casez_tmp_240 = ldq_9_bits_uop_stq_idx;
      5'b01010:
        casez_tmp_240 = ldq_10_bits_uop_stq_idx;
      5'b01011:
        casez_tmp_240 = ldq_11_bits_uop_stq_idx;
      5'b01100:
        casez_tmp_240 = ldq_12_bits_uop_stq_idx;
      5'b01101:
        casez_tmp_240 = ldq_13_bits_uop_stq_idx;
      5'b01110:
        casez_tmp_240 = ldq_14_bits_uop_stq_idx;
      5'b01111:
        casez_tmp_240 = ldq_15_bits_uop_stq_idx;
      5'b10000:
        casez_tmp_240 = ldq_16_bits_uop_stq_idx;
      5'b10001:
        casez_tmp_240 = ldq_17_bits_uop_stq_idx;
      5'b10010:
        casez_tmp_240 = ldq_18_bits_uop_stq_idx;
      5'b10011:
        casez_tmp_240 = ldq_19_bits_uop_stq_idx;
      5'b10100:
        casez_tmp_240 = ldq_20_bits_uop_stq_idx;
      5'b10101:
        casez_tmp_240 = ldq_21_bits_uop_stq_idx;
      5'b10110:
        casez_tmp_240 = ldq_22_bits_uop_stq_idx;
      5'b10111:
        casez_tmp_240 = ldq_23_bits_uop_stq_idx;
      5'b11000:
        casez_tmp_240 = ldq_24_bits_uop_stq_idx;
      5'b11001:
        casez_tmp_240 = ldq_25_bits_uop_stq_idx;
      5'b11010:
        casez_tmp_240 = ldq_26_bits_uop_stq_idx;
      5'b11011:
        casez_tmp_240 = ldq_27_bits_uop_stq_idx;
      5'b11100:
        casez_tmp_240 = ldq_28_bits_uop_stq_idx;
      5'b11101:
        casez_tmp_240 = ldq_29_bits_uop_stq_idx;
      5'b11110:
        casez_tmp_240 = ldq_30_bits_uop_stq_idx;
      default:
        casez_tmp_240 = ldq_31_bits_uop_stq_idx;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_241 = ldq_0_bits_uop_pdst;
      5'b00001:
        casez_tmp_241 = ldq_1_bits_uop_pdst;
      5'b00010:
        casez_tmp_241 = ldq_2_bits_uop_pdst;
      5'b00011:
        casez_tmp_241 = ldq_3_bits_uop_pdst;
      5'b00100:
        casez_tmp_241 = ldq_4_bits_uop_pdst;
      5'b00101:
        casez_tmp_241 = ldq_5_bits_uop_pdst;
      5'b00110:
        casez_tmp_241 = ldq_6_bits_uop_pdst;
      5'b00111:
        casez_tmp_241 = ldq_7_bits_uop_pdst;
      5'b01000:
        casez_tmp_241 = ldq_8_bits_uop_pdst;
      5'b01001:
        casez_tmp_241 = ldq_9_bits_uop_pdst;
      5'b01010:
        casez_tmp_241 = ldq_10_bits_uop_pdst;
      5'b01011:
        casez_tmp_241 = ldq_11_bits_uop_pdst;
      5'b01100:
        casez_tmp_241 = ldq_12_bits_uop_pdst;
      5'b01101:
        casez_tmp_241 = ldq_13_bits_uop_pdst;
      5'b01110:
        casez_tmp_241 = ldq_14_bits_uop_pdst;
      5'b01111:
        casez_tmp_241 = ldq_15_bits_uop_pdst;
      5'b10000:
        casez_tmp_241 = ldq_16_bits_uop_pdst;
      5'b10001:
        casez_tmp_241 = ldq_17_bits_uop_pdst;
      5'b10010:
        casez_tmp_241 = ldq_18_bits_uop_pdst;
      5'b10011:
        casez_tmp_241 = ldq_19_bits_uop_pdst;
      5'b10100:
        casez_tmp_241 = ldq_20_bits_uop_pdst;
      5'b10101:
        casez_tmp_241 = ldq_21_bits_uop_pdst;
      5'b10110:
        casez_tmp_241 = ldq_22_bits_uop_pdst;
      5'b10111:
        casez_tmp_241 = ldq_23_bits_uop_pdst;
      5'b11000:
        casez_tmp_241 = ldq_24_bits_uop_pdst;
      5'b11001:
        casez_tmp_241 = ldq_25_bits_uop_pdst;
      5'b11010:
        casez_tmp_241 = ldq_26_bits_uop_pdst;
      5'b11011:
        casez_tmp_241 = ldq_27_bits_uop_pdst;
      5'b11100:
        casez_tmp_241 = ldq_28_bits_uop_pdst;
      5'b11101:
        casez_tmp_241 = ldq_29_bits_uop_pdst;
      5'b11110:
        casez_tmp_241 = ldq_30_bits_uop_pdst;
      default:
        casez_tmp_241 = ldq_31_bits_uop_pdst;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_242 = ldq_0_bits_uop_mem_signed;
      5'b00001:
        casez_tmp_242 = ldq_1_bits_uop_mem_signed;
      5'b00010:
        casez_tmp_242 = ldq_2_bits_uop_mem_signed;
      5'b00011:
        casez_tmp_242 = ldq_3_bits_uop_mem_signed;
      5'b00100:
        casez_tmp_242 = ldq_4_bits_uop_mem_signed;
      5'b00101:
        casez_tmp_242 = ldq_5_bits_uop_mem_signed;
      5'b00110:
        casez_tmp_242 = ldq_6_bits_uop_mem_signed;
      5'b00111:
        casez_tmp_242 = ldq_7_bits_uop_mem_signed;
      5'b01000:
        casez_tmp_242 = ldq_8_bits_uop_mem_signed;
      5'b01001:
        casez_tmp_242 = ldq_9_bits_uop_mem_signed;
      5'b01010:
        casez_tmp_242 = ldq_10_bits_uop_mem_signed;
      5'b01011:
        casez_tmp_242 = ldq_11_bits_uop_mem_signed;
      5'b01100:
        casez_tmp_242 = ldq_12_bits_uop_mem_signed;
      5'b01101:
        casez_tmp_242 = ldq_13_bits_uop_mem_signed;
      5'b01110:
        casez_tmp_242 = ldq_14_bits_uop_mem_signed;
      5'b01111:
        casez_tmp_242 = ldq_15_bits_uop_mem_signed;
      5'b10000:
        casez_tmp_242 = ldq_16_bits_uop_mem_signed;
      5'b10001:
        casez_tmp_242 = ldq_17_bits_uop_mem_signed;
      5'b10010:
        casez_tmp_242 = ldq_18_bits_uop_mem_signed;
      5'b10011:
        casez_tmp_242 = ldq_19_bits_uop_mem_signed;
      5'b10100:
        casez_tmp_242 = ldq_20_bits_uop_mem_signed;
      5'b10101:
        casez_tmp_242 = ldq_21_bits_uop_mem_signed;
      5'b10110:
        casez_tmp_242 = ldq_22_bits_uop_mem_signed;
      5'b10111:
        casez_tmp_242 = ldq_23_bits_uop_mem_signed;
      5'b11000:
        casez_tmp_242 = ldq_24_bits_uop_mem_signed;
      5'b11001:
        casez_tmp_242 = ldq_25_bits_uop_mem_signed;
      5'b11010:
        casez_tmp_242 = ldq_26_bits_uop_mem_signed;
      5'b11011:
        casez_tmp_242 = ldq_27_bits_uop_mem_signed;
      5'b11100:
        casez_tmp_242 = ldq_28_bits_uop_mem_signed;
      5'b11101:
        casez_tmp_242 = ldq_29_bits_uop_mem_signed;
      5'b11110:
        casez_tmp_242 = ldq_30_bits_uop_mem_signed;
      default:
        casez_tmp_242 = ldq_31_bits_uop_mem_signed;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_243 = ldq_0_bits_uop_is_amo;
      5'b00001:
        casez_tmp_243 = ldq_1_bits_uop_is_amo;
      5'b00010:
        casez_tmp_243 = ldq_2_bits_uop_is_amo;
      5'b00011:
        casez_tmp_243 = ldq_3_bits_uop_is_amo;
      5'b00100:
        casez_tmp_243 = ldq_4_bits_uop_is_amo;
      5'b00101:
        casez_tmp_243 = ldq_5_bits_uop_is_amo;
      5'b00110:
        casez_tmp_243 = ldq_6_bits_uop_is_amo;
      5'b00111:
        casez_tmp_243 = ldq_7_bits_uop_is_amo;
      5'b01000:
        casez_tmp_243 = ldq_8_bits_uop_is_amo;
      5'b01001:
        casez_tmp_243 = ldq_9_bits_uop_is_amo;
      5'b01010:
        casez_tmp_243 = ldq_10_bits_uop_is_amo;
      5'b01011:
        casez_tmp_243 = ldq_11_bits_uop_is_amo;
      5'b01100:
        casez_tmp_243 = ldq_12_bits_uop_is_amo;
      5'b01101:
        casez_tmp_243 = ldq_13_bits_uop_is_amo;
      5'b01110:
        casez_tmp_243 = ldq_14_bits_uop_is_amo;
      5'b01111:
        casez_tmp_243 = ldq_15_bits_uop_is_amo;
      5'b10000:
        casez_tmp_243 = ldq_16_bits_uop_is_amo;
      5'b10001:
        casez_tmp_243 = ldq_17_bits_uop_is_amo;
      5'b10010:
        casez_tmp_243 = ldq_18_bits_uop_is_amo;
      5'b10011:
        casez_tmp_243 = ldq_19_bits_uop_is_amo;
      5'b10100:
        casez_tmp_243 = ldq_20_bits_uop_is_amo;
      5'b10101:
        casez_tmp_243 = ldq_21_bits_uop_is_amo;
      5'b10110:
        casez_tmp_243 = ldq_22_bits_uop_is_amo;
      5'b10111:
        casez_tmp_243 = ldq_23_bits_uop_is_amo;
      5'b11000:
        casez_tmp_243 = ldq_24_bits_uop_is_amo;
      5'b11001:
        casez_tmp_243 = ldq_25_bits_uop_is_amo;
      5'b11010:
        casez_tmp_243 = ldq_26_bits_uop_is_amo;
      5'b11011:
        casez_tmp_243 = ldq_27_bits_uop_is_amo;
      5'b11100:
        casez_tmp_243 = ldq_28_bits_uop_is_amo;
      5'b11101:
        casez_tmp_243 = ldq_29_bits_uop_is_amo;
      5'b11110:
        casez_tmp_243 = ldq_30_bits_uop_is_amo;
      default:
        casez_tmp_243 = ldq_31_bits_uop_is_amo;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_244 = ldq_0_bits_uop_uses_stq;
      5'b00001:
        casez_tmp_244 = ldq_1_bits_uop_uses_stq;
      5'b00010:
        casez_tmp_244 = ldq_2_bits_uop_uses_stq;
      5'b00011:
        casez_tmp_244 = ldq_3_bits_uop_uses_stq;
      5'b00100:
        casez_tmp_244 = ldq_4_bits_uop_uses_stq;
      5'b00101:
        casez_tmp_244 = ldq_5_bits_uop_uses_stq;
      5'b00110:
        casez_tmp_244 = ldq_6_bits_uop_uses_stq;
      5'b00111:
        casez_tmp_244 = ldq_7_bits_uop_uses_stq;
      5'b01000:
        casez_tmp_244 = ldq_8_bits_uop_uses_stq;
      5'b01001:
        casez_tmp_244 = ldq_9_bits_uop_uses_stq;
      5'b01010:
        casez_tmp_244 = ldq_10_bits_uop_uses_stq;
      5'b01011:
        casez_tmp_244 = ldq_11_bits_uop_uses_stq;
      5'b01100:
        casez_tmp_244 = ldq_12_bits_uop_uses_stq;
      5'b01101:
        casez_tmp_244 = ldq_13_bits_uop_uses_stq;
      5'b01110:
        casez_tmp_244 = ldq_14_bits_uop_uses_stq;
      5'b01111:
        casez_tmp_244 = ldq_15_bits_uop_uses_stq;
      5'b10000:
        casez_tmp_244 = ldq_16_bits_uop_uses_stq;
      5'b10001:
        casez_tmp_244 = ldq_17_bits_uop_uses_stq;
      5'b10010:
        casez_tmp_244 = ldq_18_bits_uop_uses_stq;
      5'b10011:
        casez_tmp_244 = ldq_19_bits_uop_uses_stq;
      5'b10100:
        casez_tmp_244 = ldq_20_bits_uop_uses_stq;
      5'b10101:
        casez_tmp_244 = ldq_21_bits_uop_uses_stq;
      5'b10110:
        casez_tmp_244 = ldq_22_bits_uop_uses_stq;
      5'b10111:
        casez_tmp_244 = ldq_23_bits_uop_uses_stq;
      5'b11000:
        casez_tmp_244 = ldq_24_bits_uop_uses_stq;
      5'b11001:
        casez_tmp_244 = ldq_25_bits_uop_uses_stq;
      5'b11010:
        casez_tmp_244 = ldq_26_bits_uop_uses_stq;
      5'b11011:
        casez_tmp_244 = ldq_27_bits_uop_uses_stq;
      5'b11100:
        casez_tmp_244 = ldq_28_bits_uop_uses_stq;
      5'b11101:
        casez_tmp_244 = ldq_29_bits_uop_uses_stq;
      5'b11110:
        casez_tmp_244 = ldq_30_bits_uop_uses_stq;
      default:
        casez_tmp_244 = ldq_31_bits_uop_uses_stq;
    endcase
  end // always @(*)
  always @(*) begin
    casez (wb_forward_ldq_idx_1)
      5'b00000:
        casez_tmp_245 = ldq_0_bits_uop_fp_val;
      5'b00001:
        casez_tmp_245 = ldq_1_bits_uop_fp_val;
      5'b00010:
        casez_tmp_245 = ldq_2_bits_uop_fp_val;
      5'b00011:
        casez_tmp_245 = ldq_3_bits_uop_fp_val;
      5'b00100:
        casez_tmp_245 = ldq_4_bits_uop_fp_val;
      5'b00101:
        casez_tmp_245 = ldq_5_bits_uop_fp_val;
      5'b00110:
        casez_tmp_245 = ldq_6_bits_uop_fp_val;
      5'b00111:
        casez_tmp_245 = ldq_7_bits_uop_fp_val;
      5'b01000:
        casez_tmp_245 = ldq_8_bits_uop_fp_val;
      5'b01001:
        casez_tmp_245 = ldq_9_bits_uop_fp_val;
      5'b01010:
        casez_tmp_245 = ldq_10_bits_uop_fp_val;
      5'b01011:
        casez_tmp_245 = ldq_11_bits_uop_fp_val;
      5'b01100:
        casez_tmp_245 = ldq_12_bits_uop_fp_val;
      5'b01101:
        casez_tmp_245 = ldq_13_bits_uop_fp_val;
      5'b01110:
        casez_tmp_245 = ldq_14_bits_uop_fp_val;
      5'b01111:
        casez_tmp_245 = ldq_15_bits_uop_fp_val;
      5'b10000:
        casez_tmp_245 = ldq_16_bits_uop_fp_val;
      5'b10001:
        casez_tmp_245 = ldq_17_bits_uop_fp_val;
      5'b10010:
        casez_tmp_245 = ldq_18_bits_uop_fp_val;
      5'b10011:
        casez_tmp_245 = ldq_19_bits_uop_fp_val;
      5'b10100:
        casez_tmp_245 = ldq_20_bits_uop_fp_val;
      5'b10101:
        casez_tmp_245 = ldq_21_bits_uop_fp_val;
      5'b10110:
        casez_tmp_245 = ldq_22_bits_uop_fp_val;
      5'b10111:
        casez_tmp_245 = ldq_23_bits_uop_fp_val;
      5'b11000:
        casez_tmp_245 = ldq_24_bits_uop_fp_val;
      5'b11001:
        casez_tmp_245 = ldq_25_bits_uop_fp_val;
      5'b11010:
        casez_tmp_245 = ldq_26_bits_uop_fp_val;
      5'b11011:
        casez_tmp_245 = ldq_27_bits_uop_fp_val;
      5'b11100:
        casez_tmp_245 = ldq_28_bits_uop_fp_val;
      5'b11101:
        casez_tmp_245 = ldq_29_bits_uop_fp_val;
      5'b11110:
        casez_tmp_245 = ldq_30_bits_uop_fp_val;
      default:
        casez_tmp_245 = ldq_31_bits_uop_fp_val;
    endcase
  end // always @(*)
  wire [31:0] io_core_exe_1_iresp_bits_data_zeroed = wb_forward_ld_addr_1[2] ? casez_tmp_233[63:32] : casez_tmp_233[31:0];
  wire        _ldq_bits_debug_wb_data_T_28 = casez_tmp_234 == 2'h2;
  wire [15:0] io_core_exe_1_iresp_bits_data_zeroed_1 = wb_forward_ld_addr_1[1] ? io_core_exe_1_iresp_bits_data_zeroed[31:16] : io_core_exe_1_iresp_bits_data_zeroed[15:0];
  wire        _ldq_bits_debug_wb_data_T_37 = casez_tmp_234 == 2'h1;
  wire [7:0]  io_core_exe_1_iresp_bits_data_zeroed_2 = wb_forward_ld_addr_1[0] ? io_core_exe_1_iresp_bits_data_zeroed_1[15:8] : io_core_exe_1_iresp_bits_data_zeroed_1[7:0];
  wire        _ldq_bits_debug_wb_data_T_46 = casez_tmp_234 == 2'h0;
  wire [31:0] io_core_exe_1_fresp_bits_data_zeroed = wb_forward_ld_addr_1[2] ? casez_tmp_233[63:32] : casez_tmp_233[31:0];
  wire [15:0] io_core_exe_1_fresp_bits_data_zeroed_1 = wb_forward_ld_addr_1[1] ? io_core_exe_1_fresp_bits_data_zeroed[31:16] : io_core_exe_1_fresp_bits_data_zeroed[15:0];
  wire [7:0]  io_core_exe_1_fresp_bits_data_zeroed_2 = wb_forward_ld_addr_1[0] ? io_core_exe_1_fresp_bits_data_zeroed_1[15:8] : io_core_exe_1_fresp_bits_data_zeroed_1[7:0];
  wire        _GEN_1185 = _GEN_1183 | ~_GEN_1184;
  wire        _io_core_exe_1_iresp_valid_output = _GEN_1185 ? io_dmem_resp_1_valid & (io_dmem_resp_1_bits_uop_uses_ldq ? send_iresp_1 : io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_is_amo) : casez_tmp_235 == 2'h0 & casez_tmp_236 & live_1;
  wire        _io_core_exe_1_fresp_valid_output = _GEN_1185 ? _GEN_1182 & send_fresp_1 : casez_tmp_235 == 2'h1 & casez_tmp_236 & live_1;
  reg         io_core_ld_miss_REG;
  reg         spec_ld_succeed_REG;
  reg  [4:0]  spec_ld_succeed_REG_1;
  reg         spec_ld_succeed_REG_2;
  reg  [4:0]  spec_ld_succeed_REG_3;
  wire [19:0] _GEN_1186 = io_core_brupdate_b1_mispredict_mask & stq_0_bits_uop_br_mask;
  wire [19:0] _GEN_1187 = io_core_brupdate_b1_mispredict_mask & stq_1_bits_uop_br_mask;
  wire [19:0] _GEN_1188 = io_core_brupdate_b1_mispredict_mask & stq_2_bits_uop_br_mask;
  wire [19:0] _GEN_1189 = io_core_brupdate_b1_mispredict_mask & stq_3_bits_uop_br_mask;
  wire [19:0] _GEN_1190 = io_core_brupdate_b1_mispredict_mask & stq_4_bits_uop_br_mask;
  wire [19:0] _GEN_1191 = io_core_brupdate_b1_mispredict_mask & stq_5_bits_uop_br_mask;
  wire [19:0] _GEN_1192 = io_core_brupdate_b1_mispredict_mask & stq_6_bits_uop_br_mask;
  wire [19:0] _GEN_1193 = io_core_brupdate_b1_mispredict_mask & stq_7_bits_uop_br_mask;
  wire [19:0] _GEN_1194 = io_core_brupdate_b1_mispredict_mask & stq_8_bits_uop_br_mask;
  wire [19:0] _GEN_1195 = io_core_brupdate_b1_mispredict_mask & stq_9_bits_uop_br_mask;
  wire [19:0] _GEN_1196 = io_core_brupdate_b1_mispredict_mask & stq_10_bits_uop_br_mask;
  wire [19:0] _GEN_1197 = io_core_brupdate_b1_mispredict_mask & stq_11_bits_uop_br_mask;
  wire [19:0] _GEN_1198 = io_core_brupdate_b1_mispredict_mask & stq_12_bits_uop_br_mask;
  wire [19:0] _GEN_1199 = io_core_brupdate_b1_mispredict_mask & stq_13_bits_uop_br_mask;
  wire [19:0] _GEN_1200 = io_core_brupdate_b1_mispredict_mask & stq_14_bits_uop_br_mask;
  wire [19:0] _GEN_1201 = io_core_brupdate_b1_mispredict_mask & stq_15_bits_uop_br_mask;
  wire [19:0] _GEN_1202 = io_core_brupdate_b1_mispredict_mask & stq_16_bits_uop_br_mask;
  wire [19:0] _GEN_1203 = io_core_brupdate_b1_mispredict_mask & stq_17_bits_uop_br_mask;
  wire [19:0] _GEN_1204 = io_core_brupdate_b1_mispredict_mask & stq_18_bits_uop_br_mask;
  wire [19:0] _GEN_1205 = io_core_brupdate_b1_mispredict_mask & stq_19_bits_uop_br_mask;
  wire [19:0] _GEN_1206 = io_core_brupdate_b1_mispredict_mask & stq_20_bits_uop_br_mask;
  wire [19:0] _GEN_1207 = io_core_brupdate_b1_mispredict_mask & stq_21_bits_uop_br_mask;
  wire [19:0] _GEN_1208 = io_core_brupdate_b1_mispredict_mask & stq_22_bits_uop_br_mask;
  wire [19:0] _GEN_1209 = io_core_brupdate_b1_mispredict_mask & stq_23_bits_uop_br_mask;
  wire [19:0] _GEN_1210 = io_core_brupdate_b1_mispredict_mask & stq_24_bits_uop_br_mask;
  wire [19:0] _GEN_1211 = io_core_brupdate_b1_mispredict_mask & stq_25_bits_uop_br_mask;
  wire [19:0] _GEN_1212 = io_core_brupdate_b1_mispredict_mask & stq_26_bits_uop_br_mask;
  wire [19:0] _GEN_1213 = io_core_brupdate_b1_mispredict_mask & stq_27_bits_uop_br_mask;
  wire [19:0] _GEN_1214 = io_core_brupdate_b1_mispredict_mask & stq_28_bits_uop_br_mask;
  wire [19:0] _GEN_1215 = io_core_brupdate_b1_mispredict_mask & stq_29_bits_uop_br_mask;
  wire [19:0] _GEN_1216 = io_core_brupdate_b1_mispredict_mask & stq_30_bits_uop_br_mask;
  wire [19:0] _GEN_1217 = io_core_brupdate_b1_mispredict_mask & stq_31_bits_uop_br_mask;
  wire        commit_store = io_core_commit_valids_0 & io_core_commit_uops_0_uses_stq;
  wire        commit_load = io_core_commit_valids_0 & io_core_commit_uops_0_uses_ldq;
  wire [4:0]  idx = commit_store ? stq_commit_head : ldq_head;
  wire [4:0]  _GEN_1218 = stq_commit_head + 5'h1;
  wire [4:0]  _GEN_1219 = commit_store ? _GEN_1218 : stq_commit_head;
  wire [4:0]  _GEN_1220 = ldq_head + 5'h1;
  wire [4:0]  _GEN_1221 = commit_load ? _GEN_1220 : ldq_head;
  wire        commit_store_1 = io_core_commit_valids_1 & io_core_commit_uops_1_uses_stq;
  wire        commit_load_1 = io_core_commit_valids_1 & io_core_commit_uops_1_uses_ldq;
  wire [4:0]  idx_1 = commit_store_1 ? _GEN_1219 : _GEN_1221;
  wire [4:0]  _GEN_1222 = _GEN_1219 + 5'h1;
  wire [4:0]  _GEN_1223 = commit_store_1 ? _GEN_1222 : _GEN_1219;
  wire [4:0]  _GEN_1224 = _GEN_1221 + 5'h1;
  wire [4:0]  _GEN_1225 = commit_load_1 ? _GEN_1224 : _GEN_1221;
  wire        commit_store_2 = io_core_commit_valids_2 & io_core_commit_uops_2_uses_stq;
  wire        commit_load_2 = io_core_commit_valids_2 & io_core_commit_uops_2_uses_ldq;
  wire [4:0]  idx_2 = commit_store_2 ? _GEN_1223 : _GEN_1225;
  wire [4:0]  _GEN_1226 = _GEN_1223 + 5'h1;
  wire [4:0]  _GEN_1227 = commit_store_2 ? _GEN_1226 : _GEN_1223;
  wire [4:0]  _GEN_1228 = _GEN_1225 + 5'h1;
  wire [4:0]  _GEN_1229 = commit_load_2 ? _GEN_1228 : _GEN_1225;
  wire        commit_store_3 = io_core_commit_valids_3 & io_core_commit_uops_3_uses_stq;
  wire        commit_load_3 = io_core_commit_valids_3 & io_core_commit_uops_3_uses_ldq;
  wire [4:0]  idx_3 = commit_store_3 ? _GEN_1227 : _GEN_1229;
  wire        _GEN_140185 = io_dmem_resp_0_valid & io_dmem_resp_0_bits_is_hella;
  wire        _GEN_1230 = io_dmem_nack_0_valid & io_dmem_nack_0_bits_is_hella;
  wire        _GEN_1231 = io_dmem_resp_1_valid & io_dmem_resp_1_bits_is_hella;
  wire        _GEN_1232 = io_dmem_nack_1_valid & io_dmem_nack_1_bits_is_hella;
  wire        _GEN_1233 = will_fire_hella_incoming_1 & dmem_req_fire_1;
  wire [2:0]  _GEN_140204 = _GEN_1177 & (_GEN_1231 | _GEN_140185) ? 3'h0 : hella_state;
  always @(*) begin
    casez (hella_state)
      3'b000:
        casez_tmp_246 = _GEN_140204;
      3'b001:
        casez_tmp_246 = io_hellacache_s1_kill ? (_GEN_1233 ? 3'h6 : 3'h0) : {2'h1, ~_GEN_1233};
      3'b010:
        casez_tmp_246 = {1'h1, |{hella_xcpt_ma_ld, hella_xcpt_ma_st, hella_xcpt_pf_ld, hella_xcpt_pf_st, hella_xcpt_gf_ld, hella_xcpt_gf_st, hella_xcpt_ae_ld, hella_xcpt_ae_st}, 1'h0};
      3'b011:
        casez_tmp_246 = 3'h0;
      3'b100:
        casez_tmp_246 = _GEN_1231 ? 3'h0 : _GEN_1232 ? 3'h5 : _GEN_140185 ? 3'h0 : _GEN_1230 ? 3'h5 : hella_state;
      3'b101:
        casez_tmp_246 = will_fire_hella_wakeup_1 & dmem_req_fire_1 ? 3'h4 : hella_state;
      3'b110:
        casez_tmp_246 = _GEN_140204;
      default:
        casez_tmp_246 = _GEN_140204;
    endcase
  end // always @(*)
  wire        _GEN_1234 = reset | io_core_exception;
  wire        _GEN_1235 = _GEN_1234 & reset;
  wire        _GEN_1236 = stq_execute_head < stq_head;
  wire [4:0]  _stq_execute_head_T_8 = stq_execute_head + 5'h1;
  wire [19:0] _clr_bsy_valid_0_T_22 = io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_0_bits_uop_br_mask;
  wire [19:0] _clr_bsy_valid_1_T_22 = io_core_brupdate_b1_mispredict_mask & mem_stq_incoming_e_1_bits_uop_br_mask;
  wire [31:0] _ldq_31_bits_st_dep_mask_T = 32'h1 << stq_head;
  wire        _GEN_1237 = stq_head == 5'h1;
  wire        _GEN_1238 = stq_head == 5'h2;
  wire        _GEN_1239 = stq_head == 5'h3;
  wire        _GEN_1240 = stq_head == 5'h4;
  wire        _GEN_1241 = stq_head == 5'h5;
  wire        _GEN_1242 = stq_head == 5'h6;
  wire        _GEN_1243 = stq_head == 5'h7;
  wire        _GEN_1244 = stq_head == 5'h8;
  wire        _GEN_1245 = stq_head == 5'h9;
  wire        _GEN_1246 = stq_head == 5'hA;
  wire        _GEN_1247 = stq_head == 5'hB;
  wire        _GEN_1248 = stq_head == 5'hC;
  wire        _GEN_1249 = stq_head == 5'hD;
  wire        _GEN_1250 = stq_head == 5'hE;
  wire        _GEN_1251 = stq_head == 5'hF;
  wire        _GEN_1252 = stq_head == 5'h10;
  wire        _GEN_1253 = stq_head == 5'h11;
  wire        _GEN_1254 = stq_head == 5'h12;
  wire        _GEN_1255 = stq_head == 5'h13;
  wire        _GEN_1256 = stq_head == 5'h14;
  wire        _GEN_1257 = stq_head == 5'h15;
  wire        _GEN_1258 = stq_head == 5'h16;
  wire        _GEN_1259 = stq_head == 5'h17;
  wire        _GEN_1260 = stq_head == 5'h18;
  wire        _GEN_1261 = stq_head == 5'h19;
  wire        _GEN_1262 = stq_head == 5'h1A;
  wire        _GEN_1263 = stq_head == 5'h1B;
  wire        _GEN_1264 = stq_head == 5'h1C;
  wire        _GEN_1265 = stq_head == 5'h1D;
  wire        _GEN_1266 = stq_head == 5'h1E;
  wire        clear_store = _GEN & (casez_tmp_2 ? io_dmem_ordered : casez_tmp_3);
  wire [31:0] _GEN_1267 = {32{~clear_store}};
  wire [31:0] next_live_store_mask = (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & live_store_mask;
  wire        _GEN_1268 = dis_ld_val | ~_GEN_2;
  wire        _GEN_1269 = dis_ld_val | ~_GEN_3;
  wire        _GEN_1270 = dis_ld_val | ~_GEN_4;
  wire        _GEN_1271 = dis_ld_val | ~_GEN_5;
  wire        _GEN_1272 = dis_ld_val | ~_GEN_6;
  wire        _GEN_1273 = dis_ld_val | ~_GEN_7;
  wire        _GEN_1274 = dis_ld_val | ~_GEN_8;
  wire        _GEN_1275 = dis_ld_val | ~_GEN_9;
  wire        _GEN_1276 = dis_ld_val | ~_GEN_10;
  wire        _GEN_1277 = dis_ld_val | ~_GEN_11;
  wire        _GEN_1278 = dis_ld_val | ~_GEN_12;
  wire        _GEN_1279 = dis_ld_val | ~_GEN_13;
  wire        _GEN_1280 = dis_ld_val | ~_GEN_14;
  wire        _GEN_1281 = dis_ld_val | ~_GEN_15;
  wire        _GEN_1282 = dis_ld_val | ~_GEN_16;
  wire        _GEN_1283 = dis_ld_val | ~_GEN_17;
  wire        _GEN_1284 = dis_ld_val | ~_GEN_18;
  wire        _GEN_1285 = dis_ld_val | ~_GEN_19;
  wire        _GEN_1286 = dis_ld_val | ~_GEN_20;
  wire        _GEN_1287 = dis_ld_val | ~_GEN_21;
  wire        _GEN_1288 = dis_ld_val | ~_GEN_22;
  wire        _GEN_1289 = dis_ld_val | ~_GEN_23;
  wire        _GEN_1290 = dis_ld_val | ~_GEN_24;
  wire        _GEN_1291 = dis_ld_val | ~_GEN_25;
  wire        _GEN_1292 = dis_ld_val | ~_GEN_26;
  wire        _GEN_1293 = dis_ld_val | ~_GEN_27;
  wire        _GEN_1294 = dis_ld_val | ~_GEN_28;
  wire        _GEN_1295 = dis_ld_val | ~_GEN_29;
  wire        _GEN_1296 = dis_ld_val | ~_GEN_30;
  wire        _GEN_1297 = dis_ld_val | ~_GEN_31;
  wire        _GEN_1298 = dis_ld_val | ~_GEN_32;
  wire        _GEN_1299 = dis_ld_val | ~_GEN_33;
  wire [31:0] _ldq_T_35_bits_st_dep_mask = {32{dis_st_val}} & 32'h1 << stq_tail | next_live_store_mask;
  wire        _GEN_1300 = _GEN_69 | _GEN_34;
  wire        _GEN_1301 = _GEN_70 | _GEN_35;
  wire        _GEN_1302 = _GEN_71 | _GEN_36;
  wire        _GEN_1303 = _GEN_72 | _GEN_37;
  wire        _GEN_1304 = _GEN_73 | _GEN_38;
  wire        _GEN_1305 = _GEN_74 | _GEN_39;
  wire        _GEN_1306 = _GEN_75 | _GEN_40;
  wire        _GEN_1307 = _GEN_76 | _GEN_41;
  wire        _GEN_1308 = _GEN_77 | _GEN_42;
  wire        _GEN_1309 = _GEN_78 | _GEN_43;
  wire        _GEN_1310 = _GEN_79 | _GEN_44;
  wire        _GEN_1311 = _GEN_80 | _GEN_45;
  wire        _GEN_1312 = _GEN_81 | _GEN_46;
  wire        _GEN_1313 = _GEN_82 | _GEN_47;
  wire        _GEN_1314 = _GEN_83 | _GEN_48;
  wire        _GEN_1315 = _GEN_84 | _GEN_49;
  wire        _GEN_1316 = _GEN_85 | _GEN_50;
  wire        _GEN_1317 = _GEN_86 | _GEN_51;
  wire        _GEN_1318 = _GEN_87 | _GEN_52;
  wire        _GEN_1319 = _GEN_88 | _GEN_53;
  wire        _GEN_1320 = _GEN_89 | _GEN_54;
  wire        _GEN_1321 = _GEN_90 | _GEN_55;
  wire        _GEN_1322 = _GEN_91 | _GEN_56;
  wire        _GEN_1323 = _GEN_92 | _GEN_57;
  wire        _GEN_1324 = _GEN_93 | _GEN_58;
  wire        _GEN_1325 = _GEN_94 | _GEN_59;
  wire        _GEN_1326 = _GEN_95 | _GEN_60;
  wire        _GEN_1327 = _GEN_96 | _GEN_61;
  wire        _GEN_1328 = _GEN_97 | _GEN_62;
  wire        _GEN_1329 = _GEN_98 | _GEN_63;
  wire        _GEN_1330 = _GEN_99 | _GEN_64;
  wire        _GEN_1331 = (&_GEN_66) | _GEN_65;
  wire        _GEN_22080 = dis_ld_val_1 ? _GEN_1300 | ldq_0_valid : _GEN_34 | ldq_0_valid;
  wire        _GEN_22081 = dis_ld_val_1 ? _GEN_1301 | ldq_1_valid : _GEN_35 | ldq_1_valid;
  wire        _GEN_22082 = dis_ld_val_1 ? _GEN_1302 | ldq_2_valid : _GEN_36 | ldq_2_valid;
  wire        _GEN_22083 = dis_ld_val_1 ? _GEN_1303 | ldq_3_valid : _GEN_37 | ldq_3_valid;
  wire        _GEN_22084 = dis_ld_val_1 ? _GEN_1304 | ldq_4_valid : _GEN_38 | ldq_4_valid;
  wire        _GEN_22085 = dis_ld_val_1 ? _GEN_1305 | ldq_5_valid : _GEN_39 | ldq_5_valid;
  wire        _GEN_22086 = dis_ld_val_1 ? _GEN_1306 | ldq_6_valid : _GEN_40 | ldq_6_valid;
  wire        _GEN_22087 = dis_ld_val_1 ? _GEN_1307 | ldq_7_valid : _GEN_41 | ldq_7_valid;
  wire        _GEN_22088 = dis_ld_val_1 ? _GEN_1308 | ldq_8_valid : _GEN_42 | ldq_8_valid;
  wire        _GEN_22089 = dis_ld_val_1 ? _GEN_1309 | ldq_9_valid : _GEN_43 | ldq_9_valid;
  wire        _GEN_22090 = dis_ld_val_1 ? _GEN_1310 | ldq_10_valid : _GEN_44 | ldq_10_valid;
  wire        _GEN_22091 = dis_ld_val_1 ? _GEN_1311 | ldq_11_valid : _GEN_45 | ldq_11_valid;
  wire        _GEN_22092 = dis_ld_val_1 ? _GEN_1312 | ldq_12_valid : _GEN_46 | ldq_12_valid;
  wire        _GEN_22093 = dis_ld_val_1 ? _GEN_1313 | ldq_13_valid : _GEN_47 | ldq_13_valid;
  wire        _GEN_22094 = dis_ld_val_1 ? _GEN_1314 | ldq_14_valid : _GEN_48 | ldq_14_valid;
  wire        _GEN_22095 = dis_ld_val_1 ? _GEN_1315 | ldq_15_valid : _GEN_49 | ldq_15_valid;
  wire        _GEN_22096 = dis_ld_val_1 ? _GEN_1316 | ldq_16_valid : _GEN_50 | ldq_16_valid;
  wire        _GEN_22097 = dis_ld_val_1 ? _GEN_1317 | ldq_17_valid : _GEN_51 | ldq_17_valid;
  wire        _GEN_22098 = dis_ld_val_1 ? _GEN_1318 | ldq_18_valid : _GEN_52 | ldq_18_valid;
  wire        _GEN_22099 = dis_ld_val_1 ? _GEN_1319 | ldq_19_valid : _GEN_53 | ldq_19_valid;
  wire        _GEN_22100 = dis_ld_val_1 ? _GEN_1320 | ldq_20_valid : _GEN_54 | ldq_20_valid;
  wire        _GEN_22101 = dis_ld_val_1 ? _GEN_1321 | ldq_21_valid : _GEN_55 | ldq_21_valid;
  wire        _GEN_22102 = dis_ld_val_1 ? _GEN_1322 | ldq_22_valid : _GEN_56 | ldq_22_valid;
  wire        _GEN_22103 = dis_ld_val_1 ? _GEN_1323 | ldq_23_valid : _GEN_57 | ldq_23_valid;
  wire        _GEN_22104 = dis_ld_val_1 ? _GEN_1324 | ldq_24_valid : _GEN_58 | ldq_24_valid;
  wire        _GEN_22105 = dis_ld_val_1 ? _GEN_1325 | ldq_25_valid : _GEN_59 | ldq_25_valid;
  wire        _GEN_22106 = dis_ld_val_1 ? _GEN_1326 | ldq_26_valid : _GEN_60 | ldq_26_valid;
  wire        _GEN_22107 = dis_ld_val_1 ? _GEN_1327 | ldq_27_valid : _GEN_61 | ldq_27_valid;
  wire        _GEN_22108 = dis_ld_val_1 ? _GEN_1328 | ldq_28_valid : _GEN_62 | ldq_28_valid;
  wire        _GEN_22109 = dis_ld_val_1 ? _GEN_1329 | ldq_29_valid : _GEN_63 | ldq_29_valid;
  wire        _GEN_22110 = dis_ld_val_1 ? _GEN_1330 | ldq_30_valid : _GEN_64 | ldq_30_valid;
  wire        _GEN_22111 = dis_ld_val_1 ? _GEN_1331 | ldq_31_valid : _GEN_65 | ldq_31_valid;
  wire        _GEN_24704 = dis_ld_val_1 ? ~_GEN_1300 & ldq_0_bits_addr_valid : ~_GEN_34 & ldq_0_bits_addr_valid;
  wire        _GEN_24705 = dis_ld_val_1 ? ~_GEN_1301 & ldq_1_bits_addr_valid : ~_GEN_35 & ldq_1_bits_addr_valid;
  wire        _GEN_24706 = dis_ld_val_1 ? ~_GEN_1302 & ldq_2_bits_addr_valid : ~_GEN_36 & ldq_2_bits_addr_valid;
  wire        _GEN_24707 = dis_ld_val_1 ? ~_GEN_1303 & ldq_3_bits_addr_valid : ~_GEN_37 & ldq_3_bits_addr_valid;
  wire        _GEN_24708 = dis_ld_val_1 ? ~_GEN_1304 & ldq_4_bits_addr_valid : ~_GEN_38 & ldq_4_bits_addr_valid;
  wire        _GEN_24709 = dis_ld_val_1 ? ~_GEN_1305 & ldq_5_bits_addr_valid : ~_GEN_39 & ldq_5_bits_addr_valid;
  wire        _GEN_24710 = dis_ld_val_1 ? ~_GEN_1306 & ldq_6_bits_addr_valid : ~_GEN_40 & ldq_6_bits_addr_valid;
  wire        _GEN_24711 = dis_ld_val_1 ? ~_GEN_1307 & ldq_7_bits_addr_valid : ~_GEN_41 & ldq_7_bits_addr_valid;
  wire        _GEN_24712 = dis_ld_val_1 ? ~_GEN_1308 & ldq_8_bits_addr_valid : ~_GEN_42 & ldq_8_bits_addr_valid;
  wire        _GEN_24713 = dis_ld_val_1 ? ~_GEN_1309 & ldq_9_bits_addr_valid : ~_GEN_43 & ldq_9_bits_addr_valid;
  wire        _GEN_24714 = dis_ld_val_1 ? ~_GEN_1310 & ldq_10_bits_addr_valid : ~_GEN_44 & ldq_10_bits_addr_valid;
  wire        _GEN_24715 = dis_ld_val_1 ? ~_GEN_1311 & ldq_11_bits_addr_valid : ~_GEN_45 & ldq_11_bits_addr_valid;
  wire        _GEN_24716 = dis_ld_val_1 ? ~_GEN_1312 & ldq_12_bits_addr_valid : ~_GEN_46 & ldq_12_bits_addr_valid;
  wire        _GEN_24717 = dis_ld_val_1 ? ~_GEN_1313 & ldq_13_bits_addr_valid : ~_GEN_47 & ldq_13_bits_addr_valid;
  wire        _GEN_24718 = dis_ld_val_1 ? ~_GEN_1314 & ldq_14_bits_addr_valid : ~_GEN_48 & ldq_14_bits_addr_valid;
  wire        _GEN_24719 = dis_ld_val_1 ? ~_GEN_1315 & ldq_15_bits_addr_valid : ~_GEN_49 & ldq_15_bits_addr_valid;
  wire        _GEN_24720 = dis_ld_val_1 ? ~_GEN_1316 & ldq_16_bits_addr_valid : ~_GEN_50 & ldq_16_bits_addr_valid;
  wire        _GEN_24721 = dis_ld_val_1 ? ~_GEN_1317 & ldq_17_bits_addr_valid : ~_GEN_51 & ldq_17_bits_addr_valid;
  wire        _GEN_24722 = dis_ld_val_1 ? ~_GEN_1318 & ldq_18_bits_addr_valid : ~_GEN_52 & ldq_18_bits_addr_valid;
  wire        _GEN_24723 = dis_ld_val_1 ? ~_GEN_1319 & ldq_19_bits_addr_valid : ~_GEN_53 & ldq_19_bits_addr_valid;
  wire        _GEN_24724 = dis_ld_val_1 ? ~_GEN_1320 & ldq_20_bits_addr_valid : ~_GEN_54 & ldq_20_bits_addr_valid;
  wire        _GEN_24725 = dis_ld_val_1 ? ~_GEN_1321 & ldq_21_bits_addr_valid : ~_GEN_55 & ldq_21_bits_addr_valid;
  wire        _GEN_24726 = dis_ld_val_1 ? ~_GEN_1322 & ldq_22_bits_addr_valid : ~_GEN_56 & ldq_22_bits_addr_valid;
  wire        _GEN_24727 = dis_ld_val_1 ? ~_GEN_1323 & ldq_23_bits_addr_valid : ~_GEN_57 & ldq_23_bits_addr_valid;
  wire        _GEN_24728 = dis_ld_val_1 ? ~_GEN_1324 & ldq_24_bits_addr_valid : ~_GEN_58 & ldq_24_bits_addr_valid;
  wire        _GEN_24729 = dis_ld_val_1 ? ~_GEN_1325 & ldq_25_bits_addr_valid : ~_GEN_59 & ldq_25_bits_addr_valid;
  wire        _GEN_24730 = dis_ld_val_1 ? ~_GEN_1326 & ldq_26_bits_addr_valid : ~_GEN_60 & ldq_26_bits_addr_valid;
  wire        _GEN_24731 = dis_ld_val_1 ? ~_GEN_1327 & ldq_27_bits_addr_valid : ~_GEN_61 & ldq_27_bits_addr_valid;
  wire        _GEN_24732 = dis_ld_val_1 ? ~_GEN_1328 & ldq_28_bits_addr_valid : ~_GEN_62 & ldq_28_bits_addr_valid;
  wire        _GEN_24733 = dis_ld_val_1 ? ~_GEN_1329 & ldq_29_bits_addr_valid : ~_GEN_63 & ldq_29_bits_addr_valid;
  wire        _GEN_24734 = dis_ld_val_1 ? ~_GEN_1330 & ldq_30_bits_addr_valid : ~_GEN_64 & ldq_30_bits_addr_valid;
  wire        _GEN_24735 = dis_ld_val_1 ? ~_GEN_1331 & ldq_31_bits_addr_valid : ~_GEN_65 & ldq_31_bits_addr_valid;
  wire        _GEN_24736 = dis_ld_val_1 ? ~_GEN_1300 & ldq_0_bits_executed : ~_GEN_34 & ldq_0_bits_executed;
  wire        _GEN_24737 = dis_ld_val_1 ? ~_GEN_1301 & ldq_1_bits_executed : ~_GEN_35 & ldq_1_bits_executed;
  wire        _GEN_24738 = dis_ld_val_1 ? ~_GEN_1302 & ldq_2_bits_executed : ~_GEN_36 & ldq_2_bits_executed;
  wire        _GEN_24739 = dis_ld_val_1 ? ~_GEN_1303 & ldq_3_bits_executed : ~_GEN_37 & ldq_3_bits_executed;
  wire        _GEN_24740 = dis_ld_val_1 ? ~_GEN_1304 & ldq_4_bits_executed : ~_GEN_38 & ldq_4_bits_executed;
  wire        _GEN_24741 = dis_ld_val_1 ? ~_GEN_1305 & ldq_5_bits_executed : ~_GEN_39 & ldq_5_bits_executed;
  wire        _GEN_24742 = dis_ld_val_1 ? ~_GEN_1306 & ldq_6_bits_executed : ~_GEN_40 & ldq_6_bits_executed;
  wire        _GEN_24743 = dis_ld_val_1 ? ~_GEN_1307 & ldq_7_bits_executed : ~_GEN_41 & ldq_7_bits_executed;
  wire        _GEN_24744 = dis_ld_val_1 ? ~_GEN_1308 & ldq_8_bits_executed : ~_GEN_42 & ldq_8_bits_executed;
  wire        _GEN_24745 = dis_ld_val_1 ? ~_GEN_1309 & ldq_9_bits_executed : ~_GEN_43 & ldq_9_bits_executed;
  wire        _GEN_24746 = dis_ld_val_1 ? ~_GEN_1310 & ldq_10_bits_executed : ~_GEN_44 & ldq_10_bits_executed;
  wire        _GEN_24747 = dis_ld_val_1 ? ~_GEN_1311 & ldq_11_bits_executed : ~_GEN_45 & ldq_11_bits_executed;
  wire        _GEN_24748 = dis_ld_val_1 ? ~_GEN_1312 & ldq_12_bits_executed : ~_GEN_46 & ldq_12_bits_executed;
  wire        _GEN_24749 = dis_ld_val_1 ? ~_GEN_1313 & ldq_13_bits_executed : ~_GEN_47 & ldq_13_bits_executed;
  wire        _GEN_24750 = dis_ld_val_1 ? ~_GEN_1314 & ldq_14_bits_executed : ~_GEN_48 & ldq_14_bits_executed;
  wire        _GEN_24751 = dis_ld_val_1 ? ~_GEN_1315 & ldq_15_bits_executed : ~_GEN_49 & ldq_15_bits_executed;
  wire        _GEN_24752 = dis_ld_val_1 ? ~_GEN_1316 & ldq_16_bits_executed : ~_GEN_50 & ldq_16_bits_executed;
  wire        _GEN_24753 = dis_ld_val_1 ? ~_GEN_1317 & ldq_17_bits_executed : ~_GEN_51 & ldq_17_bits_executed;
  wire        _GEN_24754 = dis_ld_val_1 ? ~_GEN_1318 & ldq_18_bits_executed : ~_GEN_52 & ldq_18_bits_executed;
  wire        _GEN_24755 = dis_ld_val_1 ? ~_GEN_1319 & ldq_19_bits_executed : ~_GEN_53 & ldq_19_bits_executed;
  wire        _GEN_24756 = dis_ld_val_1 ? ~_GEN_1320 & ldq_20_bits_executed : ~_GEN_54 & ldq_20_bits_executed;
  wire        _GEN_24757 = dis_ld_val_1 ? ~_GEN_1321 & ldq_21_bits_executed : ~_GEN_55 & ldq_21_bits_executed;
  wire        _GEN_24758 = dis_ld_val_1 ? ~_GEN_1322 & ldq_22_bits_executed : ~_GEN_56 & ldq_22_bits_executed;
  wire        _GEN_24759 = dis_ld_val_1 ? ~_GEN_1323 & ldq_23_bits_executed : ~_GEN_57 & ldq_23_bits_executed;
  wire        _GEN_24760 = dis_ld_val_1 ? ~_GEN_1324 & ldq_24_bits_executed : ~_GEN_58 & ldq_24_bits_executed;
  wire        _GEN_24761 = dis_ld_val_1 ? ~_GEN_1325 & ldq_25_bits_executed : ~_GEN_59 & ldq_25_bits_executed;
  wire        _GEN_24762 = dis_ld_val_1 ? ~_GEN_1326 & ldq_26_bits_executed : ~_GEN_60 & ldq_26_bits_executed;
  wire        _GEN_24763 = dis_ld_val_1 ? ~_GEN_1327 & ldq_27_bits_executed : ~_GEN_61 & ldq_27_bits_executed;
  wire        _GEN_24764 = dis_ld_val_1 ? ~_GEN_1328 & ldq_28_bits_executed : ~_GEN_62 & ldq_28_bits_executed;
  wire        _GEN_24765 = dis_ld_val_1 ? ~_GEN_1329 & ldq_29_bits_executed : ~_GEN_63 & ldq_29_bits_executed;
  wire        _GEN_24766 = dis_ld_val_1 ? ~_GEN_1330 & ldq_30_bits_executed : ~_GEN_64 & ldq_30_bits_executed;
  wire        _GEN_24767 = dis_ld_val_1 ? ~_GEN_1331 & ldq_31_bits_executed : ~_GEN_65 & ldq_31_bits_executed;
  wire        _GEN_24768 = dis_ld_val_1 ? ~_GEN_1300 & ldq_0_bits_succeeded : ~_GEN_34 & ldq_0_bits_succeeded;
  wire        _GEN_24769 = dis_ld_val_1 ? ~_GEN_1301 & ldq_1_bits_succeeded : ~_GEN_35 & ldq_1_bits_succeeded;
  wire        _GEN_24770 = dis_ld_val_1 ? ~_GEN_1302 & ldq_2_bits_succeeded : ~_GEN_36 & ldq_2_bits_succeeded;
  wire        _GEN_24771 = dis_ld_val_1 ? ~_GEN_1303 & ldq_3_bits_succeeded : ~_GEN_37 & ldq_3_bits_succeeded;
  wire        _GEN_24772 = dis_ld_val_1 ? ~_GEN_1304 & ldq_4_bits_succeeded : ~_GEN_38 & ldq_4_bits_succeeded;
  wire        _GEN_24773 = dis_ld_val_1 ? ~_GEN_1305 & ldq_5_bits_succeeded : ~_GEN_39 & ldq_5_bits_succeeded;
  wire        _GEN_24774 = dis_ld_val_1 ? ~_GEN_1306 & ldq_6_bits_succeeded : ~_GEN_40 & ldq_6_bits_succeeded;
  wire        _GEN_24775 = dis_ld_val_1 ? ~_GEN_1307 & ldq_7_bits_succeeded : ~_GEN_41 & ldq_7_bits_succeeded;
  wire        _GEN_24776 = dis_ld_val_1 ? ~_GEN_1308 & ldq_8_bits_succeeded : ~_GEN_42 & ldq_8_bits_succeeded;
  wire        _GEN_24777 = dis_ld_val_1 ? ~_GEN_1309 & ldq_9_bits_succeeded : ~_GEN_43 & ldq_9_bits_succeeded;
  wire        _GEN_24778 = dis_ld_val_1 ? ~_GEN_1310 & ldq_10_bits_succeeded : ~_GEN_44 & ldq_10_bits_succeeded;
  wire        _GEN_24779 = dis_ld_val_1 ? ~_GEN_1311 & ldq_11_bits_succeeded : ~_GEN_45 & ldq_11_bits_succeeded;
  wire        _GEN_24780 = dis_ld_val_1 ? ~_GEN_1312 & ldq_12_bits_succeeded : ~_GEN_46 & ldq_12_bits_succeeded;
  wire        _GEN_24781 = dis_ld_val_1 ? ~_GEN_1313 & ldq_13_bits_succeeded : ~_GEN_47 & ldq_13_bits_succeeded;
  wire        _GEN_24782 = dis_ld_val_1 ? ~_GEN_1314 & ldq_14_bits_succeeded : ~_GEN_48 & ldq_14_bits_succeeded;
  wire        _GEN_24783 = dis_ld_val_1 ? ~_GEN_1315 & ldq_15_bits_succeeded : ~_GEN_49 & ldq_15_bits_succeeded;
  wire        _GEN_24784 = dis_ld_val_1 ? ~_GEN_1316 & ldq_16_bits_succeeded : ~_GEN_50 & ldq_16_bits_succeeded;
  wire        _GEN_24785 = dis_ld_val_1 ? ~_GEN_1317 & ldq_17_bits_succeeded : ~_GEN_51 & ldq_17_bits_succeeded;
  wire        _GEN_24786 = dis_ld_val_1 ? ~_GEN_1318 & ldq_18_bits_succeeded : ~_GEN_52 & ldq_18_bits_succeeded;
  wire        _GEN_24787 = dis_ld_val_1 ? ~_GEN_1319 & ldq_19_bits_succeeded : ~_GEN_53 & ldq_19_bits_succeeded;
  wire        _GEN_24788 = dis_ld_val_1 ? ~_GEN_1320 & ldq_20_bits_succeeded : ~_GEN_54 & ldq_20_bits_succeeded;
  wire        _GEN_24789 = dis_ld_val_1 ? ~_GEN_1321 & ldq_21_bits_succeeded : ~_GEN_55 & ldq_21_bits_succeeded;
  wire        _GEN_24790 = dis_ld_val_1 ? ~_GEN_1322 & ldq_22_bits_succeeded : ~_GEN_56 & ldq_22_bits_succeeded;
  wire        _GEN_24791 = dis_ld_val_1 ? ~_GEN_1323 & ldq_23_bits_succeeded : ~_GEN_57 & ldq_23_bits_succeeded;
  wire        _GEN_24792 = dis_ld_val_1 ? ~_GEN_1324 & ldq_24_bits_succeeded : ~_GEN_58 & ldq_24_bits_succeeded;
  wire        _GEN_24793 = dis_ld_val_1 ? ~_GEN_1325 & ldq_25_bits_succeeded : ~_GEN_59 & ldq_25_bits_succeeded;
  wire        _GEN_24794 = dis_ld_val_1 ? ~_GEN_1326 & ldq_26_bits_succeeded : ~_GEN_60 & ldq_26_bits_succeeded;
  wire        _GEN_24795 = dis_ld_val_1 ? ~_GEN_1327 & ldq_27_bits_succeeded : ~_GEN_61 & ldq_27_bits_succeeded;
  wire        _GEN_24796 = dis_ld_val_1 ? ~_GEN_1328 & ldq_28_bits_succeeded : ~_GEN_62 & ldq_28_bits_succeeded;
  wire        _GEN_24797 = dis_ld_val_1 ? ~_GEN_1329 & ldq_29_bits_succeeded : ~_GEN_63 & ldq_29_bits_succeeded;
  wire        _GEN_24798 = dis_ld_val_1 ? ~_GEN_1330 & ldq_30_bits_succeeded : ~_GEN_64 & ldq_30_bits_succeeded;
  wire        _GEN_24799 = dis_ld_val_1 ? ~_GEN_1331 & ldq_31_bits_succeeded : ~_GEN_65 & ldq_31_bits_succeeded;
  wire        _GEN_24800 = dis_ld_val_1 ? ~_GEN_1300 & ldq_0_bits_order_fail : ~_GEN_34 & ldq_0_bits_order_fail;
  wire        _GEN_24801 = dis_ld_val_1 ? ~_GEN_1301 & ldq_1_bits_order_fail : ~_GEN_35 & ldq_1_bits_order_fail;
  wire        _GEN_24802 = dis_ld_val_1 ? ~_GEN_1302 & ldq_2_bits_order_fail : ~_GEN_36 & ldq_2_bits_order_fail;
  wire        _GEN_24803 = dis_ld_val_1 ? ~_GEN_1303 & ldq_3_bits_order_fail : ~_GEN_37 & ldq_3_bits_order_fail;
  wire        _GEN_24804 = dis_ld_val_1 ? ~_GEN_1304 & ldq_4_bits_order_fail : ~_GEN_38 & ldq_4_bits_order_fail;
  wire        _GEN_24805 = dis_ld_val_1 ? ~_GEN_1305 & ldq_5_bits_order_fail : ~_GEN_39 & ldq_5_bits_order_fail;
  wire        _GEN_24806 = dis_ld_val_1 ? ~_GEN_1306 & ldq_6_bits_order_fail : ~_GEN_40 & ldq_6_bits_order_fail;
  wire        _GEN_24807 = dis_ld_val_1 ? ~_GEN_1307 & ldq_7_bits_order_fail : ~_GEN_41 & ldq_7_bits_order_fail;
  wire        _GEN_24808 = dis_ld_val_1 ? ~_GEN_1308 & ldq_8_bits_order_fail : ~_GEN_42 & ldq_8_bits_order_fail;
  wire        _GEN_24809 = dis_ld_val_1 ? ~_GEN_1309 & ldq_9_bits_order_fail : ~_GEN_43 & ldq_9_bits_order_fail;
  wire        _GEN_24810 = dis_ld_val_1 ? ~_GEN_1310 & ldq_10_bits_order_fail : ~_GEN_44 & ldq_10_bits_order_fail;
  wire        _GEN_24811 = dis_ld_val_1 ? ~_GEN_1311 & ldq_11_bits_order_fail : ~_GEN_45 & ldq_11_bits_order_fail;
  wire        _GEN_24812 = dis_ld_val_1 ? ~_GEN_1312 & ldq_12_bits_order_fail : ~_GEN_46 & ldq_12_bits_order_fail;
  wire        _GEN_24813 = dis_ld_val_1 ? ~_GEN_1313 & ldq_13_bits_order_fail : ~_GEN_47 & ldq_13_bits_order_fail;
  wire        _GEN_24814 = dis_ld_val_1 ? ~_GEN_1314 & ldq_14_bits_order_fail : ~_GEN_48 & ldq_14_bits_order_fail;
  wire        _GEN_24815 = dis_ld_val_1 ? ~_GEN_1315 & ldq_15_bits_order_fail : ~_GEN_49 & ldq_15_bits_order_fail;
  wire        _GEN_24816 = dis_ld_val_1 ? ~_GEN_1316 & ldq_16_bits_order_fail : ~_GEN_50 & ldq_16_bits_order_fail;
  wire        _GEN_24817 = dis_ld_val_1 ? ~_GEN_1317 & ldq_17_bits_order_fail : ~_GEN_51 & ldq_17_bits_order_fail;
  wire        _GEN_24818 = dis_ld_val_1 ? ~_GEN_1318 & ldq_18_bits_order_fail : ~_GEN_52 & ldq_18_bits_order_fail;
  wire        _GEN_24819 = dis_ld_val_1 ? ~_GEN_1319 & ldq_19_bits_order_fail : ~_GEN_53 & ldq_19_bits_order_fail;
  wire        _GEN_24820 = dis_ld_val_1 ? ~_GEN_1320 & ldq_20_bits_order_fail : ~_GEN_54 & ldq_20_bits_order_fail;
  wire        _GEN_24821 = dis_ld_val_1 ? ~_GEN_1321 & ldq_21_bits_order_fail : ~_GEN_55 & ldq_21_bits_order_fail;
  wire        _GEN_24822 = dis_ld_val_1 ? ~_GEN_1322 & ldq_22_bits_order_fail : ~_GEN_56 & ldq_22_bits_order_fail;
  wire        _GEN_24823 = dis_ld_val_1 ? ~_GEN_1323 & ldq_23_bits_order_fail : ~_GEN_57 & ldq_23_bits_order_fail;
  wire        _GEN_24824 = dis_ld_val_1 ? ~_GEN_1324 & ldq_24_bits_order_fail : ~_GEN_58 & ldq_24_bits_order_fail;
  wire        _GEN_24825 = dis_ld_val_1 ? ~_GEN_1325 & ldq_25_bits_order_fail : ~_GEN_59 & ldq_25_bits_order_fail;
  wire        _GEN_24826 = dis_ld_val_1 ? ~_GEN_1326 & ldq_26_bits_order_fail : ~_GEN_60 & ldq_26_bits_order_fail;
  wire        _GEN_24827 = dis_ld_val_1 ? ~_GEN_1327 & ldq_27_bits_order_fail : ~_GEN_61 & ldq_27_bits_order_fail;
  wire        _GEN_24828 = dis_ld_val_1 ? ~_GEN_1328 & ldq_28_bits_order_fail : ~_GEN_62 & ldq_28_bits_order_fail;
  wire        _GEN_24829 = dis_ld_val_1 ? ~_GEN_1329 & ldq_29_bits_order_fail : ~_GEN_63 & ldq_29_bits_order_fail;
  wire        _GEN_24830 = dis_ld_val_1 ? ~_GEN_1330 & ldq_30_bits_order_fail : ~_GEN_64 & ldq_30_bits_order_fail;
  wire        _GEN_24831 = dis_ld_val_1 ? ~_GEN_1331 & ldq_31_bits_order_fail : ~_GEN_65 & ldq_31_bits_order_fail;
  wire        _GEN_24832 = dis_ld_val_1 ? ~_GEN_1300 & ldq_0_bits_observed : ~_GEN_34 & ldq_0_bits_observed;
  wire        _GEN_24833 = dis_ld_val_1 ? ~_GEN_1301 & ldq_1_bits_observed : ~_GEN_35 & ldq_1_bits_observed;
  wire        _GEN_24834 = dis_ld_val_1 ? ~_GEN_1302 & ldq_2_bits_observed : ~_GEN_36 & ldq_2_bits_observed;
  wire        _GEN_24835 = dis_ld_val_1 ? ~_GEN_1303 & ldq_3_bits_observed : ~_GEN_37 & ldq_3_bits_observed;
  wire        _GEN_24836 = dis_ld_val_1 ? ~_GEN_1304 & ldq_4_bits_observed : ~_GEN_38 & ldq_4_bits_observed;
  wire        _GEN_24837 = dis_ld_val_1 ? ~_GEN_1305 & ldq_5_bits_observed : ~_GEN_39 & ldq_5_bits_observed;
  wire        _GEN_24838 = dis_ld_val_1 ? ~_GEN_1306 & ldq_6_bits_observed : ~_GEN_40 & ldq_6_bits_observed;
  wire        _GEN_24839 = dis_ld_val_1 ? ~_GEN_1307 & ldq_7_bits_observed : ~_GEN_41 & ldq_7_bits_observed;
  wire        _GEN_24840 = dis_ld_val_1 ? ~_GEN_1308 & ldq_8_bits_observed : ~_GEN_42 & ldq_8_bits_observed;
  wire        _GEN_24841 = dis_ld_val_1 ? ~_GEN_1309 & ldq_9_bits_observed : ~_GEN_43 & ldq_9_bits_observed;
  wire        _GEN_24842 = dis_ld_val_1 ? ~_GEN_1310 & ldq_10_bits_observed : ~_GEN_44 & ldq_10_bits_observed;
  wire        _GEN_24843 = dis_ld_val_1 ? ~_GEN_1311 & ldq_11_bits_observed : ~_GEN_45 & ldq_11_bits_observed;
  wire        _GEN_24844 = dis_ld_val_1 ? ~_GEN_1312 & ldq_12_bits_observed : ~_GEN_46 & ldq_12_bits_observed;
  wire        _GEN_24845 = dis_ld_val_1 ? ~_GEN_1313 & ldq_13_bits_observed : ~_GEN_47 & ldq_13_bits_observed;
  wire        _GEN_24846 = dis_ld_val_1 ? ~_GEN_1314 & ldq_14_bits_observed : ~_GEN_48 & ldq_14_bits_observed;
  wire        _GEN_24847 = dis_ld_val_1 ? ~_GEN_1315 & ldq_15_bits_observed : ~_GEN_49 & ldq_15_bits_observed;
  wire        _GEN_24848 = dis_ld_val_1 ? ~_GEN_1316 & ldq_16_bits_observed : ~_GEN_50 & ldq_16_bits_observed;
  wire        _GEN_24849 = dis_ld_val_1 ? ~_GEN_1317 & ldq_17_bits_observed : ~_GEN_51 & ldq_17_bits_observed;
  wire        _GEN_24850 = dis_ld_val_1 ? ~_GEN_1318 & ldq_18_bits_observed : ~_GEN_52 & ldq_18_bits_observed;
  wire        _GEN_24851 = dis_ld_val_1 ? ~_GEN_1319 & ldq_19_bits_observed : ~_GEN_53 & ldq_19_bits_observed;
  wire        _GEN_24852 = dis_ld_val_1 ? ~_GEN_1320 & ldq_20_bits_observed : ~_GEN_54 & ldq_20_bits_observed;
  wire        _GEN_24853 = dis_ld_val_1 ? ~_GEN_1321 & ldq_21_bits_observed : ~_GEN_55 & ldq_21_bits_observed;
  wire        _GEN_24854 = dis_ld_val_1 ? ~_GEN_1322 & ldq_22_bits_observed : ~_GEN_56 & ldq_22_bits_observed;
  wire        _GEN_24855 = dis_ld_val_1 ? ~_GEN_1323 & ldq_23_bits_observed : ~_GEN_57 & ldq_23_bits_observed;
  wire        _GEN_24856 = dis_ld_val_1 ? ~_GEN_1324 & ldq_24_bits_observed : ~_GEN_58 & ldq_24_bits_observed;
  wire        _GEN_24857 = dis_ld_val_1 ? ~_GEN_1325 & ldq_25_bits_observed : ~_GEN_59 & ldq_25_bits_observed;
  wire        _GEN_24858 = dis_ld_val_1 ? ~_GEN_1326 & ldq_26_bits_observed : ~_GEN_60 & ldq_26_bits_observed;
  wire        _GEN_24859 = dis_ld_val_1 ? ~_GEN_1327 & ldq_27_bits_observed : ~_GEN_61 & ldq_27_bits_observed;
  wire        _GEN_24860 = dis_ld_val_1 ? ~_GEN_1328 & ldq_28_bits_observed : ~_GEN_62 & ldq_28_bits_observed;
  wire        _GEN_24861 = dis_ld_val_1 ? ~_GEN_1329 & ldq_29_bits_observed : ~_GEN_63 & ldq_29_bits_observed;
  wire        _GEN_24862 = dis_ld_val_1 ? ~_GEN_1330 & ldq_30_bits_observed : ~_GEN_64 & ldq_30_bits_observed;
  wire        _GEN_24863 = dis_ld_val_1 ? ~_GEN_1331 & ldq_31_bits_observed : ~_GEN_65 & ldq_31_bits_observed;
  wire        _GEN_24864 = dis_ld_val_1 ? ~_GEN_1300 & ldq_0_bits_forward_std_val : ~_GEN_34 & ldq_0_bits_forward_std_val;
  wire        _GEN_24865 = dis_ld_val_1 ? ~_GEN_1301 & ldq_1_bits_forward_std_val : ~_GEN_35 & ldq_1_bits_forward_std_val;
  wire        _GEN_24866 = dis_ld_val_1 ? ~_GEN_1302 & ldq_2_bits_forward_std_val : ~_GEN_36 & ldq_2_bits_forward_std_val;
  wire        _GEN_24867 = dis_ld_val_1 ? ~_GEN_1303 & ldq_3_bits_forward_std_val : ~_GEN_37 & ldq_3_bits_forward_std_val;
  wire        _GEN_24868 = dis_ld_val_1 ? ~_GEN_1304 & ldq_4_bits_forward_std_val : ~_GEN_38 & ldq_4_bits_forward_std_val;
  wire        _GEN_24869 = dis_ld_val_1 ? ~_GEN_1305 & ldq_5_bits_forward_std_val : ~_GEN_39 & ldq_5_bits_forward_std_val;
  wire        _GEN_24870 = dis_ld_val_1 ? ~_GEN_1306 & ldq_6_bits_forward_std_val : ~_GEN_40 & ldq_6_bits_forward_std_val;
  wire        _GEN_24871 = dis_ld_val_1 ? ~_GEN_1307 & ldq_7_bits_forward_std_val : ~_GEN_41 & ldq_7_bits_forward_std_val;
  wire        _GEN_24872 = dis_ld_val_1 ? ~_GEN_1308 & ldq_8_bits_forward_std_val : ~_GEN_42 & ldq_8_bits_forward_std_val;
  wire        _GEN_24873 = dis_ld_val_1 ? ~_GEN_1309 & ldq_9_bits_forward_std_val : ~_GEN_43 & ldq_9_bits_forward_std_val;
  wire        _GEN_24874 = dis_ld_val_1 ? ~_GEN_1310 & ldq_10_bits_forward_std_val : ~_GEN_44 & ldq_10_bits_forward_std_val;
  wire        _GEN_24875 = dis_ld_val_1 ? ~_GEN_1311 & ldq_11_bits_forward_std_val : ~_GEN_45 & ldq_11_bits_forward_std_val;
  wire        _GEN_24876 = dis_ld_val_1 ? ~_GEN_1312 & ldq_12_bits_forward_std_val : ~_GEN_46 & ldq_12_bits_forward_std_val;
  wire        _GEN_24877 = dis_ld_val_1 ? ~_GEN_1313 & ldq_13_bits_forward_std_val : ~_GEN_47 & ldq_13_bits_forward_std_val;
  wire        _GEN_24878 = dis_ld_val_1 ? ~_GEN_1314 & ldq_14_bits_forward_std_val : ~_GEN_48 & ldq_14_bits_forward_std_val;
  wire        _GEN_24879 = dis_ld_val_1 ? ~_GEN_1315 & ldq_15_bits_forward_std_val : ~_GEN_49 & ldq_15_bits_forward_std_val;
  wire        _GEN_24880 = dis_ld_val_1 ? ~_GEN_1316 & ldq_16_bits_forward_std_val : ~_GEN_50 & ldq_16_bits_forward_std_val;
  wire        _GEN_24881 = dis_ld_val_1 ? ~_GEN_1317 & ldq_17_bits_forward_std_val : ~_GEN_51 & ldq_17_bits_forward_std_val;
  wire        _GEN_24882 = dis_ld_val_1 ? ~_GEN_1318 & ldq_18_bits_forward_std_val : ~_GEN_52 & ldq_18_bits_forward_std_val;
  wire        _GEN_24883 = dis_ld_val_1 ? ~_GEN_1319 & ldq_19_bits_forward_std_val : ~_GEN_53 & ldq_19_bits_forward_std_val;
  wire        _GEN_24884 = dis_ld_val_1 ? ~_GEN_1320 & ldq_20_bits_forward_std_val : ~_GEN_54 & ldq_20_bits_forward_std_val;
  wire        _GEN_24885 = dis_ld_val_1 ? ~_GEN_1321 & ldq_21_bits_forward_std_val : ~_GEN_55 & ldq_21_bits_forward_std_val;
  wire        _GEN_24886 = dis_ld_val_1 ? ~_GEN_1322 & ldq_22_bits_forward_std_val : ~_GEN_56 & ldq_22_bits_forward_std_val;
  wire        _GEN_24887 = dis_ld_val_1 ? ~_GEN_1323 & ldq_23_bits_forward_std_val : ~_GEN_57 & ldq_23_bits_forward_std_val;
  wire        _GEN_24888 = dis_ld_val_1 ? ~_GEN_1324 & ldq_24_bits_forward_std_val : ~_GEN_58 & ldq_24_bits_forward_std_val;
  wire        _GEN_24889 = dis_ld_val_1 ? ~_GEN_1325 & ldq_25_bits_forward_std_val : ~_GEN_59 & ldq_25_bits_forward_std_val;
  wire        _GEN_24890 = dis_ld_val_1 ? ~_GEN_1326 & ldq_26_bits_forward_std_val : ~_GEN_60 & ldq_26_bits_forward_std_val;
  wire        _GEN_24891 = dis_ld_val_1 ? ~_GEN_1327 & ldq_27_bits_forward_std_val : ~_GEN_61 & ldq_27_bits_forward_std_val;
  wire        _GEN_24892 = dis_ld_val_1 ? ~_GEN_1328 & ldq_28_bits_forward_std_val : ~_GEN_62 & ldq_28_bits_forward_std_val;
  wire        _GEN_24893 = dis_ld_val_1 ? ~_GEN_1329 & ldq_29_bits_forward_std_val : ~_GEN_63 & ldq_29_bits_forward_std_val;
  wire        _GEN_24894 = dis_ld_val_1 ? ~_GEN_1330 & ldq_30_bits_forward_std_val : ~_GEN_64 & ldq_30_bits_forward_std_val;
  wire        _GEN_24895 = dis_ld_val_1 ? ~_GEN_1331 & ldq_31_bits_forward_std_val : ~_GEN_65 & ldq_31_bits_forward_std_val;
  wire        _GEN_1332 = dis_ld_val_1 | ~_GEN_100;
  wire        _GEN_1333 = dis_ld_val_1 | ~_GEN_101;
  wire        _GEN_1334 = dis_ld_val_1 | ~_GEN_102;
  wire        _GEN_1335 = dis_ld_val_1 | ~_GEN_103;
  wire        _GEN_1336 = dis_ld_val_1 | ~_GEN_104;
  wire        _GEN_1337 = dis_ld_val_1 | ~_GEN_105;
  wire        _GEN_1338 = dis_ld_val_1 | ~_GEN_106;
  wire        _GEN_1339 = dis_ld_val_1 | ~_GEN_107;
  wire        _GEN_1340 = dis_ld_val_1 | ~_GEN_108;
  wire        _GEN_1341 = dis_ld_val_1 | ~_GEN_109;
  wire        _GEN_1342 = dis_ld_val_1 | ~_GEN_110;
  wire        _GEN_1343 = dis_ld_val_1 | ~_GEN_111;
  wire        _GEN_1344 = dis_ld_val_1 | ~_GEN_112;
  wire        _GEN_1345 = dis_ld_val_1 | ~_GEN_113;
  wire        _GEN_1346 = dis_ld_val_1 | ~_GEN_114;
  wire        _GEN_1347 = dis_ld_val_1 | ~_GEN_115;
  wire        _GEN_1348 = dis_ld_val_1 | ~_GEN_116;
  wire        _GEN_1349 = dis_ld_val_1 | ~_GEN_117;
  wire        _GEN_1350 = dis_ld_val_1 | ~_GEN_118;
  wire        _GEN_1351 = dis_ld_val_1 | ~_GEN_119;
  wire        _GEN_1352 = dis_ld_val_1 | ~_GEN_120;
  wire        _GEN_1353 = dis_ld_val_1 | ~_GEN_121;
  wire        _GEN_1354 = dis_ld_val_1 | ~_GEN_122;
  wire        _GEN_1355 = dis_ld_val_1 | ~_GEN_123;
  wire        _GEN_1356 = dis_ld_val_1 | ~_GEN_124;
  wire        _GEN_1357 = dis_ld_val_1 | ~_GEN_125;
  wire        _GEN_1358 = dis_ld_val_1 | ~_GEN_126;
  wire        _GEN_1359 = dis_ld_val_1 | ~_GEN_127;
  wire        _GEN_1360 = dis_ld_val_1 | ~_GEN_128;
  wire        _GEN_1361 = dis_ld_val_1 | ~_GEN_129;
  wire        _GEN_1362 = dis_ld_val_1 | ~_GEN_130;
  wire        _GEN_1363 = dis_ld_val_1 | ~_GEN_131;
  wire [31:0] _ldq_T_75_bits_st_dep_mask = {32{dis_st_val_1}} & 32'h1 << _ldq_T_35_bits_youngest_stq_idx | _ldq_T_35_bits_st_dep_mask;
  wire        _GEN_1364 = dis_ld_val_2 | ~_GEN_167;
  wire        _GEN_1365 = dis_ld_val_2 | ~_GEN_168;
  wire        _GEN_1366 = dis_ld_val_2 | ~_GEN_169;
  wire        _GEN_1367 = dis_ld_val_2 | ~_GEN_170;
  wire        _GEN_1368 = dis_ld_val_2 | ~_GEN_171;
  wire        _GEN_1369 = dis_ld_val_2 | ~_GEN_172;
  wire        _GEN_1370 = dis_ld_val_2 | ~_GEN_173;
  wire        _GEN_1371 = dis_ld_val_2 | ~_GEN_174;
  wire        _GEN_1372 = dis_ld_val_2 | ~_GEN_175;
  wire        _GEN_1373 = dis_ld_val_2 | ~_GEN_176;
  wire        _GEN_1374 = dis_ld_val_2 | ~_GEN_177;
  wire        _GEN_1375 = dis_ld_val_2 | ~_GEN_178;
  wire        _GEN_1376 = dis_ld_val_2 | ~_GEN_179;
  wire        _GEN_1377 = dis_ld_val_2 | ~_GEN_180;
  wire        _GEN_1378 = dis_ld_val_2 | ~_GEN_181;
  wire        _GEN_1379 = dis_ld_val_2 | ~_GEN_182;
  wire        _GEN_1380 = dis_ld_val_2 | ~_GEN_183;
  wire        _GEN_1381 = dis_ld_val_2 | ~_GEN_184;
  wire        _GEN_1382 = dis_ld_val_2 | ~_GEN_185;
  wire        _GEN_1383 = dis_ld_val_2 | ~_GEN_186;
  wire        _GEN_1384 = dis_ld_val_2 | ~_GEN_187;
  wire        _GEN_1385 = dis_ld_val_2 | ~_GEN_188;
  wire        _GEN_1386 = dis_ld_val_2 | ~_GEN_189;
  wire        _GEN_1387 = dis_ld_val_2 | ~_GEN_190;
  wire        _GEN_1388 = dis_ld_val_2 | ~_GEN_191;
  wire        _GEN_1389 = dis_ld_val_2 | ~_GEN_192;
  wire        _GEN_1390 = dis_ld_val_2 | ~_GEN_193;
  wire        _GEN_1391 = dis_ld_val_2 | ~_GEN_194;
  wire        _GEN_1392 = dis_ld_val_2 | ~_GEN_195;
  wire        _GEN_1393 = dis_ld_val_2 | ~_GEN_196;
  wire        _GEN_1394 = dis_ld_val_2 | ~_GEN_197;
  wire        _GEN_1395 = dis_ld_val_2 | ~_GEN_198;
  wire [31:0] _ldq_T_115_bits_st_dep_mask = {32{dis_st_val_2}} & 32'h1 << _ldq_T_75_bits_youngest_stq_idx | _ldq_T_75_bits_st_dep_mask;
  wire        _GEN_1396 = _GEN_234 | _GEN_199;
  wire        _GEN_1397 = _GEN_235 | _GEN_200;
  wire        _GEN_1398 = _GEN_236 | _GEN_201;
  wire        _GEN_1399 = _GEN_237 | _GEN_202;
  wire        _GEN_1400 = _GEN_238 | _GEN_203;
  wire        _GEN_1401 = _GEN_239 | _GEN_204;
  wire        _GEN_1402 = _GEN_240 | _GEN_205;
  wire        _GEN_1403 = _GEN_241 | _GEN_206;
  wire        _GEN_1404 = _GEN_242 | _GEN_207;
  wire        _GEN_1405 = _GEN_243 | _GEN_208;
  wire        _GEN_1406 = _GEN_244 | _GEN_209;
  wire        _GEN_1407 = _GEN_245 | _GEN_210;
  wire        _GEN_1408 = _GEN_246 | _GEN_211;
  wire        _GEN_1409 = _GEN_247 | _GEN_212;
  wire        _GEN_1410 = _GEN_248 | _GEN_213;
  wire        _GEN_1411 = _GEN_249 | _GEN_214;
  wire        _GEN_1412 = _GEN_250 | _GEN_215;
  wire        _GEN_1413 = _GEN_251 | _GEN_216;
  wire        _GEN_1414 = _GEN_252 | _GEN_217;
  wire        _GEN_1415 = _GEN_253 | _GEN_218;
  wire        _GEN_1416 = _GEN_254 | _GEN_219;
  wire        _GEN_1417 = _GEN_255 | _GEN_220;
  wire        _GEN_1418 = _GEN_256 | _GEN_221;
  wire        _GEN_1419 = _GEN_257 | _GEN_222;
  wire        _GEN_1420 = _GEN_258 | _GEN_223;
  wire        _GEN_1421 = _GEN_259 | _GEN_224;
  wire        _GEN_1422 = _GEN_260 | _GEN_225;
  wire        _GEN_1423 = _GEN_261 | _GEN_226;
  wire        _GEN_1424 = _GEN_262 | _GEN_227;
  wire        _GEN_1425 = _GEN_263 | _GEN_228;
  wire        _GEN_1426 = _GEN_264 | _GEN_229;
  wire        _GEN_1427 = (&_GEN_231) | _GEN_230;
  wire        _GEN_49600 = dis_ld_val_3 ? _GEN_1396 | _GEN_22080 : _GEN_199 | _GEN_22080;
  wire        _GEN_49601 = dis_ld_val_3 ? _GEN_1397 | _GEN_22081 : _GEN_200 | _GEN_22081;
  wire        _GEN_49602 = dis_ld_val_3 ? _GEN_1398 | _GEN_22082 : _GEN_201 | _GEN_22082;
  wire        _GEN_49603 = dis_ld_val_3 ? _GEN_1399 | _GEN_22083 : _GEN_202 | _GEN_22083;
  wire        _GEN_49604 = dis_ld_val_3 ? _GEN_1400 | _GEN_22084 : _GEN_203 | _GEN_22084;
  wire        _GEN_49605 = dis_ld_val_3 ? _GEN_1401 | _GEN_22085 : _GEN_204 | _GEN_22085;
  wire        _GEN_49606 = dis_ld_val_3 ? _GEN_1402 | _GEN_22086 : _GEN_205 | _GEN_22086;
  wire        _GEN_49607 = dis_ld_val_3 ? _GEN_1403 | _GEN_22087 : _GEN_206 | _GEN_22087;
  wire        _GEN_49608 = dis_ld_val_3 ? _GEN_1404 | _GEN_22088 : _GEN_207 | _GEN_22088;
  wire        _GEN_49609 = dis_ld_val_3 ? _GEN_1405 | _GEN_22089 : _GEN_208 | _GEN_22089;
  wire        _GEN_49610 = dis_ld_val_3 ? _GEN_1406 | _GEN_22090 : _GEN_209 | _GEN_22090;
  wire        _GEN_49611 = dis_ld_val_3 ? _GEN_1407 | _GEN_22091 : _GEN_210 | _GEN_22091;
  wire        _GEN_49612 = dis_ld_val_3 ? _GEN_1408 | _GEN_22092 : _GEN_211 | _GEN_22092;
  wire        _GEN_49613 = dis_ld_val_3 ? _GEN_1409 | _GEN_22093 : _GEN_212 | _GEN_22093;
  wire        _GEN_49614 = dis_ld_val_3 ? _GEN_1410 | _GEN_22094 : _GEN_213 | _GEN_22094;
  wire        _GEN_49615 = dis_ld_val_3 ? _GEN_1411 | _GEN_22095 : _GEN_214 | _GEN_22095;
  wire        _GEN_49616 = dis_ld_val_3 ? _GEN_1412 | _GEN_22096 : _GEN_215 | _GEN_22096;
  wire        _GEN_49617 = dis_ld_val_3 ? _GEN_1413 | _GEN_22097 : _GEN_216 | _GEN_22097;
  wire        _GEN_49618 = dis_ld_val_3 ? _GEN_1414 | _GEN_22098 : _GEN_217 | _GEN_22098;
  wire        _GEN_49619 = dis_ld_val_3 ? _GEN_1415 | _GEN_22099 : _GEN_218 | _GEN_22099;
  wire        _GEN_49620 = dis_ld_val_3 ? _GEN_1416 | _GEN_22100 : _GEN_219 | _GEN_22100;
  wire        _GEN_49621 = dis_ld_val_3 ? _GEN_1417 | _GEN_22101 : _GEN_220 | _GEN_22101;
  wire        _GEN_49622 = dis_ld_val_3 ? _GEN_1418 | _GEN_22102 : _GEN_221 | _GEN_22102;
  wire        _GEN_49623 = dis_ld_val_3 ? _GEN_1419 | _GEN_22103 : _GEN_222 | _GEN_22103;
  wire        _GEN_49624 = dis_ld_val_3 ? _GEN_1420 | _GEN_22104 : _GEN_223 | _GEN_22104;
  wire        _GEN_49625 = dis_ld_val_3 ? _GEN_1421 | _GEN_22105 : _GEN_224 | _GEN_22105;
  wire        _GEN_49626 = dis_ld_val_3 ? _GEN_1422 | _GEN_22106 : _GEN_225 | _GEN_22106;
  wire        _GEN_49627 = dis_ld_val_3 ? _GEN_1423 | _GEN_22107 : _GEN_226 | _GEN_22107;
  wire        _GEN_49628 = dis_ld_val_3 ? _GEN_1424 | _GEN_22108 : _GEN_227 | _GEN_22108;
  wire        _GEN_49629 = dis_ld_val_3 ? _GEN_1425 | _GEN_22109 : _GEN_228 | _GEN_22109;
  wire        _GEN_49630 = dis_ld_val_3 ? _GEN_1426 | _GEN_22110 : _GEN_229 | _GEN_22110;
  wire        _GEN_49631 = dis_ld_val_3 ? _GEN_1427 | _GEN_22111 : _GEN_230 | _GEN_22111;
  wire        _GEN_52224 = dis_ld_val_3 ? ~_GEN_1396 & _GEN_24704 : ~_GEN_199 & _GEN_24704;
  wire        _GEN_52225 = dis_ld_val_3 ? ~_GEN_1397 & _GEN_24705 : ~_GEN_200 & _GEN_24705;
  wire        _GEN_52226 = dis_ld_val_3 ? ~_GEN_1398 & _GEN_24706 : ~_GEN_201 & _GEN_24706;
  wire        _GEN_52227 = dis_ld_val_3 ? ~_GEN_1399 & _GEN_24707 : ~_GEN_202 & _GEN_24707;
  wire        _GEN_52228 = dis_ld_val_3 ? ~_GEN_1400 & _GEN_24708 : ~_GEN_203 & _GEN_24708;
  wire        _GEN_52229 = dis_ld_val_3 ? ~_GEN_1401 & _GEN_24709 : ~_GEN_204 & _GEN_24709;
  wire        _GEN_52230 = dis_ld_val_3 ? ~_GEN_1402 & _GEN_24710 : ~_GEN_205 & _GEN_24710;
  wire        _GEN_52231 = dis_ld_val_3 ? ~_GEN_1403 & _GEN_24711 : ~_GEN_206 & _GEN_24711;
  wire        _GEN_52232 = dis_ld_val_3 ? ~_GEN_1404 & _GEN_24712 : ~_GEN_207 & _GEN_24712;
  wire        _GEN_52233 = dis_ld_val_3 ? ~_GEN_1405 & _GEN_24713 : ~_GEN_208 & _GEN_24713;
  wire        _GEN_52234 = dis_ld_val_3 ? ~_GEN_1406 & _GEN_24714 : ~_GEN_209 & _GEN_24714;
  wire        _GEN_52235 = dis_ld_val_3 ? ~_GEN_1407 & _GEN_24715 : ~_GEN_210 & _GEN_24715;
  wire        _GEN_52236 = dis_ld_val_3 ? ~_GEN_1408 & _GEN_24716 : ~_GEN_211 & _GEN_24716;
  wire        _GEN_52237 = dis_ld_val_3 ? ~_GEN_1409 & _GEN_24717 : ~_GEN_212 & _GEN_24717;
  wire        _GEN_52238 = dis_ld_val_3 ? ~_GEN_1410 & _GEN_24718 : ~_GEN_213 & _GEN_24718;
  wire        _GEN_52239 = dis_ld_val_3 ? ~_GEN_1411 & _GEN_24719 : ~_GEN_214 & _GEN_24719;
  wire        _GEN_52240 = dis_ld_val_3 ? ~_GEN_1412 & _GEN_24720 : ~_GEN_215 & _GEN_24720;
  wire        _GEN_52241 = dis_ld_val_3 ? ~_GEN_1413 & _GEN_24721 : ~_GEN_216 & _GEN_24721;
  wire        _GEN_52242 = dis_ld_val_3 ? ~_GEN_1414 & _GEN_24722 : ~_GEN_217 & _GEN_24722;
  wire        _GEN_52243 = dis_ld_val_3 ? ~_GEN_1415 & _GEN_24723 : ~_GEN_218 & _GEN_24723;
  wire        _GEN_52244 = dis_ld_val_3 ? ~_GEN_1416 & _GEN_24724 : ~_GEN_219 & _GEN_24724;
  wire        _GEN_52245 = dis_ld_val_3 ? ~_GEN_1417 & _GEN_24725 : ~_GEN_220 & _GEN_24725;
  wire        _GEN_52246 = dis_ld_val_3 ? ~_GEN_1418 & _GEN_24726 : ~_GEN_221 & _GEN_24726;
  wire        _GEN_52247 = dis_ld_val_3 ? ~_GEN_1419 & _GEN_24727 : ~_GEN_222 & _GEN_24727;
  wire        _GEN_52248 = dis_ld_val_3 ? ~_GEN_1420 & _GEN_24728 : ~_GEN_223 & _GEN_24728;
  wire        _GEN_52249 = dis_ld_val_3 ? ~_GEN_1421 & _GEN_24729 : ~_GEN_224 & _GEN_24729;
  wire        _GEN_52250 = dis_ld_val_3 ? ~_GEN_1422 & _GEN_24730 : ~_GEN_225 & _GEN_24730;
  wire        _GEN_52251 = dis_ld_val_3 ? ~_GEN_1423 & _GEN_24731 : ~_GEN_226 & _GEN_24731;
  wire        _GEN_52252 = dis_ld_val_3 ? ~_GEN_1424 & _GEN_24732 : ~_GEN_227 & _GEN_24732;
  wire        _GEN_52253 = dis_ld_val_3 ? ~_GEN_1425 & _GEN_24733 : ~_GEN_228 & _GEN_24733;
  wire        _GEN_52254 = dis_ld_val_3 ? ~_GEN_1426 & _GEN_24734 : ~_GEN_229 & _GEN_24734;
  wire        _GEN_52255 = dis_ld_val_3 ? ~_GEN_1427 & _GEN_24735 : ~_GEN_230 & _GEN_24735;
  wire        _GEN_52320 = dis_ld_val_3 ? ~_GEN_1396 & _GEN_24800 : ~_GEN_199 & _GEN_24800;
  wire        _GEN_52321 = dis_ld_val_3 ? ~_GEN_1397 & _GEN_24801 : ~_GEN_200 & _GEN_24801;
  wire        _GEN_52322 = dis_ld_val_3 ? ~_GEN_1398 & _GEN_24802 : ~_GEN_201 & _GEN_24802;
  wire        _GEN_52323 = dis_ld_val_3 ? ~_GEN_1399 & _GEN_24803 : ~_GEN_202 & _GEN_24803;
  wire        _GEN_52324 = dis_ld_val_3 ? ~_GEN_1400 & _GEN_24804 : ~_GEN_203 & _GEN_24804;
  wire        _GEN_52325 = dis_ld_val_3 ? ~_GEN_1401 & _GEN_24805 : ~_GEN_204 & _GEN_24805;
  wire        _GEN_52326 = dis_ld_val_3 ? ~_GEN_1402 & _GEN_24806 : ~_GEN_205 & _GEN_24806;
  wire        _GEN_52327 = dis_ld_val_3 ? ~_GEN_1403 & _GEN_24807 : ~_GEN_206 & _GEN_24807;
  wire        _GEN_52328 = dis_ld_val_3 ? ~_GEN_1404 & _GEN_24808 : ~_GEN_207 & _GEN_24808;
  wire        _GEN_52329 = dis_ld_val_3 ? ~_GEN_1405 & _GEN_24809 : ~_GEN_208 & _GEN_24809;
  wire        _GEN_52330 = dis_ld_val_3 ? ~_GEN_1406 & _GEN_24810 : ~_GEN_209 & _GEN_24810;
  wire        _GEN_52331 = dis_ld_val_3 ? ~_GEN_1407 & _GEN_24811 : ~_GEN_210 & _GEN_24811;
  wire        _GEN_52332 = dis_ld_val_3 ? ~_GEN_1408 & _GEN_24812 : ~_GEN_211 & _GEN_24812;
  wire        _GEN_52333 = dis_ld_val_3 ? ~_GEN_1409 & _GEN_24813 : ~_GEN_212 & _GEN_24813;
  wire        _GEN_52334 = dis_ld_val_3 ? ~_GEN_1410 & _GEN_24814 : ~_GEN_213 & _GEN_24814;
  wire        _GEN_52335 = dis_ld_val_3 ? ~_GEN_1411 & _GEN_24815 : ~_GEN_214 & _GEN_24815;
  wire        _GEN_52336 = dis_ld_val_3 ? ~_GEN_1412 & _GEN_24816 : ~_GEN_215 & _GEN_24816;
  wire        _GEN_52337 = dis_ld_val_3 ? ~_GEN_1413 & _GEN_24817 : ~_GEN_216 & _GEN_24817;
  wire        _GEN_52338 = dis_ld_val_3 ? ~_GEN_1414 & _GEN_24818 : ~_GEN_217 & _GEN_24818;
  wire        _GEN_52339 = dis_ld_val_3 ? ~_GEN_1415 & _GEN_24819 : ~_GEN_218 & _GEN_24819;
  wire        _GEN_52340 = dis_ld_val_3 ? ~_GEN_1416 & _GEN_24820 : ~_GEN_219 & _GEN_24820;
  wire        _GEN_52341 = dis_ld_val_3 ? ~_GEN_1417 & _GEN_24821 : ~_GEN_220 & _GEN_24821;
  wire        _GEN_52342 = dis_ld_val_3 ? ~_GEN_1418 & _GEN_24822 : ~_GEN_221 & _GEN_24822;
  wire        _GEN_52343 = dis_ld_val_3 ? ~_GEN_1419 & _GEN_24823 : ~_GEN_222 & _GEN_24823;
  wire        _GEN_52344 = dis_ld_val_3 ? ~_GEN_1420 & _GEN_24824 : ~_GEN_223 & _GEN_24824;
  wire        _GEN_52345 = dis_ld_val_3 ? ~_GEN_1421 & _GEN_24825 : ~_GEN_224 & _GEN_24825;
  wire        _GEN_52346 = dis_ld_val_3 ? ~_GEN_1422 & _GEN_24826 : ~_GEN_225 & _GEN_24826;
  wire        _GEN_52347 = dis_ld_val_3 ? ~_GEN_1423 & _GEN_24827 : ~_GEN_226 & _GEN_24827;
  wire        _GEN_52348 = dis_ld_val_3 ? ~_GEN_1424 & _GEN_24828 : ~_GEN_227 & _GEN_24828;
  wire        _GEN_52349 = dis_ld_val_3 ? ~_GEN_1425 & _GEN_24829 : ~_GEN_228 & _GEN_24829;
  wire        _GEN_52350 = dis_ld_val_3 ? ~_GEN_1426 & _GEN_24830 : ~_GEN_229 & _GEN_24830;
  wire        _GEN_52351 = dis_ld_val_3 ? ~_GEN_1427 & _GEN_24831 : ~_GEN_230 & _GEN_24831;
  wire        _GEN_52416 = ~dis_ld_val_3 & _GEN_265 | ~dis_ld_val_2 & _GEN_167 | ~dis_ld_val_1 & _GEN_100 | ~dis_ld_val & _GEN_2 | stq_0_valid;
  wire        _GEN_52417 = ~dis_ld_val_3 & _GEN_266 | ~dis_ld_val_2 & _GEN_168 | ~dis_ld_val_1 & _GEN_101 | ~dis_ld_val & _GEN_3 | stq_1_valid;
  wire        _GEN_52418 = ~dis_ld_val_3 & _GEN_267 | ~dis_ld_val_2 & _GEN_169 | ~dis_ld_val_1 & _GEN_102 | ~dis_ld_val & _GEN_4 | stq_2_valid;
  wire        _GEN_52419 = ~dis_ld_val_3 & _GEN_268 | ~dis_ld_val_2 & _GEN_170 | ~dis_ld_val_1 & _GEN_103 | ~dis_ld_val & _GEN_5 | stq_3_valid;
  wire        _GEN_52420 = ~dis_ld_val_3 & _GEN_269 | ~dis_ld_val_2 & _GEN_171 | ~dis_ld_val_1 & _GEN_104 | ~dis_ld_val & _GEN_6 | stq_4_valid;
  wire        _GEN_52421 = ~dis_ld_val_3 & _GEN_270 | ~dis_ld_val_2 & _GEN_172 | ~dis_ld_val_1 & _GEN_105 | ~dis_ld_val & _GEN_7 | stq_5_valid;
  wire        _GEN_52422 = ~dis_ld_val_3 & _GEN_271 | ~dis_ld_val_2 & _GEN_173 | ~dis_ld_val_1 & _GEN_106 | ~dis_ld_val & _GEN_8 | stq_6_valid;
  wire        _GEN_52423 = ~dis_ld_val_3 & _GEN_272 | ~dis_ld_val_2 & _GEN_174 | ~dis_ld_val_1 & _GEN_107 | ~dis_ld_val & _GEN_9 | stq_7_valid;
  wire        _GEN_52424 = ~dis_ld_val_3 & _GEN_273 | ~dis_ld_val_2 & _GEN_175 | ~dis_ld_val_1 & _GEN_108 | ~dis_ld_val & _GEN_10 | stq_8_valid;
  wire        _GEN_52425 = ~dis_ld_val_3 & _GEN_274 | ~dis_ld_val_2 & _GEN_176 | ~dis_ld_val_1 & _GEN_109 | ~dis_ld_val & _GEN_11 | stq_9_valid;
  wire        _GEN_52426 = ~dis_ld_val_3 & _GEN_275 | ~dis_ld_val_2 & _GEN_177 | ~dis_ld_val_1 & _GEN_110 | ~dis_ld_val & _GEN_12 | stq_10_valid;
  wire        _GEN_52427 = ~dis_ld_val_3 & _GEN_276 | ~dis_ld_val_2 & _GEN_178 | ~dis_ld_val_1 & _GEN_111 | ~dis_ld_val & _GEN_13 | stq_11_valid;
  wire        _GEN_52428 = ~dis_ld_val_3 & _GEN_277 | ~dis_ld_val_2 & _GEN_179 | ~dis_ld_val_1 & _GEN_112 | ~dis_ld_val & _GEN_14 | stq_12_valid;
  wire        _GEN_52429 = ~dis_ld_val_3 & _GEN_278 | ~dis_ld_val_2 & _GEN_180 | ~dis_ld_val_1 & _GEN_113 | ~dis_ld_val & _GEN_15 | stq_13_valid;
  wire        _GEN_52430 = ~dis_ld_val_3 & _GEN_279 | ~dis_ld_val_2 & _GEN_181 | ~dis_ld_val_1 & _GEN_114 | ~dis_ld_val & _GEN_16 | stq_14_valid;
  wire        _GEN_52431 = ~dis_ld_val_3 & _GEN_280 | ~dis_ld_val_2 & _GEN_182 | ~dis_ld_val_1 & _GEN_115 | ~dis_ld_val & _GEN_17 | stq_15_valid;
  wire        _GEN_52432 = ~dis_ld_val_3 & _GEN_281 | ~dis_ld_val_2 & _GEN_183 | ~dis_ld_val_1 & _GEN_116 | ~dis_ld_val & _GEN_18 | stq_16_valid;
  wire        _GEN_52433 = ~dis_ld_val_3 & _GEN_282 | ~dis_ld_val_2 & _GEN_184 | ~dis_ld_val_1 & _GEN_117 | ~dis_ld_val & _GEN_19 | stq_17_valid;
  wire        _GEN_52434 = ~dis_ld_val_3 & _GEN_283 | ~dis_ld_val_2 & _GEN_185 | ~dis_ld_val_1 & _GEN_118 | ~dis_ld_val & _GEN_20 | stq_18_valid;
  wire        _GEN_52435 = ~dis_ld_val_3 & _GEN_284 | ~dis_ld_val_2 & _GEN_186 | ~dis_ld_val_1 & _GEN_119 | ~dis_ld_val & _GEN_21 | stq_19_valid;
  wire        _GEN_52436 = ~dis_ld_val_3 & _GEN_285 | ~dis_ld_val_2 & _GEN_187 | ~dis_ld_val_1 & _GEN_120 | ~dis_ld_val & _GEN_22 | stq_20_valid;
  wire        _GEN_52437 = ~dis_ld_val_3 & _GEN_286 | ~dis_ld_val_2 & _GEN_188 | ~dis_ld_val_1 & _GEN_121 | ~dis_ld_val & _GEN_23 | stq_21_valid;
  wire        _GEN_52438 = ~dis_ld_val_3 & _GEN_287 | ~dis_ld_val_2 & _GEN_189 | ~dis_ld_val_1 & _GEN_122 | ~dis_ld_val & _GEN_24 | stq_22_valid;
  wire        _GEN_52439 = ~dis_ld_val_3 & _GEN_288 | ~dis_ld_val_2 & _GEN_190 | ~dis_ld_val_1 & _GEN_123 | ~dis_ld_val & _GEN_25 | stq_23_valid;
  wire        _GEN_52440 = ~dis_ld_val_3 & _GEN_289 | ~dis_ld_val_2 & _GEN_191 | ~dis_ld_val_1 & _GEN_124 | ~dis_ld_val & _GEN_26 | stq_24_valid;
  wire        _GEN_52441 = ~dis_ld_val_3 & _GEN_290 | ~dis_ld_val_2 & _GEN_192 | ~dis_ld_val_1 & _GEN_125 | ~dis_ld_val & _GEN_27 | stq_25_valid;
  wire        _GEN_52442 = ~dis_ld_val_3 & _GEN_291 | ~dis_ld_val_2 & _GEN_193 | ~dis_ld_val_1 & _GEN_126 | ~dis_ld_val & _GEN_28 | stq_26_valid;
  wire        _GEN_52443 = ~dis_ld_val_3 & _GEN_292 | ~dis_ld_val_2 & _GEN_194 | ~dis_ld_val_1 & _GEN_127 | ~dis_ld_val & _GEN_29 | stq_27_valid;
  wire        _GEN_52444 = ~dis_ld_val_3 & _GEN_293 | ~dis_ld_val_2 & _GEN_195 | ~dis_ld_val_1 & _GEN_128 | ~dis_ld_val & _GEN_30 | stq_28_valid;
  wire        _GEN_52445 = ~dis_ld_val_3 & _GEN_294 | ~dis_ld_val_2 & _GEN_196 | ~dis_ld_val_1 & _GEN_129 | ~dis_ld_val & _GEN_31 | stq_29_valid;
  wire        _GEN_52446 = ~dis_ld_val_3 & _GEN_295 | ~dis_ld_val_2 & _GEN_197 | ~dis_ld_val_1 & _GEN_130 | ~dis_ld_val & _GEN_32 | stq_30_valid;
  wire        _GEN_52447 = ~dis_ld_val_3 & _GEN_296 | ~dis_ld_val_2 & _GEN_198 | ~dis_ld_val_1 & _GEN_131 | ~dis_ld_val & _GEN_33 | stq_31_valid;
  wire        _GEN_1428 = dis_ld_val_3 | ~_GEN_265;
  wire        _GEN_1429 = dis_ld_val_3 | ~_GEN_266;
  wire        _GEN_1430 = dis_ld_val_3 | ~_GEN_267;
  wire        _GEN_1431 = dis_ld_val_3 | ~_GEN_268;
  wire        _GEN_1432 = dis_ld_val_3 | ~_GEN_269;
  wire        _GEN_1433 = dis_ld_val_3 | ~_GEN_270;
  wire        _GEN_1434 = dis_ld_val_3 | ~_GEN_271;
  wire        _GEN_1435 = dis_ld_val_3 | ~_GEN_272;
  wire        _GEN_1436 = dis_ld_val_3 | ~_GEN_273;
  wire        _GEN_1437 = dis_ld_val_3 | ~_GEN_274;
  wire        _GEN_1438 = dis_ld_val_3 | ~_GEN_275;
  wire        _GEN_1439 = dis_ld_val_3 | ~_GEN_276;
  wire        _GEN_1440 = dis_ld_val_3 | ~_GEN_277;
  wire        _GEN_1441 = dis_ld_val_3 | ~_GEN_278;
  wire        _GEN_1442 = dis_ld_val_3 | ~_GEN_279;
  wire        _GEN_1443 = dis_ld_val_3 | ~_GEN_280;
  wire        _GEN_1444 = dis_ld_val_3 | ~_GEN_281;
  wire        _GEN_1445 = dis_ld_val_3 | ~_GEN_282;
  wire        _GEN_1446 = dis_ld_val_3 | ~_GEN_283;
  wire        _GEN_1447 = dis_ld_val_3 | ~_GEN_284;
  wire        _GEN_1448 = dis_ld_val_3 | ~_GEN_285;
  wire        _GEN_1449 = dis_ld_val_3 | ~_GEN_286;
  wire        _GEN_1450 = dis_ld_val_3 | ~_GEN_287;
  wire        _GEN_1451 = dis_ld_val_3 | ~_GEN_288;
  wire        _GEN_1452 = dis_ld_val_3 | ~_GEN_289;
  wire        _GEN_1453 = dis_ld_val_3 | ~_GEN_290;
  wire        _GEN_1454 = dis_ld_val_3 | ~_GEN_291;
  wire        _GEN_1455 = dis_ld_val_3 | ~_GEN_292;
  wire        _GEN_1456 = dis_ld_val_3 | ~_GEN_293;
  wire        _GEN_1457 = dis_ld_val_3 | ~_GEN_294;
  wire        _GEN_1458 = dis_ld_val_3 | ~_GEN_295;
  wire        _GEN_1459 = dis_ld_val_3 | ~_GEN_296;
  wire        _GEN_55008 = _GEN_1428 & _GEN_1364 & _GEN_1332 & _GEN_1268 & stq_0_bits_data_valid;
  wire        _GEN_55009 = _GEN_1429 & _GEN_1365 & _GEN_1333 & _GEN_1269 & stq_1_bits_data_valid;
  wire        _GEN_55010 = _GEN_1430 & _GEN_1366 & _GEN_1334 & _GEN_1270 & stq_2_bits_data_valid;
  wire        _GEN_55011 = _GEN_1431 & _GEN_1367 & _GEN_1335 & _GEN_1271 & stq_3_bits_data_valid;
  wire        _GEN_55012 = _GEN_1432 & _GEN_1368 & _GEN_1336 & _GEN_1272 & stq_4_bits_data_valid;
  wire        _GEN_55013 = _GEN_1433 & _GEN_1369 & _GEN_1337 & _GEN_1273 & stq_5_bits_data_valid;
  wire        _GEN_55014 = _GEN_1434 & _GEN_1370 & _GEN_1338 & _GEN_1274 & stq_6_bits_data_valid;
  wire        _GEN_55015 = _GEN_1435 & _GEN_1371 & _GEN_1339 & _GEN_1275 & stq_7_bits_data_valid;
  wire        _GEN_55016 = _GEN_1436 & _GEN_1372 & _GEN_1340 & _GEN_1276 & stq_8_bits_data_valid;
  wire        _GEN_55017 = _GEN_1437 & _GEN_1373 & _GEN_1341 & _GEN_1277 & stq_9_bits_data_valid;
  wire        _GEN_55018 = _GEN_1438 & _GEN_1374 & _GEN_1342 & _GEN_1278 & stq_10_bits_data_valid;
  wire        _GEN_55019 = _GEN_1439 & _GEN_1375 & _GEN_1343 & _GEN_1279 & stq_11_bits_data_valid;
  wire        _GEN_55020 = _GEN_1440 & _GEN_1376 & _GEN_1344 & _GEN_1280 & stq_12_bits_data_valid;
  wire        _GEN_55021 = _GEN_1441 & _GEN_1377 & _GEN_1345 & _GEN_1281 & stq_13_bits_data_valid;
  wire        _GEN_55022 = _GEN_1442 & _GEN_1378 & _GEN_1346 & _GEN_1282 & stq_14_bits_data_valid;
  wire        _GEN_55023 = _GEN_1443 & _GEN_1379 & _GEN_1347 & _GEN_1283 & stq_15_bits_data_valid;
  wire        _GEN_55024 = _GEN_1444 & _GEN_1380 & _GEN_1348 & _GEN_1284 & stq_16_bits_data_valid;
  wire        _GEN_55025 = _GEN_1445 & _GEN_1381 & _GEN_1349 & _GEN_1285 & stq_17_bits_data_valid;
  wire        _GEN_55026 = _GEN_1446 & _GEN_1382 & _GEN_1350 & _GEN_1286 & stq_18_bits_data_valid;
  wire        _GEN_55027 = _GEN_1447 & _GEN_1383 & _GEN_1351 & _GEN_1287 & stq_19_bits_data_valid;
  wire        _GEN_55028 = _GEN_1448 & _GEN_1384 & _GEN_1352 & _GEN_1288 & stq_20_bits_data_valid;
  wire        _GEN_55029 = _GEN_1449 & _GEN_1385 & _GEN_1353 & _GEN_1289 & stq_21_bits_data_valid;
  wire        _GEN_55030 = _GEN_1450 & _GEN_1386 & _GEN_1354 & _GEN_1290 & stq_22_bits_data_valid;
  wire        _GEN_55031 = _GEN_1451 & _GEN_1387 & _GEN_1355 & _GEN_1291 & stq_23_bits_data_valid;
  wire        _GEN_55032 = _GEN_1452 & _GEN_1388 & _GEN_1356 & _GEN_1292 & stq_24_bits_data_valid;
  wire        _GEN_55033 = _GEN_1453 & _GEN_1389 & _GEN_1357 & _GEN_1293 & stq_25_bits_data_valid;
  wire        _GEN_55034 = _GEN_1454 & _GEN_1390 & _GEN_1358 & _GEN_1294 & stq_26_bits_data_valid;
  wire        _GEN_55035 = _GEN_1455 & _GEN_1391 & _GEN_1359 & _GEN_1295 & stq_27_bits_data_valid;
  wire        _GEN_55036 = _GEN_1456 & _GEN_1392 & _GEN_1360 & _GEN_1296 & stq_28_bits_data_valid;
  wire        _GEN_55037 = _GEN_1457 & _GEN_1393 & _GEN_1361 & _GEN_1297 & stq_29_bits_data_valid;
  wire        _GEN_55038 = _GEN_1458 & _GEN_1394 & _GEN_1362 & _GEN_1298 & stq_30_bits_data_valid;
  wire        _GEN_55039 = _GEN_1459 & _GEN_1395 & _GEN_1363 & _GEN_1299 & stq_31_bits_data_valid;
  wire        _GEN_55040 = _GEN_1428 & _GEN_1364 & _GEN_1332 & _GEN_1268 & stq_0_bits_committed;
  wire        _GEN_55041 = _GEN_1429 & _GEN_1365 & _GEN_1333 & _GEN_1269 & stq_1_bits_committed;
  wire        _GEN_55042 = _GEN_1430 & _GEN_1366 & _GEN_1334 & _GEN_1270 & stq_2_bits_committed;
  wire        _GEN_55043 = _GEN_1431 & _GEN_1367 & _GEN_1335 & _GEN_1271 & stq_3_bits_committed;
  wire        _GEN_55044 = _GEN_1432 & _GEN_1368 & _GEN_1336 & _GEN_1272 & stq_4_bits_committed;
  wire        _GEN_55045 = _GEN_1433 & _GEN_1369 & _GEN_1337 & _GEN_1273 & stq_5_bits_committed;
  wire        _GEN_55046 = _GEN_1434 & _GEN_1370 & _GEN_1338 & _GEN_1274 & stq_6_bits_committed;
  wire        _GEN_55047 = _GEN_1435 & _GEN_1371 & _GEN_1339 & _GEN_1275 & stq_7_bits_committed;
  wire        _GEN_55048 = _GEN_1436 & _GEN_1372 & _GEN_1340 & _GEN_1276 & stq_8_bits_committed;
  wire        _GEN_55049 = _GEN_1437 & _GEN_1373 & _GEN_1341 & _GEN_1277 & stq_9_bits_committed;
  wire        _GEN_55050 = _GEN_1438 & _GEN_1374 & _GEN_1342 & _GEN_1278 & stq_10_bits_committed;
  wire        _GEN_55051 = _GEN_1439 & _GEN_1375 & _GEN_1343 & _GEN_1279 & stq_11_bits_committed;
  wire        _GEN_55052 = _GEN_1440 & _GEN_1376 & _GEN_1344 & _GEN_1280 & stq_12_bits_committed;
  wire        _GEN_55053 = _GEN_1441 & _GEN_1377 & _GEN_1345 & _GEN_1281 & stq_13_bits_committed;
  wire        _GEN_55054 = _GEN_1442 & _GEN_1378 & _GEN_1346 & _GEN_1282 & stq_14_bits_committed;
  wire        _GEN_55055 = _GEN_1443 & _GEN_1379 & _GEN_1347 & _GEN_1283 & stq_15_bits_committed;
  wire        _GEN_55056 = _GEN_1444 & _GEN_1380 & _GEN_1348 & _GEN_1284 & stq_16_bits_committed;
  wire        _GEN_55057 = _GEN_1445 & _GEN_1381 & _GEN_1349 & _GEN_1285 & stq_17_bits_committed;
  wire        _GEN_55058 = _GEN_1446 & _GEN_1382 & _GEN_1350 & _GEN_1286 & stq_18_bits_committed;
  wire        _GEN_55059 = _GEN_1447 & _GEN_1383 & _GEN_1351 & _GEN_1287 & stq_19_bits_committed;
  wire        _GEN_55060 = _GEN_1448 & _GEN_1384 & _GEN_1352 & _GEN_1288 & stq_20_bits_committed;
  wire        _GEN_55061 = _GEN_1449 & _GEN_1385 & _GEN_1353 & _GEN_1289 & stq_21_bits_committed;
  wire        _GEN_55062 = _GEN_1450 & _GEN_1386 & _GEN_1354 & _GEN_1290 & stq_22_bits_committed;
  wire        _GEN_55063 = _GEN_1451 & _GEN_1387 & _GEN_1355 & _GEN_1291 & stq_23_bits_committed;
  wire        _GEN_55064 = _GEN_1452 & _GEN_1388 & _GEN_1356 & _GEN_1292 & stq_24_bits_committed;
  wire        _GEN_55065 = _GEN_1453 & _GEN_1389 & _GEN_1357 & _GEN_1293 & stq_25_bits_committed;
  wire        _GEN_55066 = _GEN_1454 & _GEN_1390 & _GEN_1358 & _GEN_1294 & stq_26_bits_committed;
  wire        _GEN_55067 = _GEN_1455 & _GEN_1391 & _GEN_1359 & _GEN_1295 & stq_27_bits_committed;
  wire        _GEN_55068 = _GEN_1456 & _GEN_1392 & _GEN_1360 & _GEN_1296 & stq_28_bits_committed;
  wire        _GEN_55069 = _GEN_1457 & _GEN_1393 & _GEN_1361 & _GEN_1297 & stq_29_bits_committed;
  wire        _GEN_55070 = _GEN_1458 & _GEN_1394 & _GEN_1362 & _GEN_1298 & stq_30_bits_committed;
  wire        _GEN_55071 = _GEN_1459 & _GEN_1395 & _GEN_1363 & _GEN_1299 & stq_31_bits_committed;
  wire        _GEN_1460 = ldq_incoming_idx_1 == 5'h1;
  wire        _GEN_1461 = ldq_incoming_idx_1 == 5'h2;
  wire        _GEN_1462 = ldq_incoming_idx_1 == 5'h3;
  wire        _GEN_1463 = ldq_incoming_idx_1 == 5'h4;
  wire        _GEN_1464 = ldq_incoming_idx_1 == 5'h5;
  wire        _GEN_1465 = ldq_incoming_idx_1 == 5'h6;
  wire        _GEN_1466 = ldq_incoming_idx_1 == 5'h7;
  wire        _GEN_1467 = ldq_incoming_idx_1 == 5'h8;
  wire        _GEN_1468 = ldq_incoming_idx_1 == 5'h9;
  wire        _GEN_1469 = ldq_incoming_idx_1 == 5'hA;
  wire        _GEN_1470 = ldq_incoming_idx_1 == 5'hB;
  wire        _GEN_1471 = ldq_incoming_idx_1 == 5'hC;
  wire        _GEN_1472 = ldq_incoming_idx_1 == 5'hD;
  wire        _GEN_1473 = ldq_incoming_idx_1 == 5'hE;
  wire        _GEN_1474 = ldq_incoming_idx_1 == 5'hF;
  wire        _GEN_1475 = ldq_incoming_idx_1 == 5'h10;
  wire        _GEN_1476 = ldq_incoming_idx_1 == 5'h11;
  wire        _GEN_1477 = ldq_incoming_idx_1 == 5'h12;
  wire        _GEN_1478 = ldq_incoming_idx_1 == 5'h13;
  wire        _GEN_1479 = ldq_incoming_idx_1 == 5'h14;
  wire        _GEN_1480 = ldq_incoming_idx_1 == 5'h15;
  wire        _GEN_1481 = ldq_incoming_idx_1 == 5'h16;
  wire        _GEN_1482 = ldq_incoming_idx_1 == 5'h17;
  wire        _GEN_1483 = ldq_incoming_idx_1 == 5'h18;
  wire        _GEN_1484 = ldq_incoming_idx_1 == 5'h19;
  wire        _GEN_1485 = ldq_incoming_idx_1 == 5'h1A;
  wire        _GEN_1486 = ldq_incoming_idx_1 == 5'h1B;
  wire        _GEN_1487 = ldq_incoming_idx_1 == 5'h1C;
  wire        _GEN_1488 = ldq_incoming_idx_1 == 5'h1D;
  wire        _GEN_1489 = ldq_incoming_idx_1 == 5'h1E;
  wire        _GEN_1490 = ldq_wakeup_idx == 5'h1;
  wire        _GEN_1491 = ldq_wakeup_idx == 5'h2;
  wire        _GEN_1492 = ldq_wakeup_idx == 5'h3;
  wire        _GEN_1493 = ldq_wakeup_idx == 5'h4;
  wire        _GEN_1494 = ldq_wakeup_idx == 5'h5;
  wire        _GEN_1495 = ldq_wakeup_idx == 5'h6;
  wire        _GEN_1496 = ldq_wakeup_idx == 5'h7;
  wire        _GEN_1497 = ldq_wakeup_idx == 5'h8;
  wire        _GEN_1498 = ldq_wakeup_idx == 5'h9;
  wire        _GEN_1499 = ldq_wakeup_idx == 5'hA;
  wire        _GEN_1500 = ldq_wakeup_idx == 5'hB;
  wire        _GEN_1501 = ldq_wakeup_idx == 5'hC;
  wire        _GEN_1502 = ldq_wakeup_idx == 5'hD;
  wire        _GEN_1503 = ldq_wakeup_idx == 5'hE;
  wire        _GEN_1504 = ldq_wakeup_idx == 5'hF;
  wire        _GEN_1505 = ldq_wakeup_idx == 5'h10;
  wire        _GEN_1506 = ldq_wakeup_idx == 5'h11;
  wire        _GEN_1507 = ldq_wakeup_idx == 5'h12;
  wire        _GEN_1508 = ldq_wakeup_idx == 5'h13;
  wire        _GEN_1509 = ldq_wakeup_idx == 5'h14;
  wire        _GEN_1510 = ldq_wakeup_idx == 5'h15;
  wire        _GEN_1511 = ldq_wakeup_idx == 5'h16;
  wire        _GEN_1512 = ldq_wakeup_idx == 5'h17;
  wire        _GEN_1513 = ldq_wakeup_idx == 5'h18;
  wire        _GEN_1514 = ldq_wakeup_idx == 5'h19;
  wire        _GEN_1515 = ldq_wakeup_idx == 5'h1A;
  wire        _GEN_1516 = ldq_wakeup_idx == 5'h1B;
  wire        _GEN_1517 = ldq_wakeup_idx == 5'h1C;
  wire        _GEN_1518 = ldq_wakeup_idx == 5'h1D;
  wire        _GEN_1519 = ldq_wakeup_idx == 5'h1E;
  wire        _GEN_1520 = ldq_retry_idx == 5'h1;
  wire        _GEN_1521 = ldq_retry_idx == 5'h2;
  wire        _GEN_1522 = ldq_retry_idx == 5'h3;
  wire        _GEN_1523 = ldq_retry_idx == 5'h4;
  wire        _GEN_1524 = ldq_retry_idx == 5'h5;
  wire        _GEN_1525 = ldq_retry_idx == 5'h6;
  wire        _GEN_1526 = ldq_retry_idx == 5'h7;
  wire        _GEN_1527 = ldq_retry_idx == 5'h8;
  wire        _GEN_1528 = ldq_retry_idx == 5'h9;
  wire        _GEN_1529 = ldq_retry_idx == 5'hA;
  wire        _GEN_1530 = ldq_retry_idx == 5'hB;
  wire        _GEN_1531 = ldq_retry_idx == 5'hC;
  wire        _GEN_1532 = ldq_retry_idx == 5'hD;
  wire        _GEN_1533 = ldq_retry_idx == 5'hE;
  wire        _GEN_1534 = ldq_retry_idx == 5'hF;
  wire        _GEN_1535 = ldq_retry_idx == 5'h10;
  wire        _GEN_1536 = ldq_retry_idx == 5'h11;
  wire        _GEN_1537 = ldq_retry_idx == 5'h12;
  wire        _GEN_1538 = ldq_retry_idx == 5'h13;
  wire        _GEN_1539 = ldq_retry_idx == 5'h14;
  wire        _GEN_1540 = ldq_retry_idx == 5'h15;
  wire        _GEN_1541 = ldq_retry_idx == 5'h16;
  wire        _GEN_1542 = ldq_retry_idx == 5'h17;
  wire        _GEN_1543 = ldq_retry_idx == 5'h18;
  wire        _GEN_1544 = ldq_retry_idx == 5'h19;
  wire        _GEN_1545 = ldq_retry_idx == 5'h1A;
  wire        _GEN_1546 = ldq_retry_idx == 5'h1B;
  wire        _GEN_1547 = ldq_retry_idx == 5'h1C;
  wire        _GEN_1548 = ldq_retry_idx == 5'h1D;
  wire        _GEN_1549 = ldq_retry_idx == 5'h1E;
  wire        _GEN_68500 = can_fire_load_incoming_0 & ~(|ldq_incoming_idx_0);
  wire        _GEN_1550 = ldq_wakeup_idx == 5'h0;
  wire        _GEN_68532 = _GEN_1550 | _GEN_68500;
  wire        _GEN_1551 = ldq_incoming_idx_1 == 5'h0;
  wire        _GEN_68564 = _GEN_1551 | _GEN_68500;
  wire        _GEN_1552 = ldq_retry_idx == 5'h0;
  wire        _GEN_68628 = will_fire_load_retry_1 & _GEN_1552 | _GEN_68500;
  wire        ldq_retry_idx_block = (will_fire_load_wakeup_1 ? _GEN_68532 : can_fire_load_incoming_1 ? _GEN_68564 : _GEN_68628) | p1_block_load_mask_0;
  wire        _ldq_retry_idx_T_2 = ldq_0_bits_addr_valid & ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;
  wire        _GEN_68501 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1;
  wire        _GEN_68533 = _GEN_1490 | _GEN_68501;
  wire        _GEN_68565 = _GEN_1460 | _GEN_68501;
  wire        _GEN_68629 = will_fire_load_retry_1 & _GEN_1520 | _GEN_68501;
  wire        ldq_retry_idx_block_1 = (will_fire_load_wakeup_1 ? _GEN_68533 : can_fire_load_incoming_1 ? _GEN_68565 : _GEN_68629) | p1_block_load_mask_1;
  wire        _ldq_retry_idx_T_5 = ldq_1_bits_addr_valid & ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;
  wire        _GEN_68502 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h2;
  wire        _GEN_68534 = _GEN_1491 | _GEN_68502;
  wire        _GEN_68566 = _GEN_1461 | _GEN_68502;
  wire        _GEN_68630 = will_fire_load_retry_1 & _GEN_1521 | _GEN_68502;
  wire        ldq_retry_idx_block_2 = (will_fire_load_wakeup_1 ? _GEN_68534 : can_fire_load_incoming_1 ? _GEN_68566 : _GEN_68630) | p1_block_load_mask_2;
  wire        _ldq_retry_idx_T_8 = ldq_2_bits_addr_valid & ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;
  wire        _GEN_68503 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h3;
  wire        _GEN_68535 = _GEN_1492 | _GEN_68503;
  wire        _GEN_68567 = _GEN_1462 | _GEN_68503;
  wire        _GEN_68631 = will_fire_load_retry_1 & _GEN_1522 | _GEN_68503;
  wire        ldq_retry_idx_block_3 = (will_fire_load_wakeup_1 ? _GEN_68535 : can_fire_load_incoming_1 ? _GEN_68567 : _GEN_68631) | p1_block_load_mask_3;
  wire        _ldq_retry_idx_T_11 = ldq_3_bits_addr_valid & ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;
  wire        _GEN_68504 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h4;
  wire        _GEN_68536 = _GEN_1493 | _GEN_68504;
  wire        _GEN_68568 = _GEN_1463 | _GEN_68504;
  wire        _GEN_68632 = will_fire_load_retry_1 & _GEN_1523 | _GEN_68504;
  wire        ldq_retry_idx_block_4 = (will_fire_load_wakeup_1 ? _GEN_68536 : can_fire_load_incoming_1 ? _GEN_68568 : _GEN_68632) | p1_block_load_mask_4;
  wire        _ldq_retry_idx_T_14 = ldq_4_bits_addr_valid & ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;
  wire        _GEN_68505 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h5;
  wire        _GEN_68537 = _GEN_1494 | _GEN_68505;
  wire        _GEN_68569 = _GEN_1464 | _GEN_68505;
  wire        _GEN_68633 = will_fire_load_retry_1 & _GEN_1524 | _GEN_68505;
  wire        ldq_retry_idx_block_5 = (will_fire_load_wakeup_1 ? _GEN_68537 : can_fire_load_incoming_1 ? _GEN_68569 : _GEN_68633) | p1_block_load_mask_5;
  wire        _ldq_retry_idx_T_17 = ldq_5_bits_addr_valid & ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;
  wire        _GEN_68506 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h6;
  wire        _GEN_68538 = _GEN_1495 | _GEN_68506;
  wire        _GEN_68570 = _GEN_1465 | _GEN_68506;
  wire        _GEN_68634 = will_fire_load_retry_1 & _GEN_1525 | _GEN_68506;
  wire        ldq_retry_idx_block_6 = (will_fire_load_wakeup_1 ? _GEN_68538 : can_fire_load_incoming_1 ? _GEN_68570 : _GEN_68634) | p1_block_load_mask_6;
  wire        _ldq_retry_idx_T_20 = ldq_6_bits_addr_valid & ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;
  wire        _GEN_68507 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h7;
  wire        _GEN_68539 = _GEN_1496 | _GEN_68507;
  wire        _GEN_68571 = _GEN_1466 | _GEN_68507;
  wire        _GEN_68635 = will_fire_load_retry_1 & _GEN_1526 | _GEN_68507;
  wire        ldq_retry_idx_block_7 = (will_fire_load_wakeup_1 ? _GEN_68539 : can_fire_load_incoming_1 ? _GEN_68571 : _GEN_68635) | p1_block_load_mask_7;
  wire        _ldq_retry_idx_T_23 = ldq_7_bits_addr_valid & ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;
  wire        _GEN_68508 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h8;
  wire        _GEN_68540 = _GEN_1497 | _GEN_68508;
  wire        _GEN_68572 = _GEN_1467 | _GEN_68508;
  wire        _GEN_68636 = will_fire_load_retry_1 & _GEN_1527 | _GEN_68508;
  wire        ldq_retry_idx_block_8 = (will_fire_load_wakeup_1 ? _GEN_68540 : can_fire_load_incoming_1 ? _GEN_68572 : _GEN_68636) | p1_block_load_mask_8;
  wire        _ldq_retry_idx_T_26 = ldq_8_bits_addr_valid & ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;
  wire        _GEN_68509 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h9;
  wire        _GEN_68541 = _GEN_1498 | _GEN_68509;
  wire        _GEN_68573 = _GEN_1468 | _GEN_68509;
  wire        _GEN_68637 = will_fire_load_retry_1 & _GEN_1528 | _GEN_68509;
  wire        ldq_retry_idx_block_9 = (will_fire_load_wakeup_1 ? _GEN_68541 : can_fire_load_incoming_1 ? _GEN_68573 : _GEN_68637) | p1_block_load_mask_9;
  wire        _ldq_retry_idx_T_29 = ldq_9_bits_addr_valid & ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;
  wire        _GEN_68510 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hA;
  wire        _GEN_68542 = _GEN_1499 | _GEN_68510;
  wire        _GEN_68574 = _GEN_1469 | _GEN_68510;
  wire        _GEN_68638 = will_fire_load_retry_1 & _GEN_1529 | _GEN_68510;
  wire        ldq_retry_idx_block_10 = (will_fire_load_wakeup_1 ? _GEN_68542 : can_fire_load_incoming_1 ? _GEN_68574 : _GEN_68638) | p1_block_load_mask_10;
  wire        _ldq_retry_idx_T_32 = ldq_10_bits_addr_valid & ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;
  wire        _GEN_68511 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hB;
  wire        _GEN_68543 = _GEN_1500 | _GEN_68511;
  wire        _GEN_68575 = _GEN_1470 | _GEN_68511;
  wire        _GEN_68639 = will_fire_load_retry_1 & _GEN_1530 | _GEN_68511;
  wire        ldq_retry_idx_block_11 = (will_fire_load_wakeup_1 ? _GEN_68543 : can_fire_load_incoming_1 ? _GEN_68575 : _GEN_68639) | p1_block_load_mask_11;
  wire        _ldq_retry_idx_T_35 = ldq_11_bits_addr_valid & ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;
  wire        _GEN_68512 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hC;
  wire        _GEN_68544 = _GEN_1501 | _GEN_68512;
  wire        _GEN_68576 = _GEN_1471 | _GEN_68512;
  wire        _GEN_68640 = will_fire_load_retry_1 & _GEN_1531 | _GEN_68512;
  wire        ldq_retry_idx_block_12 = (will_fire_load_wakeup_1 ? _GEN_68544 : can_fire_load_incoming_1 ? _GEN_68576 : _GEN_68640) | p1_block_load_mask_12;
  wire        _ldq_retry_idx_T_38 = ldq_12_bits_addr_valid & ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;
  wire        _GEN_68513 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hD;
  wire        _GEN_68545 = _GEN_1502 | _GEN_68513;
  wire        _GEN_68577 = _GEN_1472 | _GEN_68513;
  wire        _GEN_68641 = will_fire_load_retry_1 & _GEN_1532 | _GEN_68513;
  wire        ldq_retry_idx_block_13 = (will_fire_load_wakeup_1 ? _GEN_68545 : can_fire_load_incoming_1 ? _GEN_68577 : _GEN_68641) | p1_block_load_mask_13;
  wire        _ldq_retry_idx_T_41 = ldq_13_bits_addr_valid & ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;
  wire        _GEN_68514 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hE;
  wire        _GEN_68546 = _GEN_1503 | _GEN_68514;
  wire        _GEN_68578 = _GEN_1473 | _GEN_68514;
  wire        _GEN_68642 = will_fire_load_retry_1 & _GEN_1533 | _GEN_68514;
  wire        ldq_retry_idx_block_14 = (will_fire_load_wakeup_1 ? _GEN_68546 : can_fire_load_incoming_1 ? _GEN_68578 : _GEN_68642) | p1_block_load_mask_14;
  wire        _ldq_retry_idx_T_44 = ldq_14_bits_addr_valid & ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;
  wire        _GEN_68515 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hF;
  wire        _GEN_68547 = _GEN_1504 | _GEN_68515;
  wire        _GEN_68579 = _GEN_1474 | _GEN_68515;
  wire        _GEN_68643 = will_fire_load_retry_1 & _GEN_1534 | _GEN_68515;
  wire        ldq_retry_idx_block_15 = (will_fire_load_wakeup_1 ? _GEN_68547 : can_fire_load_incoming_1 ? _GEN_68579 : _GEN_68643) | p1_block_load_mask_15;
  wire        _ldq_retry_idx_T_47 = ldq_15_bits_addr_valid & ldq_15_bits_addr_is_virtual & ~ldq_retry_idx_block_15;
  wire        _GEN_68516 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h10;
  wire        _GEN_68548 = _GEN_1505 | _GEN_68516;
  wire        _GEN_68580 = _GEN_1475 | _GEN_68516;
  wire        _GEN_68644 = will_fire_load_retry_1 & _GEN_1535 | _GEN_68516;
  wire        ldq_retry_idx_block_16 = (will_fire_load_wakeup_1 ? _GEN_68548 : can_fire_load_incoming_1 ? _GEN_68580 : _GEN_68644) | p1_block_load_mask_16;
  wire        _ldq_retry_idx_T_50 = ldq_16_bits_addr_valid & ldq_16_bits_addr_is_virtual & ~ldq_retry_idx_block_16;
  wire        _GEN_68517 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h11;
  wire        _GEN_68549 = _GEN_1506 | _GEN_68517;
  wire        _GEN_68581 = _GEN_1476 | _GEN_68517;
  wire        _GEN_68645 = will_fire_load_retry_1 & _GEN_1536 | _GEN_68517;
  wire        ldq_retry_idx_block_17 = (will_fire_load_wakeup_1 ? _GEN_68549 : can_fire_load_incoming_1 ? _GEN_68581 : _GEN_68645) | p1_block_load_mask_17;
  wire        _ldq_retry_idx_T_53 = ldq_17_bits_addr_valid & ldq_17_bits_addr_is_virtual & ~ldq_retry_idx_block_17;
  wire        _GEN_68518 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h12;
  wire        _GEN_68550 = _GEN_1507 | _GEN_68518;
  wire        _GEN_68582 = _GEN_1477 | _GEN_68518;
  wire        _GEN_68646 = will_fire_load_retry_1 & _GEN_1537 | _GEN_68518;
  wire        ldq_retry_idx_block_18 = (will_fire_load_wakeup_1 ? _GEN_68550 : can_fire_load_incoming_1 ? _GEN_68582 : _GEN_68646) | p1_block_load_mask_18;
  wire        _ldq_retry_idx_T_56 = ldq_18_bits_addr_valid & ldq_18_bits_addr_is_virtual & ~ldq_retry_idx_block_18;
  wire        _GEN_68519 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h13;
  wire        _GEN_68551 = _GEN_1508 | _GEN_68519;
  wire        _GEN_68583 = _GEN_1478 | _GEN_68519;
  wire        _GEN_68647 = will_fire_load_retry_1 & _GEN_1538 | _GEN_68519;
  wire        ldq_retry_idx_block_19 = (will_fire_load_wakeup_1 ? _GEN_68551 : can_fire_load_incoming_1 ? _GEN_68583 : _GEN_68647) | p1_block_load_mask_19;
  wire        _ldq_retry_idx_T_59 = ldq_19_bits_addr_valid & ldq_19_bits_addr_is_virtual & ~ldq_retry_idx_block_19;
  wire        _GEN_68520 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h14;
  wire        _GEN_68552 = _GEN_1509 | _GEN_68520;
  wire        _GEN_68584 = _GEN_1479 | _GEN_68520;
  wire        _GEN_68648 = will_fire_load_retry_1 & _GEN_1539 | _GEN_68520;
  wire        ldq_retry_idx_block_20 = (will_fire_load_wakeup_1 ? _GEN_68552 : can_fire_load_incoming_1 ? _GEN_68584 : _GEN_68648) | p1_block_load_mask_20;
  wire        _ldq_retry_idx_T_62 = ldq_20_bits_addr_valid & ldq_20_bits_addr_is_virtual & ~ldq_retry_idx_block_20;
  wire        _GEN_68521 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h15;
  wire        _GEN_68553 = _GEN_1510 | _GEN_68521;
  wire        _GEN_68585 = _GEN_1480 | _GEN_68521;
  wire        _GEN_68649 = will_fire_load_retry_1 & _GEN_1540 | _GEN_68521;
  wire        ldq_retry_idx_block_21 = (will_fire_load_wakeup_1 ? _GEN_68553 : can_fire_load_incoming_1 ? _GEN_68585 : _GEN_68649) | p1_block_load_mask_21;
  wire        _ldq_retry_idx_T_65 = ldq_21_bits_addr_valid & ldq_21_bits_addr_is_virtual & ~ldq_retry_idx_block_21;
  wire        _GEN_68522 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h16;
  wire        _GEN_68554 = _GEN_1511 | _GEN_68522;
  wire        _GEN_68586 = _GEN_1481 | _GEN_68522;
  wire        _GEN_68650 = will_fire_load_retry_1 & _GEN_1541 | _GEN_68522;
  wire        ldq_retry_idx_block_22 = (will_fire_load_wakeup_1 ? _GEN_68554 : can_fire_load_incoming_1 ? _GEN_68586 : _GEN_68650) | p1_block_load_mask_22;
  wire        _ldq_retry_idx_T_68 = ldq_22_bits_addr_valid & ldq_22_bits_addr_is_virtual & ~ldq_retry_idx_block_22;
  wire        _GEN_68523 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h17;
  wire        _GEN_68555 = _GEN_1512 | _GEN_68523;
  wire        _GEN_68587 = _GEN_1482 | _GEN_68523;
  wire        _GEN_68651 = will_fire_load_retry_1 & _GEN_1542 | _GEN_68523;
  wire        ldq_retry_idx_block_23 = (will_fire_load_wakeup_1 ? _GEN_68555 : can_fire_load_incoming_1 ? _GEN_68587 : _GEN_68651) | p1_block_load_mask_23;
  wire        _ldq_retry_idx_T_71 = ldq_23_bits_addr_valid & ldq_23_bits_addr_is_virtual & ~ldq_retry_idx_block_23;
  wire        _GEN_68524 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h18;
  wire        _GEN_68556 = _GEN_1513 | _GEN_68524;
  wire        _GEN_68588 = _GEN_1483 | _GEN_68524;
  wire        _GEN_68652 = will_fire_load_retry_1 & _GEN_1543 | _GEN_68524;
  wire        ldq_retry_idx_block_24 = (will_fire_load_wakeup_1 ? _GEN_68556 : can_fire_load_incoming_1 ? _GEN_68588 : _GEN_68652) | p1_block_load_mask_24;
  wire        _ldq_retry_idx_T_74 = ldq_24_bits_addr_valid & ldq_24_bits_addr_is_virtual & ~ldq_retry_idx_block_24;
  wire        _GEN_68525 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h19;
  wire        _GEN_68557 = _GEN_1514 | _GEN_68525;
  wire        _GEN_68589 = _GEN_1484 | _GEN_68525;
  wire        _GEN_68653 = will_fire_load_retry_1 & _GEN_1544 | _GEN_68525;
  wire        ldq_retry_idx_block_25 = (will_fire_load_wakeup_1 ? _GEN_68557 : can_fire_load_incoming_1 ? _GEN_68589 : _GEN_68653) | p1_block_load_mask_25;
  wire        _ldq_retry_idx_T_77 = ldq_25_bits_addr_valid & ldq_25_bits_addr_is_virtual & ~ldq_retry_idx_block_25;
  wire        _GEN_68526 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1A;
  wire        _GEN_68558 = _GEN_1515 | _GEN_68526;
  wire        _GEN_68590 = _GEN_1485 | _GEN_68526;
  wire        _GEN_68654 = will_fire_load_retry_1 & _GEN_1545 | _GEN_68526;
  wire        ldq_retry_idx_block_26 = (will_fire_load_wakeup_1 ? _GEN_68558 : can_fire_load_incoming_1 ? _GEN_68590 : _GEN_68654) | p1_block_load_mask_26;
  wire        _ldq_retry_idx_T_80 = ldq_26_bits_addr_valid & ldq_26_bits_addr_is_virtual & ~ldq_retry_idx_block_26;
  wire        _GEN_68527 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1B;
  wire        _GEN_68559 = _GEN_1516 | _GEN_68527;
  wire        _GEN_68591 = _GEN_1486 | _GEN_68527;
  wire        _GEN_68655 = will_fire_load_retry_1 & _GEN_1546 | _GEN_68527;
  wire        ldq_retry_idx_block_27 = (will_fire_load_wakeup_1 ? _GEN_68559 : can_fire_load_incoming_1 ? _GEN_68591 : _GEN_68655) | p1_block_load_mask_27;
  wire        _ldq_retry_idx_T_83 = ldq_27_bits_addr_valid & ldq_27_bits_addr_is_virtual & ~ldq_retry_idx_block_27;
  wire        _GEN_68528 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1C;
  wire        _GEN_68560 = _GEN_1517 | _GEN_68528;
  wire        _GEN_68592 = _GEN_1487 | _GEN_68528;
  wire        _GEN_68656 = will_fire_load_retry_1 & _GEN_1547 | _GEN_68528;
  wire        ldq_retry_idx_block_28 = (will_fire_load_wakeup_1 ? _GEN_68560 : can_fire_load_incoming_1 ? _GEN_68592 : _GEN_68656) | p1_block_load_mask_28;
  wire        _ldq_retry_idx_T_86 = ldq_28_bits_addr_valid & ldq_28_bits_addr_is_virtual & ~ldq_retry_idx_block_28;
  wire        _GEN_68529 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1D;
  wire        _GEN_68561 = _GEN_1518 | _GEN_68529;
  wire        _GEN_68593 = _GEN_1488 | _GEN_68529;
  wire        _GEN_68657 = will_fire_load_retry_1 & _GEN_1548 | _GEN_68529;
  wire        ldq_retry_idx_block_29 = (will_fire_load_wakeup_1 ? _GEN_68561 : can_fire_load_incoming_1 ? _GEN_68593 : _GEN_68657) | p1_block_load_mask_29;
  wire        _ldq_retry_idx_T_89 = ldq_29_bits_addr_valid & ldq_29_bits_addr_is_virtual & ~ldq_retry_idx_block_29;
  wire        _GEN_68530 = can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1E;
  wire        _GEN_68562 = _GEN_1519 | _GEN_68530;
  wire        _GEN_68594 = _GEN_1489 | _GEN_68530;
  wire        _GEN_68658 = will_fire_load_retry_1 & _GEN_1549 | _GEN_68530;
  wire        ldq_retry_idx_block_30 = (will_fire_load_wakeup_1 ? _GEN_68562 : can_fire_load_incoming_1 ? _GEN_68594 : _GEN_68658) | p1_block_load_mask_30;
  wire        _ldq_retry_idx_T_92 = ldq_30_bits_addr_valid & ldq_30_bits_addr_is_virtual & ~ldq_retry_idx_block_30;
  wire        _GEN_68531 = can_fire_load_incoming_0 & (&ldq_incoming_idx_0);
  wire        _GEN_68563 = (&ldq_wakeup_idx) | _GEN_68531;
  wire        _GEN_68595 = (&ldq_incoming_idx_1) | _GEN_68531;
  wire        _GEN_68659 = will_fire_load_retry_1 & (&ldq_retry_idx) | _GEN_68531;
  wire        ldq_retry_idx_block_31 = (will_fire_load_wakeup_1 ? _GEN_68563 : can_fire_load_incoming_1 ? _GEN_68595 : _GEN_68659) | p1_block_load_mask_31;
  wire        _stq_retry_idx_T = stq_0_bits_addr_valid & stq_0_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_1 = stq_1_bits_addr_valid & stq_1_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_2 = stq_2_bits_addr_valid & stq_2_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_3 = stq_3_bits_addr_valid & stq_3_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_4 = stq_4_bits_addr_valid & stq_4_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_5 = stq_5_bits_addr_valid & stq_5_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_6 = stq_6_bits_addr_valid & stq_6_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_7 = stq_7_bits_addr_valid & stq_7_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_8 = stq_8_bits_addr_valid & stq_8_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_9 = stq_9_bits_addr_valid & stq_9_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_10 = stq_10_bits_addr_valid & stq_10_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_11 = stq_11_bits_addr_valid & stq_11_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_12 = stq_12_bits_addr_valid & stq_12_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_13 = stq_13_bits_addr_valid & stq_13_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_14 = stq_14_bits_addr_valid & stq_14_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_15 = stq_15_bits_addr_valid & stq_15_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_16 = stq_16_bits_addr_valid & stq_16_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_17 = stq_17_bits_addr_valid & stq_17_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_18 = stq_18_bits_addr_valid & stq_18_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_19 = stq_19_bits_addr_valid & stq_19_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_20 = stq_20_bits_addr_valid & stq_20_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_21 = stq_21_bits_addr_valid & stq_21_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_22 = stq_22_bits_addr_valid & stq_22_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_23 = stq_23_bits_addr_valid & stq_23_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_24 = stq_24_bits_addr_valid & stq_24_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_25 = stq_25_bits_addr_valid & stq_25_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_26 = stq_26_bits_addr_valid & stq_26_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_27 = stq_27_bits_addr_valid & stq_27_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_28 = stq_28_bits_addr_valid & stq_28_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_29 = stq_29_bits_addr_valid & stq_29_bits_addr_is_virtual;
  wire        _stq_retry_idx_T_30 = stq_30_bits_addr_valid & stq_30_bits_addr_is_virtual;
  wire        _ldq_wakeup_idx_T_7 = ldq_0_bits_addr_valid & ~ldq_0_bits_executed & ~ldq_0_bits_succeeded & ~ldq_0_bits_addr_is_virtual & ~ldq_retry_idx_block;
  wire        _ldq_wakeup_idx_T_15 = ldq_1_bits_addr_valid & ~ldq_1_bits_executed & ~ldq_1_bits_succeeded & ~ldq_1_bits_addr_is_virtual & ~ldq_retry_idx_block_1;
  wire        _ldq_wakeup_idx_T_23 = ldq_2_bits_addr_valid & ~ldq_2_bits_executed & ~ldq_2_bits_succeeded & ~ldq_2_bits_addr_is_virtual & ~ldq_retry_idx_block_2;
  wire        _ldq_wakeup_idx_T_31 = ldq_3_bits_addr_valid & ~ldq_3_bits_executed & ~ldq_3_bits_succeeded & ~ldq_3_bits_addr_is_virtual & ~ldq_retry_idx_block_3;
  wire        _ldq_wakeup_idx_T_39 = ldq_4_bits_addr_valid & ~ldq_4_bits_executed & ~ldq_4_bits_succeeded & ~ldq_4_bits_addr_is_virtual & ~ldq_retry_idx_block_4;
  wire        _ldq_wakeup_idx_T_47 = ldq_5_bits_addr_valid & ~ldq_5_bits_executed & ~ldq_5_bits_succeeded & ~ldq_5_bits_addr_is_virtual & ~ldq_retry_idx_block_5;
  wire        _ldq_wakeup_idx_T_55 = ldq_6_bits_addr_valid & ~ldq_6_bits_executed & ~ldq_6_bits_succeeded & ~ldq_6_bits_addr_is_virtual & ~ldq_retry_idx_block_6;
  wire        _ldq_wakeup_idx_T_63 = ldq_7_bits_addr_valid & ~ldq_7_bits_executed & ~ldq_7_bits_succeeded & ~ldq_7_bits_addr_is_virtual & ~ldq_retry_idx_block_7;
  wire        _ldq_wakeup_idx_T_71 = ldq_8_bits_addr_valid & ~ldq_8_bits_executed & ~ldq_8_bits_succeeded & ~ldq_8_bits_addr_is_virtual & ~ldq_retry_idx_block_8;
  wire        _ldq_wakeup_idx_T_79 = ldq_9_bits_addr_valid & ~ldq_9_bits_executed & ~ldq_9_bits_succeeded & ~ldq_9_bits_addr_is_virtual & ~ldq_retry_idx_block_9;
  wire        _ldq_wakeup_idx_T_87 = ldq_10_bits_addr_valid & ~ldq_10_bits_executed & ~ldq_10_bits_succeeded & ~ldq_10_bits_addr_is_virtual & ~ldq_retry_idx_block_10;
  wire        _ldq_wakeup_idx_T_95 = ldq_11_bits_addr_valid & ~ldq_11_bits_executed & ~ldq_11_bits_succeeded & ~ldq_11_bits_addr_is_virtual & ~ldq_retry_idx_block_11;
  wire        _ldq_wakeup_idx_T_103 = ldq_12_bits_addr_valid & ~ldq_12_bits_executed & ~ldq_12_bits_succeeded & ~ldq_12_bits_addr_is_virtual & ~ldq_retry_idx_block_12;
  wire        _ldq_wakeup_idx_T_111 = ldq_13_bits_addr_valid & ~ldq_13_bits_executed & ~ldq_13_bits_succeeded & ~ldq_13_bits_addr_is_virtual & ~ldq_retry_idx_block_13;
  wire        _ldq_wakeup_idx_T_119 = ldq_14_bits_addr_valid & ~ldq_14_bits_executed & ~ldq_14_bits_succeeded & ~ldq_14_bits_addr_is_virtual & ~ldq_retry_idx_block_14;
  wire        _ldq_wakeup_idx_T_127 = ldq_15_bits_addr_valid & ~ldq_15_bits_executed & ~ldq_15_bits_succeeded & ~ldq_15_bits_addr_is_virtual & ~ldq_retry_idx_block_15;
  wire        _ldq_wakeup_idx_T_135 = ldq_16_bits_addr_valid & ~ldq_16_bits_executed & ~ldq_16_bits_succeeded & ~ldq_16_bits_addr_is_virtual & ~ldq_retry_idx_block_16;
  wire        _ldq_wakeup_idx_T_143 = ldq_17_bits_addr_valid & ~ldq_17_bits_executed & ~ldq_17_bits_succeeded & ~ldq_17_bits_addr_is_virtual & ~ldq_retry_idx_block_17;
  wire        _ldq_wakeup_idx_T_151 = ldq_18_bits_addr_valid & ~ldq_18_bits_executed & ~ldq_18_bits_succeeded & ~ldq_18_bits_addr_is_virtual & ~ldq_retry_idx_block_18;
  wire        _ldq_wakeup_idx_T_159 = ldq_19_bits_addr_valid & ~ldq_19_bits_executed & ~ldq_19_bits_succeeded & ~ldq_19_bits_addr_is_virtual & ~ldq_retry_idx_block_19;
  wire        _ldq_wakeup_idx_T_167 = ldq_20_bits_addr_valid & ~ldq_20_bits_executed & ~ldq_20_bits_succeeded & ~ldq_20_bits_addr_is_virtual & ~ldq_retry_idx_block_20;
  wire        _ldq_wakeup_idx_T_175 = ldq_21_bits_addr_valid & ~ldq_21_bits_executed & ~ldq_21_bits_succeeded & ~ldq_21_bits_addr_is_virtual & ~ldq_retry_idx_block_21;
  wire        _ldq_wakeup_idx_T_183 = ldq_22_bits_addr_valid & ~ldq_22_bits_executed & ~ldq_22_bits_succeeded & ~ldq_22_bits_addr_is_virtual & ~ldq_retry_idx_block_22;
  wire        _ldq_wakeup_idx_T_191 = ldq_23_bits_addr_valid & ~ldq_23_bits_executed & ~ldq_23_bits_succeeded & ~ldq_23_bits_addr_is_virtual & ~ldq_retry_idx_block_23;
  wire        _ldq_wakeup_idx_T_199 = ldq_24_bits_addr_valid & ~ldq_24_bits_executed & ~ldq_24_bits_succeeded & ~ldq_24_bits_addr_is_virtual & ~ldq_retry_idx_block_24;
  wire        _ldq_wakeup_idx_T_207 = ldq_25_bits_addr_valid & ~ldq_25_bits_executed & ~ldq_25_bits_succeeded & ~ldq_25_bits_addr_is_virtual & ~ldq_retry_idx_block_25;
  wire        _ldq_wakeup_idx_T_215 = ldq_26_bits_addr_valid & ~ldq_26_bits_executed & ~ldq_26_bits_succeeded & ~ldq_26_bits_addr_is_virtual & ~ldq_retry_idx_block_26;
  wire        _ldq_wakeup_idx_T_223 = ldq_27_bits_addr_valid & ~ldq_27_bits_executed & ~ldq_27_bits_succeeded & ~ldq_27_bits_addr_is_virtual & ~ldq_retry_idx_block_27;
  wire        _ldq_wakeup_idx_T_231 = ldq_28_bits_addr_valid & ~ldq_28_bits_executed & ~ldq_28_bits_succeeded & ~ldq_28_bits_addr_is_virtual & ~ldq_retry_idx_block_28;
  wire        _ldq_wakeup_idx_T_239 = ldq_29_bits_addr_valid & ~ldq_29_bits_executed & ~ldq_29_bits_succeeded & ~ldq_29_bits_addr_is_virtual & ~ldq_retry_idx_block_29;
  wire        _ldq_wakeup_idx_T_247 = ldq_30_bits_addr_valid & ~ldq_30_bits_executed & ~ldq_30_bits_succeeded & ~ldq_30_bits_addr_is_virtual & ~ldq_retry_idx_block_30;
  wire        ma_ld_0 = can_fire_load_incoming_0 & exe_req_0_bits_mxcpt_valid;
  wire        ma_ld_1 = can_fire_load_incoming_1 & exe_req_1_bits_mxcpt_valid;
  wire        ma_st_0 = _stq_idx_T & exe_req_0_bits_mxcpt_valid;
  wire        ma_st_1 = _stq_idx_T_1 & exe_req_1_bits_mxcpt_valid;
  wire        pf_ld_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_ld & exe_tlb_uop_0_uses_ldq;
  wire        pf_ld_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_pf_ld & exe_tlb_uop_1_uses_ldq;
  wire        pf_st_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_pf_st & exe_tlb_uop_0_uses_stq;
  wire        pf_st_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_pf_st & exe_tlb_uop_1_uses_stq;
  wire        ae_ld_0 = ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_ae_ld & exe_tlb_uop_0_uses_ldq;
  wire        ae_ld_1 = ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_ae_ld & exe_tlb_uop_1_uses_ldq;
  wire        is_older = mem_xcpt_valids_1 & (mem_xcpt_uops_1_rob_idx < mem_xcpt_uops_0_rob_idx ^ mem_xcpt_uops_1_rob_idx < io_core_rob_head_idx ^ mem_xcpt_uops_0_rob_idx < io_core_rob_head_idx | ~mem_xcpt_valids_0);
  wire [6:0]  mem_xcpt_uop_rob_idx = is_older ? mem_xcpt_uops_1_rob_idx : mem_xcpt_uops_0_rob_idx;
  wire        dmem_req_fire_0 = dmem_req_0_valid & _dmem_req_fire_T_2;
  wire [4:0]  ldq_idx = can_fire_load_incoming_0 ? ldq_incoming_idx_0 : ldq_retry_idx;
  wire        _ldq_T_340_bits_addr_is_uncacheable = ~_dtlb_io_resp_0_cacheable & ~exe_tlb_miss_0;
  wire        _GEN_1553 = can_fire_load_incoming_0 & ldq_idx == 5'h0;
  wire        _GEN_1554 = can_fire_load_incoming_0 & ldq_idx == 5'h1;
  wire        _GEN_1555 = can_fire_load_incoming_0 & ldq_idx == 5'h2;
  wire        _GEN_1556 = can_fire_load_incoming_0 & ldq_idx == 5'h3;
  wire        _GEN_1557 = can_fire_load_incoming_0 & ldq_idx == 5'h4;
  wire        _GEN_1558 = can_fire_load_incoming_0 & ldq_idx == 5'h5;
  wire        _GEN_1559 = can_fire_load_incoming_0 & ldq_idx == 5'h6;
  wire        _GEN_1560 = can_fire_load_incoming_0 & ldq_idx == 5'h7;
  wire        _GEN_1561 = can_fire_load_incoming_0 & ldq_idx == 5'h8;
  wire        _GEN_1562 = can_fire_load_incoming_0 & ldq_idx == 5'h9;
  wire        _GEN_1563 = can_fire_load_incoming_0 & ldq_idx == 5'hA;
  wire        _GEN_1564 = can_fire_load_incoming_0 & ldq_idx == 5'hB;
  wire        _GEN_1565 = can_fire_load_incoming_0 & ldq_idx == 5'hC;
  wire        _GEN_1566 = can_fire_load_incoming_0 & ldq_idx == 5'hD;
  wire        _GEN_1567 = can_fire_load_incoming_0 & ldq_idx == 5'hE;
  wire        _GEN_1568 = can_fire_load_incoming_0 & ldq_idx == 5'hF;
  wire        _GEN_1569 = can_fire_load_incoming_0 & ldq_idx == 5'h10;
  wire        _GEN_1570 = can_fire_load_incoming_0 & ldq_idx == 5'h11;
  wire        _GEN_1571 = can_fire_load_incoming_0 & ldq_idx == 5'h12;
  wire        _GEN_1572 = can_fire_load_incoming_0 & ldq_idx == 5'h13;
  wire        _GEN_1573 = can_fire_load_incoming_0 & ldq_idx == 5'h14;
  wire        _GEN_1574 = can_fire_load_incoming_0 & ldq_idx == 5'h15;
  wire        _GEN_1575 = can_fire_load_incoming_0 & ldq_idx == 5'h16;
  wire        _GEN_1576 = can_fire_load_incoming_0 & ldq_idx == 5'h17;
  wire        _GEN_1577 = can_fire_load_incoming_0 & ldq_idx == 5'h18;
  wire        _GEN_1578 = can_fire_load_incoming_0 & ldq_idx == 5'h19;
  wire        _GEN_1579 = can_fire_load_incoming_0 & ldq_idx == 5'h1A;
  wire        _GEN_1580 = can_fire_load_incoming_0 & ldq_idx == 5'h1B;
  wire        _GEN_1581 = can_fire_load_incoming_0 & ldq_idx == 5'h1C;
  wire        _GEN_1582 = can_fire_load_incoming_0 & ldq_idx == 5'h1D;
  wire        _GEN_1583 = can_fire_load_incoming_0 & ldq_idx == 5'h1E;
  wire        _GEN_1584 = can_fire_load_incoming_0 & (&ldq_idx);
  wire [4:0]  stq_idx = _stq_idx_T ? stq_incoming_idx_0 : stq_retry_idx;
  wire        _GEN_1585 = _stq_idx_T & stq_idx == 5'h0;
  wire        _GEN_1586 = _stq_idx_T & stq_idx == 5'h1;
  wire        _GEN_1587 = _stq_idx_T & stq_idx == 5'h2;
  wire        _GEN_1588 = _stq_idx_T & stq_idx == 5'h3;
  wire        _GEN_1589 = _stq_idx_T & stq_idx == 5'h4;
  wire        _GEN_1590 = _stq_idx_T & stq_idx == 5'h5;
  wire        _GEN_1591 = _stq_idx_T & stq_idx == 5'h6;
  wire        _GEN_1592 = _stq_idx_T & stq_idx == 5'h7;
  wire        _GEN_1593 = _stq_idx_T & stq_idx == 5'h8;
  wire        _GEN_1594 = _stq_idx_T & stq_idx == 5'h9;
  wire        _GEN_1595 = _stq_idx_T & stq_idx == 5'hA;
  wire        _GEN_1596 = _stq_idx_T & stq_idx == 5'hB;
  wire        _GEN_1597 = _stq_idx_T & stq_idx == 5'hC;
  wire        _GEN_1598 = _stq_idx_T & stq_idx == 5'hD;
  wire        _GEN_1599 = _stq_idx_T & stq_idx == 5'hE;
  wire        _GEN_1600 = _stq_idx_T & stq_idx == 5'hF;
  wire        _GEN_1601 = _stq_idx_T & stq_idx == 5'h10;
  wire        _GEN_1602 = _stq_idx_T & stq_idx == 5'h11;
  wire        _GEN_1603 = _stq_idx_T & stq_idx == 5'h12;
  wire        _GEN_1604 = _stq_idx_T & stq_idx == 5'h13;
  wire        _GEN_1605 = _stq_idx_T & stq_idx == 5'h14;
  wire        _GEN_1606 = _stq_idx_T & stq_idx == 5'h15;
  wire        _GEN_1607 = _stq_idx_T & stq_idx == 5'h16;
  wire        _GEN_1608 = _stq_idx_T & stq_idx == 5'h17;
  wire        _GEN_1609 = _stq_idx_T & stq_idx == 5'h18;
  wire        _GEN_1610 = _stq_idx_T & stq_idx == 5'h19;
  wire        _GEN_1611 = _stq_idx_T & stq_idx == 5'h1A;
  wire        _GEN_1612 = _stq_idx_T & stq_idx == 5'h1B;
  wire        _GEN_1613 = _stq_idx_T & stq_idx == 5'h1C;
  wire        _GEN_1614 = _stq_idx_T & stq_idx == 5'h1D;
  wire        _GEN_1615 = _stq_idx_T & stq_idx == 5'h1E;
  wire        _GEN_1616 = _stq_idx_T & (&stq_idx);
  wire        _GEN_1617 = _GEN_335 & sidx == 5'h0;
  wire        _GEN_1618 = _GEN_335 & sidx == 5'h1;
  wire        _GEN_1619 = _GEN_335 & sidx == 5'h2;
  wire        _GEN_1620 = _GEN_335 & sidx == 5'h3;
  wire        _GEN_1621 = _GEN_335 & sidx == 5'h4;
  wire        _GEN_1622 = _GEN_335 & sidx == 5'h5;
  wire        _GEN_1623 = _GEN_335 & sidx == 5'h6;
  wire        _GEN_1624 = _GEN_335 & sidx == 5'h7;
  wire        _GEN_1625 = _GEN_335 & sidx == 5'h8;
  wire        _GEN_1626 = _GEN_335 & sidx == 5'h9;
  wire        _GEN_1627 = _GEN_335 & sidx == 5'hA;
  wire        _GEN_1628 = _GEN_335 & sidx == 5'hB;
  wire        _GEN_1629 = _GEN_335 & sidx == 5'hC;
  wire        _GEN_1630 = _GEN_335 & sidx == 5'hD;
  wire        _GEN_1631 = _GEN_335 & sidx == 5'hE;
  wire        _GEN_1632 = _GEN_335 & sidx == 5'hF;
  wire        _GEN_1633 = _GEN_335 & sidx == 5'h10;
  wire        _GEN_1634 = _GEN_335 & sidx == 5'h11;
  wire        _GEN_1635 = _GEN_335 & sidx == 5'h12;
  wire        _GEN_1636 = _GEN_335 & sidx == 5'h13;
  wire        _GEN_1637 = _GEN_335 & sidx == 5'h14;
  wire        _GEN_1638 = _GEN_335 & sidx == 5'h15;
  wire        _GEN_1639 = _GEN_335 & sidx == 5'h16;
  wire        _GEN_1640 = _GEN_335 & sidx == 5'h17;
  wire        _GEN_1641 = _GEN_335 & sidx == 5'h18;
  wire        _GEN_1642 = _GEN_335 & sidx == 5'h19;
  wire        _GEN_1643 = _GEN_335 & sidx == 5'h1A;
  wire        _GEN_1644 = _GEN_335 & sidx == 5'h1B;
  wire        _GEN_1645 = _GEN_335 & sidx == 5'h1C;
  wire        _GEN_1646 = _GEN_335 & sidx == 5'h1D;
  wire        _GEN_1647 = _GEN_335 & sidx == 5'h1E;
  wire        _GEN_1648 = _GEN_335 & (&sidx);
  wire [4:0]  ldq_idx_1 = can_fire_load_incoming_1 ? ldq_incoming_idx_1 : ldq_retry_idx;
  wire        _GEN_1649 = ldq_idx_1 == 5'h0;
  wire        _GEN_1650 = ldq_idx_1 == 5'h1;
  wire        _GEN_1651 = ldq_idx_1 == 5'h2;
  wire        _GEN_1652 = ldq_idx_1 == 5'h3;
  wire        _GEN_1653 = ldq_idx_1 == 5'h4;
  wire        _GEN_1654 = ldq_idx_1 == 5'h5;
  wire        _GEN_1655 = ldq_idx_1 == 5'h6;
  wire        _GEN_1656 = ldq_idx_1 == 5'h7;
  wire        _GEN_1657 = ldq_idx_1 == 5'h8;
  wire        _GEN_1658 = ldq_idx_1 == 5'h9;
  wire        _GEN_1659 = ldq_idx_1 == 5'hA;
  wire        _GEN_1660 = ldq_idx_1 == 5'hB;
  wire        _GEN_1661 = ldq_idx_1 == 5'hC;
  wire        _GEN_1662 = ldq_idx_1 == 5'hD;
  wire        _GEN_1663 = ldq_idx_1 == 5'hE;
  wire        _GEN_1664 = ldq_idx_1 == 5'hF;
  wire        _GEN_1665 = ldq_idx_1 == 5'h10;
  wire        _GEN_1666 = ldq_idx_1 == 5'h11;
  wire        _GEN_1667 = ldq_idx_1 == 5'h12;
  wire        _GEN_1668 = ldq_idx_1 == 5'h13;
  wire        _GEN_1669 = ldq_idx_1 == 5'h14;
  wire        _GEN_1670 = ldq_idx_1 == 5'h15;
  wire        _GEN_1671 = ldq_idx_1 == 5'h16;
  wire        _GEN_1672 = ldq_idx_1 == 5'h17;
  wire        _GEN_1673 = ldq_idx_1 == 5'h18;
  wire        _GEN_1674 = ldq_idx_1 == 5'h19;
  wire        _GEN_1675 = ldq_idx_1 == 5'h1A;
  wire        _GEN_1676 = ldq_idx_1 == 5'h1B;
  wire        _GEN_1677 = ldq_idx_1 == 5'h1C;
  wire        _GEN_1678 = ldq_idx_1 == 5'h1D;
  wire        _GEN_1679 = ldq_idx_1 == 5'h1E;
  wire        _ldq_T_403_bits_addr_is_uncacheable = ~_dtlb_io_resp_1_cacheable & ~exe_tlb_miss_1;
  wire        _GEN_81718 = _GEN_341 ? _GEN_1649 | _GEN_1553 | _GEN_52224 : _GEN_1553 | _GEN_52224;
  wire        _GEN_81719 = _GEN_341 ? _GEN_1650 | _GEN_1554 | _GEN_52225 : _GEN_1554 | _GEN_52225;
  wire        _GEN_81720 = _GEN_341 ? _GEN_1651 | _GEN_1555 | _GEN_52226 : _GEN_1555 | _GEN_52226;
  wire        _GEN_81721 = _GEN_341 ? _GEN_1652 | _GEN_1556 | _GEN_52227 : _GEN_1556 | _GEN_52227;
  wire        _GEN_81722 = _GEN_341 ? _GEN_1653 | _GEN_1557 | _GEN_52228 : _GEN_1557 | _GEN_52228;
  wire        _GEN_81723 = _GEN_341 ? _GEN_1654 | _GEN_1558 | _GEN_52229 : _GEN_1558 | _GEN_52229;
  wire        _GEN_81724 = _GEN_341 ? _GEN_1655 | _GEN_1559 | _GEN_52230 : _GEN_1559 | _GEN_52230;
  wire        _GEN_81725 = _GEN_341 ? _GEN_1656 | _GEN_1560 | _GEN_52231 : _GEN_1560 | _GEN_52231;
  wire        _GEN_81726 = _GEN_341 ? _GEN_1657 | _GEN_1561 | _GEN_52232 : _GEN_1561 | _GEN_52232;
  wire        _GEN_81727 = _GEN_341 ? _GEN_1658 | _GEN_1562 | _GEN_52233 : _GEN_1562 | _GEN_52233;
  wire        _GEN_81728 = _GEN_341 ? _GEN_1659 | _GEN_1563 | _GEN_52234 : _GEN_1563 | _GEN_52234;
  wire        _GEN_81729 = _GEN_341 ? _GEN_1660 | _GEN_1564 | _GEN_52235 : _GEN_1564 | _GEN_52235;
  wire        _GEN_81730 = _GEN_341 ? _GEN_1661 | _GEN_1565 | _GEN_52236 : _GEN_1565 | _GEN_52236;
  wire        _GEN_81731 = _GEN_341 ? _GEN_1662 | _GEN_1566 | _GEN_52237 : _GEN_1566 | _GEN_52237;
  wire        _GEN_81732 = _GEN_341 ? _GEN_1663 | _GEN_1567 | _GEN_52238 : _GEN_1567 | _GEN_52238;
  wire        _GEN_81733 = _GEN_341 ? _GEN_1664 | _GEN_1568 | _GEN_52239 : _GEN_1568 | _GEN_52239;
  wire        _GEN_81734 = _GEN_341 ? _GEN_1665 | _GEN_1569 | _GEN_52240 : _GEN_1569 | _GEN_52240;
  wire        _GEN_81735 = _GEN_341 ? _GEN_1666 | _GEN_1570 | _GEN_52241 : _GEN_1570 | _GEN_52241;
  wire        _GEN_81736 = _GEN_341 ? _GEN_1667 | _GEN_1571 | _GEN_52242 : _GEN_1571 | _GEN_52242;
  wire        _GEN_81737 = _GEN_341 ? _GEN_1668 | _GEN_1572 | _GEN_52243 : _GEN_1572 | _GEN_52243;
  wire        _GEN_81738 = _GEN_341 ? _GEN_1669 | _GEN_1573 | _GEN_52244 : _GEN_1573 | _GEN_52244;
  wire        _GEN_81739 = _GEN_341 ? _GEN_1670 | _GEN_1574 | _GEN_52245 : _GEN_1574 | _GEN_52245;
  wire        _GEN_81740 = _GEN_341 ? _GEN_1671 | _GEN_1575 | _GEN_52246 : _GEN_1575 | _GEN_52246;
  wire        _GEN_81741 = _GEN_341 ? _GEN_1672 | _GEN_1576 | _GEN_52247 : _GEN_1576 | _GEN_52247;
  wire        _GEN_81742 = _GEN_341 ? _GEN_1673 | _GEN_1577 | _GEN_52248 : _GEN_1577 | _GEN_52248;
  wire        _GEN_81743 = _GEN_341 ? _GEN_1674 | _GEN_1578 | _GEN_52249 : _GEN_1578 | _GEN_52249;
  wire        _GEN_81744 = _GEN_341 ? _GEN_1675 | _GEN_1579 | _GEN_52250 : _GEN_1579 | _GEN_52250;
  wire        _GEN_81745 = _GEN_341 ? _GEN_1676 | _GEN_1580 | _GEN_52251 : _GEN_1580 | _GEN_52251;
  wire        _GEN_81746 = _GEN_341 ? _GEN_1677 | _GEN_1581 | _GEN_52252 : _GEN_1581 | _GEN_52252;
  wire        _GEN_81747 = _GEN_341 ? _GEN_1678 | _GEN_1582 | _GEN_52253 : _GEN_1582 | _GEN_52253;
  wire        _GEN_81748 = _GEN_341 ? _GEN_1679 | _GEN_1583 | _GEN_52254 : _GEN_1583 | _GEN_52254;
  wire        _GEN_81749 = _GEN_341 ? (&ldq_idx_1) | _GEN_1584 | _GEN_52255 : _GEN_1584 | _GEN_52255;
  wire [4:0]  stq_idx_1 = _stq_idx_T_1 ? stq_incoming_idx_1 : stq_retry_idx;
  wire        _GEN_1680 = _GEN_342 & stq_idx_1 == 5'h0;
  wire        _GEN_82006 = _GEN_1680 ? ~pf_st_1 : _GEN_1585 ? ~pf_st_0 : _GEN_1428 & _GEN_1364 & _GEN_1332 & _GEN_1268 & stq_0_bits_addr_valid;
  wire        _GEN_1681 = _GEN_342 & stq_idx_1 == 5'h1;
  wire        _GEN_82007 = _GEN_1681 ? ~pf_st_1 : _GEN_1586 ? ~pf_st_0 : _GEN_1429 & _GEN_1365 & _GEN_1333 & _GEN_1269 & stq_1_bits_addr_valid;
  wire        _GEN_1682 = _GEN_342 & stq_idx_1 == 5'h2;
  wire        _GEN_82008 = _GEN_1682 ? ~pf_st_1 : _GEN_1587 ? ~pf_st_0 : _GEN_1430 & _GEN_1366 & _GEN_1334 & _GEN_1270 & stq_2_bits_addr_valid;
  wire        _GEN_1683 = _GEN_342 & stq_idx_1 == 5'h3;
  wire        _GEN_82009 = _GEN_1683 ? ~pf_st_1 : _GEN_1588 ? ~pf_st_0 : _GEN_1431 & _GEN_1367 & _GEN_1335 & _GEN_1271 & stq_3_bits_addr_valid;
  wire        _GEN_1684 = _GEN_342 & stq_idx_1 == 5'h4;
  wire        _GEN_82010 = _GEN_1684 ? ~pf_st_1 : _GEN_1589 ? ~pf_st_0 : _GEN_1432 & _GEN_1368 & _GEN_1336 & _GEN_1272 & stq_4_bits_addr_valid;
  wire        _GEN_1685 = _GEN_342 & stq_idx_1 == 5'h5;
  wire        _GEN_82011 = _GEN_1685 ? ~pf_st_1 : _GEN_1590 ? ~pf_st_0 : _GEN_1433 & _GEN_1369 & _GEN_1337 & _GEN_1273 & stq_5_bits_addr_valid;
  wire        _GEN_1686 = _GEN_342 & stq_idx_1 == 5'h6;
  wire        _GEN_82012 = _GEN_1686 ? ~pf_st_1 : _GEN_1591 ? ~pf_st_0 : _GEN_1434 & _GEN_1370 & _GEN_1338 & _GEN_1274 & stq_6_bits_addr_valid;
  wire        _GEN_1687 = _GEN_342 & stq_idx_1 == 5'h7;
  wire        _GEN_82013 = _GEN_1687 ? ~pf_st_1 : _GEN_1592 ? ~pf_st_0 : _GEN_1435 & _GEN_1371 & _GEN_1339 & _GEN_1275 & stq_7_bits_addr_valid;
  wire        _GEN_1688 = _GEN_342 & stq_idx_1 == 5'h8;
  wire        _GEN_82014 = _GEN_1688 ? ~pf_st_1 : _GEN_1593 ? ~pf_st_0 : _GEN_1436 & _GEN_1372 & _GEN_1340 & _GEN_1276 & stq_8_bits_addr_valid;
  wire        _GEN_1689 = _GEN_342 & stq_idx_1 == 5'h9;
  wire        _GEN_82015 = _GEN_1689 ? ~pf_st_1 : _GEN_1594 ? ~pf_st_0 : _GEN_1437 & _GEN_1373 & _GEN_1341 & _GEN_1277 & stq_9_bits_addr_valid;
  wire        _GEN_1690 = _GEN_342 & stq_idx_1 == 5'hA;
  wire        _GEN_82016 = _GEN_1690 ? ~pf_st_1 : _GEN_1595 ? ~pf_st_0 : _GEN_1438 & _GEN_1374 & _GEN_1342 & _GEN_1278 & stq_10_bits_addr_valid;
  wire        _GEN_1691 = _GEN_342 & stq_idx_1 == 5'hB;
  wire        _GEN_82017 = _GEN_1691 ? ~pf_st_1 : _GEN_1596 ? ~pf_st_0 : _GEN_1439 & _GEN_1375 & _GEN_1343 & _GEN_1279 & stq_11_bits_addr_valid;
  wire        _GEN_1692 = _GEN_342 & stq_idx_1 == 5'hC;
  wire        _GEN_82018 = _GEN_1692 ? ~pf_st_1 : _GEN_1597 ? ~pf_st_0 : _GEN_1440 & _GEN_1376 & _GEN_1344 & _GEN_1280 & stq_12_bits_addr_valid;
  wire        _GEN_1693 = _GEN_342 & stq_idx_1 == 5'hD;
  wire        _GEN_82019 = _GEN_1693 ? ~pf_st_1 : _GEN_1598 ? ~pf_st_0 : _GEN_1441 & _GEN_1377 & _GEN_1345 & _GEN_1281 & stq_13_bits_addr_valid;
  wire        _GEN_1694 = _GEN_342 & stq_idx_1 == 5'hE;
  wire        _GEN_82020 = _GEN_1694 ? ~pf_st_1 : _GEN_1599 ? ~pf_st_0 : _GEN_1442 & _GEN_1378 & _GEN_1346 & _GEN_1282 & stq_14_bits_addr_valid;
  wire        _GEN_1695 = _GEN_342 & stq_idx_1 == 5'hF;
  wire        _GEN_82021 = _GEN_1695 ? ~pf_st_1 : _GEN_1600 ? ~pf_st_0 : _GEN_1443 & _GEN_1379 & _GEN_1347 & _GEN_1283 & stq_15_bits_addr_valid;
  wire        _GEN_1696 = _GEN_342 & stq_idx_1 == 5'h10;
  wire        _GEN_82022 = _GEN_1696 ? ~pf_st_1 : _GEN_1601 ? ~pf_st_0 : _GEN_1444 & _GEN_1380 & _GEN_1348 & _GEN_1284 & stq_16_bits_addr_valid;
  wire        _GEN_1697 = _GEN_342 & stq_idx_1 == 5'h11;
  wire        _GEN_82023 = _GEN_1697 ? ~pf_st_1 : _GEN_1602 ? ~pf_st_0 : _GEN_1445 & _GEN_1381 & _GEN_1349 & _GEN_1285 & stq_17_bits_addr_valid;
  wire        _GEN_1698 = _GEN_342 & stq_idx_1 == 5'h12;
  wire        _GEN_82024 = _GEN_1698 ? ~pf_st_1 : _GEN_1603 ? ~pf_st_0 : _GEN_1446 & _GEN_1382 & _GEN_1350 & _GEN_1286 & stq_18_bits_addr_valid;
  wire        _GEN_1699 = _GEN_342 & stq_idx_1 == 5'h13;
  wire        _GEN_82025 = _GEN_1699 ? ~pf_st_1 : _GEN_1604 ? ~pf_st_0 : _GEN_1447 & _GEN_1383 & _GEN_1351 & _GEN_1287 & stq_19_bits_addr_valid;
  wire        _GEN_1700 = _GEN_342 & stq_idx_1 == 5'h14;
  wire        _GEN_82026 = _GEN_1700 ? ~pf_st_1 : _GEN_1605 ? ~pf_st_0 : _GEN_1448 & _GEN_1384 & _GEN_1352 & _GEN_1288 & stq_20_bits_addr_valid;
  wire        _GEN_1701 = _GEN_342 & stq_idx_1 == 5'h15;
  wire        _GEN_82027 = _GEN_1701 ? ~pf_st_1 : _GEN_1606 ? ~pf_st_0 : _GEN_1449 & _GEN_1385 & _GEN_1353 & _GEN_1289 & stq_21_bits_addr_valid;
  wire        _GEN_1702 = _GEN_342 & stq_idx_1 == 5'h16;
  wire        _GEN_82028 = _GEN_1702 ? ~pf_st_1 : _GEN_1607 ? ~pf_st_0 : _GEN_1450 & _GEN_1386 & _GEN_1354 & _GEN_1290 & stq_22_bits_addr_valid;
  wire        _GEN_1703 = _GEN_342 & stq_idx_1 == 5'h17;
  wire        _GEN_82029 = _GEN_1703 ? ~pf_st_1 : _GEN_1608 ? ~pf_st_0 : _GEN_1451 & _GEN_1387 & _GEN_1355 & _GEN_1291 & stq_23_bits_addr_valid;
  wire        _GEN_1704 = _GEN_342 & stq_idx_1 == 5'h18;
  wire        _GEN_82030 = _GEN_1704 ? ~pf_st_1 : _GEN_1609 ? ~pf_st_0 : _GEN_1452 & _GEN_1388 & _GEN_1356 & _GEN_1292 & stq_24_bits_addr_valid;
  wire        _GEN_1705 = _GEN_342 & stq_idx_1 == 5'h19;
  wire        _GEN_82031 = _GEN_1705 ? ~pf_st_1 : _GEN_1610 ? ~pf_st_0 : _GEN_1453 & _GEN_1389 & _GEN_1357 & _GEN_1293 & stq_25_bits_addr_valid;
  wire        _GEN_1706 = _GEN_342 & stq_idx_1 == 5'h1A;
  wire        _GEN_82032 = _GEN_1706 ? ~pf_st_1 : _GEN_1611 ? ~pf_st_0 : _GEN_1454 & _GEN_1390 & _GEN_1358 & _GEN_1294 & stq_26_bits_addr_valid;
  wire        _GEN_1707 = _GEN_342 & stq_idx_1 == 5'h1B;
  wire        _GEN_82033 = _GEN_1707 ? ~pf_st_1 : _GEN_1612 ? ~pf_st_0 : _GEN_1455 & _GEN_1391 & _GEN_1359 & _GEN_1295 & stq_27_bits_addr_valid;
  wire        _GEN_1708 = _GEN_342 & stq_idx_1 == 5'h1C;
  wire        _GEN_82034 = _GEN_1708 ? ~pf_st_1 : _GEN_1613 ? ~pf_st_0 : _GEN_1456 & _GEN_1392 & _GEN_1360 & _GEN_1296 & stq_28_bits_addr_valid;
  wire        _GEN_1709 = _GEN_342 & stq_idx_1 == 5'h1D;
  wire        _GEN_82035 = _GEN_1709 ? ~pf_st_1 : _GEN_1614 ? ~pf_st_0 : _GEN_1457 & _GEN_1393 & _GEN_1361 & _GEN_1297 & stq_29_bits_addr_valid;
  wire        _GEN_1710 = _GEN_342 & stq_idx_1 == 5'h1E;
  wire        _GEN_82036 = _GEN_1710 ? ~pf_st_1 : _GEN_1615 ? ~pf_st_0 : _GEN_1458 & _GEN_1394 & _GEN_1362 & _GEN_1298 & stq_30_bits_addr_valid;
  wire        _GEN_1711 = _GEN_342 & (&stq_idx_1);
  wire        _GEN_82037 = _GEN_1711 ? ~pf_st_1 : _GEN_1616 ? ~pf_st_0 : _GEN_1459 & _GEN_1395 & _GEN_1363 & _GEN_1299 & stq_31_bits_addr_valid;
  wire        _GEN_1712 = sidx_1 == 5'h0;
  wire        _GEN_1713 = sidx_1 == 5'h1;
  wire        _GEN_1714 = sidx_1 == 5'h2;
  wire        _GEN_1715 = sidx_1 == 5'h3;
  wire        _GEN_1716 = sidx_1 == 5'h4;
  wire        _GEN_1717 = sidx_1 == 5'h5;
  wire        _GEN_1718 = sidx_1 == 5'h6;
  wire        _GEN_1719 = sidx_1 == 5'h7;
  wire        _GEN_1720 = sidx_1 == 5'h8;
  wire        _GEN_1721 = sidx_1 == 5'h9;
  wire        _GEN_1722 = sidx_1 == 5'hA;
  wire        _GEN_1723 = sidx_1 == 5'hB;
  wire        _GEN_1724 = sidx_1 == 5'hC;
  wire        _GEN_1725 = sidx_1 == 5'hD;
  wire        _GEN_1726 = sidx_1 == 5'hE;
  wire        _GEN_1727 = sidx_1 == 5'hF;
  wire        _GEN_1728 = sidx_1 == 5'h10;
  wire        _GEN_1729 = sidx_1 == 5'h11;
  wire        _GEN_1730 = sidx_1 == 5'h12;
  wire        _GEN_1731 = sidx_1 == 5'h13;
  wire        _GEN_1732 = sidx_1 == 5'h14;
  wire        _GEN_1733 = sidx_1 == 5'h15;
  wire        _GEN_1734 = sidx_1 == 5'h16;
  wire        _GEN_1735 = sidx_1 == 5'h17;
  wire        _GEN_1736 = sidx_1 == 5'h18;
  wire        _GEN_1737 = sidx_1 == 5'h19;
  wire        _GEN_1738 = sidx_1 == 5'h1A;
  wire        _GEN_1739 = sidx_1 == 5'h1B;
  wire        _GEN_1740 = sidx_1 == 5'h1C;
  wire        _GEN_1741 = sidx_1 == 5'h1D;
  wire        _GEN_1742 = sidx_1 == 5'h1E;
  wire        _GEN_82230 = _stq_bits_data_bits_T_2 ? _GEN_1712 | _GEN_1617 | _GEN_55008 : _GEN_1617 | _GEN_55008;
  wire        _GEN_82231 = _stq_bits_data_bits_T_2 ? _GEN_1713 | _GEN_1618 | _GEN_55009 : _GEN_1618 | _GEN_55009;
  wire        _GEN_82232 = _stq_bits_data_bits_T_2 ? _GEN_1714 | _GEN_1619 | _GEN_55010 : _GEN_1619 | _GEN_55010;
  wire        _GEN_82233 = _stq_bits_data_bits_T_2 ? _GEN_1715 | _GEN_1620 | _GEN_55011 : _GEN_1620 | _GEN_55011;
  wire        _GEN_82234 = _stq_bits_data_bits_T_2 ? _GEN_1716 | _GEN_1621 | _GEN_55012 : _GEN_1621 | _GEN_55012;
  wire        _GEN_82235 = _stq_bits_data_bits_T_2 ? _GEN_1717 | _GEN_1622 | _GEN_55013 : _GEN_1622 | _GEN_55013;
  wire        _GEN_82236 = _stq_bits_data_bits_T_2 ? _GEN_1718 | _GEN_1623 | _GEN_55014 : _GEN_1623 | _GEN_55014;
  wire        _GEN_82237 = _stq_bits_data_bits_T_2 ? _GEN_1719 | _GEN_1624 | _GEN_55015 : _GEN_1624 | _GEN_55015;
  wire        _GEN_82238 = _stq_bits_data_bits_T_2 ? _GEN_1720 | _GEN_1625 | _GEN_55016 : _GEN_1625 | _GEN_55016;
  wire        _GEN_82239 = _stq_bits_data_bits_T_2 ? _GEN_1721 | _GEN_1626 | _GEN_55017 : _GEN_1626 | _GEN_55017;
  wire        _GEN_82240 = _stq_bits_data_bits_T_2 ? _GEN_1722 | _GEN_1627 | _GEN_55018 : _GEN_1627 | _GEN_55018;
  wire        _GEN_82241 = _stq_bits_data_bits_T_2 ? _GEN_1723 | _GEN_1628 | _GEN_55019 : _GEN_1628 | _GEN_55019;
  wire        _GEN_82242 = _stq_bits_data_bits_T_2 ? _GEN_1724 | _GEN_1629 | _GEN_55020 : _GEN_1629 | _GEN_55020;
  wire        _GEN_82243 = _stq_bits_data_bits_T_2 ? _GEN_1725 | _GEN_1630 | _GEN_55021 : _GEN_1630 | _GEN_55021;
  wire        _GEN_82244 = _stq_bits_data_bits_T_2 ? _GEN_1726 | _GEN_1631 | _GEN_55022 : _GEN_1631 | _GEN_55022;
  wire        _GEN_82245 = _stq_bits_data_bits_T_2 ? _GEN_1727 | _GEN_1632 | _GEN_55023 : _GEN_1632 | _GEN_55023;
  wire        _GEN_82246 = _stq_bits_data_bits_T_2 ? _GEN_1728 | _GEN_1633 | _GEN_55024 : _GEN_1633 | _GEN_55024;
  wire        _GEN_82247 = _stq_bits_data_bits_T_2 ? _GEN_1729 | _GEN_1634 | _GEN_55025 : _GEN_1634 | _GEN_55025;
  wire        _GEN_82248 = _stq_bits_data_bits_T_2 ? _GEN_1730 | _GEN_1635 | _GEN_55026 : _GEN_1635 | _GEN_55026;
  wire        _GEN_82249 = _stq_bits_data_bits_T_2 ? _GEN_1731 | _GEN_1636 | _GEN_55027 : _GEN_1636 | _GEN_55027;
  wire        _GEN_82250 = _stq_bits_data_bits_T_2 ? _GEN_1732 | _GEN_1637 | _GEN_55028 : _GEN_1637 | _GEN_55028;
  wire        _GEN_82251 = _stq_bits_data_bits_T_2 ? _GEN_1733 | _GEN_1638 | _GEN_55029 : _GEN_1638 | _GEN_55029;
  wire        _GEN_82252 = _stq_bits_data_bits_T_2 ? _GEN_1734 | _GEN_1639 | _GEN_55030 : _GEN_1639 | _GEN_55030;
  wire        _GEN_82253 = _stq_bits_data_bits_T_2 ? _GEN_1735 | _GEN_1640 | _GEN_55031 : _GEN_1640 | _GEN_55031;
  wire        _GEN_82254 = _stq_bits_data_bits_T_2 ? _GEN_1736 | _GEN_1641 | _GEN_55032 : _GEN_1641 | _GEN_55032;
  wire        _GEN_82255 = _stq_bits_data_bits_T_2 ? _GEN_1737 | _GEN_1642 | _GEN_55033 : _GEN_1642 | _GEN_55033;
  wire        _GEN_82256 = _stq_bits_data_bits_T_2 ? _GEN_1738 | _GEN_1643 | _GEN_55034 : _GEN_1643 | _GEN_55034;
  wire        _GEN_82257 = _stq_bits_data_bits_T_2 ? _GEN_1739 | _GEN_1644 | _GEN_55035 : _GEN_1644 | _GEN_55035;
  wire        _GEN_82258 = _stq_bits_data_bits_T_2 ? _GEN_1740 | _GEN_1645 | _GEN_55036 : _GEN_1645 | _GEN_55036;
  wire        _GEN_82259 = _stq_bits_data_bits_T_2 ? _GEN_1741 | _GEN_1646 | _GEN_55037 : _GEN_1646 | _GEN_55037;
  wire        _GEN_82260 = _stq_bits_data_bits_T_2 ? _GEN_1742 | _GEN_1647 | _GEN_55038 : _GEN_1647 | _GEN_55038;
  wire        _GEN_82261 = _stq_bits_data_bits_T_2 ? (&sidx_1) | _GEN_1648 | _GEN_55039 : _GEN_1648 | _GEN_55039;
  wire        _fired_std_incoming_T = (io_core_brupdate_b1_mispredict_mask & exe_req_0_bits_uop_br_mask) == 20'h0;
  wire        _fired_std_incoming_T_2 = (io_core_brupdate_b1_mispredict_mask & exe_req_1_bits_uop_br_mask) == 20'h0;
  wire        _GEN_1743 = lcam_ldq_idx_0 == 5'h1;
  wire        _GEN_1744 = lcam_ldq_idx_0 == 5'h2;
  wire        _GEN_1745 = lcam_ldq_idx_0 == 5'h3;
  wire        _GEN_1746 = lcam_ldq_idx_0 == 5'h4;
  wire        _GEN_1747 = lcam_ldq_idx_0 == 5'h5;
  wire        _GEN_1748 = lcam_ldq_idx_0 == 5'h6;
  wire        _GEN_1749 = lcam_ldq_idx_0 == 5'h7;
  wire        _GEN_1750 = lcam_ldq_idx_0 == 5'h8;
  wire        _GEN_1751 = lcam_ldq_idx_0 == 5'h9;
  wire        _GEN_1752 = lcam_ldq_idx_0 == 5'hA;
  wire        _GEN_1753 = lcam_ldq_idx_0 == 5'hB;
  wire        _GEN_1754 = lcam_ldq_idx_0 == 5'hC;
  wire        _GEN_1755 = lcam_ldq_idx_0 == 5'hD;
  wire        _GEN_1756 = lcam_ldq_idx_0 == 5'hE;
  wire        _GEN_1757 = lcam_ldq_idx_0 == 5'hF;
  wire        _GEN_1758 = lcam_ldq_idx_0 == 5'h10;
  wire        _GEN_1759 = lcam_ldq_idx_0 == 5'h11;
  wire        _GEN_1760 = lcam_ldq_idx_0 == 5'h12;
  wire        _GEN_1761 = lcam_ldq_idx_0 == 5'h13;
  wire        _GEN_1762 = lcam_ldq_idx_0 == 5'h14;
  wire        _GEN_1763 = lcam_ldq_idx_0 == 5'h15;
  wire        _GEN_1764 = lcam_ldq_idx_0 == 5'h16;
  wire        _GEN_1765 = lcam_ldq_idx_0 == 5'h17;
  wire        _GEN_1766 = lcam_ldq_idx_0 == 5'h18;
  wire        _GEN_1767 = lcam_ldq_idx_0 == 5'h19;
  wire        _GEN_1768 = lcam_ldq_idx_0 == 5'h1A;
  wire        _GEN_1769 = lcam_ldq_idx_0 == 5'h1B;
  wire        _GEN_1770 = lcam_ldq_idx_0 == 5'h1C;
  wire        _GEN_1771 = lcam_ldq_idx_0 == 5'h1D;
  wire        _GEN_1772 = lcam_ldq_idx_0 == 5'h1E;
  wire        _GEN_1773 = lcam_ldq_idx_1 == 5'h1;
  wire        _GEN_1774 = lcam_ldq_idx_1 == 5'h2;
  wire        _GEN_1775 = lcam_ldq_idx_1 == 5'h3;
  wire        _GEN_1776 = lcam_ldq_idx_1 == 5'h4;
  wire        _GEN_1777 = lcam_ldq_idx_1 == 5'h5;
  wire        _GEN_1778 = lcam_ldq_idx_1 == 5'h6;
  wire        _GEN_1779 = lcam_ldq_idx_1 == 5'h7;
  wire        _GEN_1780 = lcam_ldq_idx_1 == 5'h8;
  wire        _GEN_1781 = lcam_ldq_idx_1 == 5'h9;
  wire        _GEN_1782 = lcam_ldq_idx_1 == 5'hA;
  wire        _GEN_1783 = lcam_ldq_idx_1 == 5'hB;
  wire        _GEN_1784 = lcam_ldq_idx_1 == 5'hC;
  wire        _GEN_1785 = lcam_ldq_idx_1 == 5'hD;
  wire        _GEN_1786 = lcam_ldq_idx_1 == 5'hE;
  wire        _GEN_1787 = lcam_ldq_idx_1 == 5'hF;
  wire        _GEN_1788 = lcam_ldq_idx_1 == 5'h10;
  wire        _GEN_1789 = lcam_ldq_idx_1 == 5'h11;
  wire        _GEN_1790 = lcam_ldq_idx_1 == 5'h12;
  wire        _GEN_1791 = lcam_ldq_idx_1 == 5'h13;
  wire        _GEN_1792 = lcam_ldq_idx_1 == 5'h14;
  wire        _GEN_1793 = lcam_ldq_idx_1 == 5'h15;
  wire        _GEN_1794 = lcam_ldq_idx_1 == 5'h16;
  wire        _GEN_1795 = lcam_ldq_idx_1 == 5'h17;
  wire        _GEN_1796 = lcam_ldq_idx_1 == 5'h18;
  wire        _GEN_1797 = lcam_ldq_idx_1 == 5'h19;
  wire        _GEN_1798 = lcam_ldq_idx_1 == 5'h1A;
  wire        _GEN_1799 = lcam_ldq_idx_1 == 5'h1B;
  wire        _GEN_1800 = lcam_ldq_idx_1 == 5'h1C;
  wire        _GEN_1801 = lcam_ldq_idx_1 == 5'h1D;
  wire        _GEN_1802 = lcam_ldq_idx_1 == 5'h1E;
  wire        _GEN_83271 = _GEN_351 ? _GEN_83096 | _GEN_52320 : _GEN_352 & searcher_is_older & _GEN_83098 | _GEN_52320;
  wire        _GEN_83769 = _GEN_370 ? _GEN_83594 | _GEN_52321 : _GEN_371 & searcher_is_older_2 & _GEN_83596 | _GEN_52321;
  wire        _GEN_84267 = _GEN_390 ? _GEN_84092 | _GEN_52322 : _GEN_391 & searcher_is_older_4 & _GEN_84094 | _GEN_52322;
  wire        _GEN_84765 = _GEN_410 ? _GEN_84590 | _GEN_52323 : _GEN_411 & searcher_is_older_6 & _GEN_84592 | _GEN_52323;
  wire        _GEN_85263 = _GEN_430 ? _GEN_85088 | _GEN_52324 : _GEN_431 & searcher_is_older_8 & _GEN_85090 | _GEN_52324;
  wire        _GEN_85761 = _GEN_450 ? _GEN_85586 | _GEN_52325 : _GEN_451 & searcher_is_older_10 & _GEN_85588 | _GEN_52325;
  wire        _GEN_86259 = _GEN_470 ? _GEN_86084 | _GEN_52326 : _GEN_471 & searcher_is_older_12 & _GEN_86086 | _GEN_52326;
  wire        _GEN_86757 = _GEN_490 ? _GEN_86582 | _GEN_52327 : _GEN_491 & searcher_is_older_14 & _GEN_86584 | _GEN_52327;
  wire        _GEN_87255 = _GEN_510 ? _GEN_87080 | _GEN_52328 : _GEN_511 & searcher_is_older_16 & _GEN_87082 | _GEN_52328;
  wire        _GEN_87753 = _GEN_530 ? _GEN_87578 | _GEN_52329 : _GEN_531 & searcher_is_older_18 & _GEN_87580 | _GEN_52329;
  wire        _GEN_88251 = _GEN_550 ? _GEN_88076 | _GEN_52330 : _GEN_551 & searcher_is_older_20 & _GEN_88078 | _GEN_52330;
  wire        _GEN_88749 = _GEN_570 ? _GEN_88574 | _GEN_52331 : _GEN_571 & searcher_is_older_22 & _GEN_88576 | _GEN_52331;
  wire        _GEN_89247 = _GEN_590 ? _GEN_89072 | _GEN_52332 : _GEN_591 & searcher_is_older_24 & _GEN_89074 | _GEN_52332;
  wire        _GEN_89745 = _GEN_610 ? _GEN_89570 | _GEN_52333 : _GEN_611 & searcher_is_older_26 & _GEN_89572 | _GEN_52333;
  wire        _GEN_90243 = _GEN_630 ? _GEN_90068 | _GEN_52334 : _GEN_631 & searcher_is_older_28 & _GEN_90070 | _GEN_52334;
  wire        _GEN_90741 = _GEN_650 ? _GEN_90566 | _GEN_52335 : _GEN_651 & searcher_is_older_30 & _GEN_90568 | _GEN_52335;
  wire        _GEN_91239 = _GEN_670 ? _GEN_91064 | _GEN_52336 : _GEN_671 & searcher_is_older_32 & _GEN_91066 | _GEN_52336;
  wire        _GEN_91737 = _GEN_690 ? _GEN_91562 | _GEN_52337 : _GEN_691 & searcher_is_older_34 & _GEN_91564 | _GEN_52337;
  wire        _GEN_92235 = _GEN_710 ? _GEN_92060 | _GEN_52338 : _GEN_711 & searcher_is_older_36 & _GEN_92062 | _GEN_52338;
  wire        _GEN_92733 = _GEN_730 ? _GEN_92558 | _GEN_52339 : _GEN_731 & searcher_is_older_38 & _GEN_92560 | _GEN_52339;
  wire        _GEN_93231 = _GEN_750 ? _GEN_93056 | _GEN_52340 : _GEN_751 & searcher_is_older_40 & _GEN_93058 | _GEN_52340;
  wire        _GEN_93729 = _GEN_770 ? _GEN_93554 | _GEN_52341 : _GEN_771 & searcher_is_older_42 & _GEN_93556 | _GEN_52341;
  wire        _GEN_94227 = _GEN_790 ? _GEN_94052 | _GEN_52342 : _GEN_791 & searcher_is_older_44 & _GEN_94054 | _GEN_52342;
  wire        _GEN_94725 = _GEN_810 ? _GEN_94550 | _GEN_52343 : _GEN_811 & searcher_is_older_46 & _GEN_94552 | _GEN_52343;
  wire        _GEN_95223 = _GEN_830 ? _GEN_95048 | _GEN_52344 : _GEN_831 & searcher_is_older_48 & _GEN_95050 | _GEN_52344;
  wire        _GEN_95721 = _GEN_850 ? _GEN_95546 | _GEN_52345 : _GEN_851 & searcher_is_older_50 & _GEN_95548 | _GEN_52345;
  wire        _GEN_96219 = _GEN_870 ? _GEN_96044 | _GEN_52346 : _GEN_871 & searcher_is_older_52 & _GEN_96046 | _GEN_52346;
  wire        _GEN_96717 = _GEN_890 ? _GEN_96542 | _GEN_52347 : _GEN_891 & searcher_is_older_54 & _GEN_96544 | _GEN_52347;
  wire        _GEN_97215 = _GEN_910 ? _GEN_97040 | _GEN_52348 : _GEN_911 & searcher_is_older_56 & _GEN_97042 | _GEN_52348;
  wire        _GEN_97713 = _GEN_930 ? _GEN_97538 | _GEN_52349 : _GEN_931 & searcher_is_older_58 & _GEN_97540 | _GEN_52349;
  wire        _GEN_98211 = _GEN_950 ? _GEN_98036 | _GEN_52350 : _GEN_951 & searcher_is_older_60 & _GEN_98038 | _GEN_52350;
  wire        _GEN_1803 =
    (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & (&lcam_ldq_idx_1))) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & (&lcam_ldq_idx_0))) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & (&lcam_ldq_idx_1))) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & (&lcam_ldq_idx_0))) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & (&lcam_ldq_idx_1))) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & (&lcam_ldq_idx_0))) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & (&lcam_ldq_idx_1))) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & (&lcam_ldq_idx_0))) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & (&lcam_ldq_idx_1))) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & (&lcam_ldq_idx_0))) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & (&lcam_ldq_idx_1))) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & (&lcam_ldq_idx_0))) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & (&lcam_ldq_idx_1))) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & (&lcam_ldq_idx_0))) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & (&lcam_ldq_idx_1))) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & (&lcam_ldq_idx_0))) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & (&lcam_ldq_idx_1))) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & (&lcam_ldq_idx_0))) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & (&lcam_ldq_idx_1))) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & (&lcam_ldq_idx_0))) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & (&lcam_ldq_idx_1))) & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & (&lcam_ldq_idx_0)))
    & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & (&lcam_ldq_idx_1))) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & (&lcam_ldq_idx_0))) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & (&lcam_ldq_idx_1))) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & (&lcam_ldq_idx_0))) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & (&lcam_ldq_idx_1))) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & (&lcam_ldq_idx_0))) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & (&lcam_ldq_idx_1))) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & (&lcam_ldq_idx_0))) & (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & (&lcam_ldq_idx_1)));
  wire        _GEN_1804 =
    (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & (&lcam_ldq_idx_0))) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & (&lcam_ldq_idx_1))) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & (&lcam_ldq_idx_0))) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & (&lcam_ldq_idx_1))) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & (&lcam_ldq_idx_0))) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & (&lcam_ldq_idx_1))) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & (&lcam_ldq_idx_0))) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & (&lcam_ldq_idx_1))) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & (&lcam_ldq_idx_0))) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & (&lcam_ldq_idx_1))) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & (&lcam_ldq_idx_0))) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & (&lcam_ldq_idx_1))) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & (&lcam_ldq_idx_0))) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & (&lcam_ldq_idx_1))) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & (&lcam_ldq_idx_0))) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & (&lcam_ldq_idx_1))) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & (&lcam_ldq_idx_0))) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & (&lcam_ldq_idx_1))) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & (&lcam_ldq_idx_0))) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & (&lcam_ldq_idx_1))) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & (&lcam_ldq_idx_0))) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & (&lcam_ldq_idx_1)))
    & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & (&lcam_ldq_idx_0))) & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & (&lcam_ldq_idx_1))) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & (&lcam_ldq_idx_0))) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & (&lcam_ldq_idx_1))) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & (&lcam_ldq_idx_0))) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & (&lcam_ldq_idx_1))) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & (&lcam_ldq_idx_0))) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & (&lcam_ldq_idx_1))) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & (&lcam_ldq_idx_0))) & s1_executing_loads_31;
  wire        _GEN_98530 = _GEN_1803 & _GEN_1804;
  wire        _GEN_98709 = _GEN_970 ? _GEN_98534 | _GEN_52351 : _GEN_971 & searcher_is_older_62 & _GEN_98536 | _GEN_52351;
  wire        _GEN_1805 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & ~(|lcam_ldq_idx_1))) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & ~(|lcam_ldq_idx_0))) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & ~(|lcam_ldq_idx_1))) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & ~(|lcam_ldq_idx_0))) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & ~(|lcam_ldq_idx_1))) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & ~(|lcam_ldq_idx_0))) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & ~(|lcam_ldq_idx_1))) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & ~(|lcam_ldq_idx_0))) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & ~(|lcam_ldq_idx_1))) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & ~(|lcam_ldq_idx_0))) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & ~(|lcam_ldq_idx_1))) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & ~(|lcam_ldq_idx_0))) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & ~(|lcam_ldq_idx_1))) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & ~(|lcam_ldq_idx_0))) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & ~(|lcam_ldq_idx_1))) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & ~(|lcam_ldq_idx_0))) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & ~(|lcam_ldq_idx_1))) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & ~(|lcam_ldq_idx_0))) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & ~(|lcam_ldq_idx_1))) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & ~(|lcam_ldq_idx_0))) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & ~(|lcam_ldq_idx_1)))
    & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & ~(|lcam_ldq_idx_0))) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & ~(|lcam_ldq_idx_1))) & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & ~(|lcam_ldq_idx_0))) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & ~(|lcam_ldq_idx_1))) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & ~(|lcam_ldq_idx_0))) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & ~(|lcam_ldq_idx_1))) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & ~(|lcam_ldq_idx_0))) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & ~(|lcam_ldq_idx_1))) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & ~(|lcam_ldq_idx_0))) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & ~(|lcam_ldq_idx_1)));
  wire        _GEN_1806 =
    (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & ~(|lcam_ldq_idx_0))) & (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & ~(|lcam_ldq_idx_1))) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & ~(|lcam_ldq_idx_0))) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & ~(|lcam_ldq_idx_1))) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & ~(|lcam_ldq_idx_0))) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & ~(|lcam_ldq_idx_1))) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & ~(|lcam_ldq_idx_0))) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & ~(|lcam_ldq_idx_1))) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & ~(|lcam_ldq_idx_0))) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & ~(|lcam_ldq_idx_1))) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & ~(|lcam_ldq_idx_0))) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & ~(|lcam_ldq_idx_1))) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & ~(|lcam_ldq_idx_0))) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & ~(|lcam_ldq_idx_1))) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & ~(|lcam_ldq_idx_0))) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & ~(|lcam_ldq_idx_1))) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & ~(|lcam_ldq_idx_0))) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & ~(|lcam_ldq_idx_1))) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & ~(|lcam_ldq_idx_0))) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & ~(|lcam_ldq_idx_1))) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & ~(|lcam_ldq_idx_0)))
    & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & ~(|lcam_ldq_idx_1))) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & ~(|lcam_ldq_idx_0))) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & ~(|lcam_ldq_idx_1))) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & ~(|lcam_ldq_idx_0))) & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & ~(|lcam_ldq_idx_1))) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & ~(|lcam_ldq_idx_0))) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & ~(|lcam_ldq_idx_1))) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & ~(|lcam_ldq_idx_0))) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & ~(|lcam_ldq_idx_1))) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & ~(|lcam_ldq_idx_0))) & s1_executing_loads_0;
  wire        _GEN_98997 = _GEN_1805 & _GEN_1806;
  wire        _GEN_1807 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1773)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1743)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1773)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1743)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1773)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1743)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1773)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1743)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1773)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1743)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1773)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1743)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1773)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1743)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1773)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1743)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1773)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1743)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1773)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1743)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1773)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1743)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1773))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1743)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1773)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1743)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1773)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1743)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1773)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1743)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1773)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1743));
  wire        _GEN_1808 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1773)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1743)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1773)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1743)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1773)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1743)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1773)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1743)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1773)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1743)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1773)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1743)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1773)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1743)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1773)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1743)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1773)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1743)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1773)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1743)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1773)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1743)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1773)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1743))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1773)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1743)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1773)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1743)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1773)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1743)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1773)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1743)) & s1_executing_loads_1;
  wire        _GEN_98998 = _GEN_1807 & _GEN_1808;
  wire        _GEN_1809 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1774)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1744)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1774)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1744)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1774)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1744)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1774)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1744)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1774)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1744)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1774)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1744)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1774)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1744)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1774)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1744)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1774)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1744)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1774)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1744)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1774)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1744)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1774))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1744)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1774)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1744)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1774)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1744)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1774)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1744)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1774)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1744));
  wire        _GEN_1810 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1774)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1744)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1774)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1744)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1774)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1744)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1774)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1744)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1774)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1744)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1774)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1744)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1774)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1744)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1774)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1744)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1774)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1744)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1774)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1744)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1774)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1744)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1774)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1744))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1774)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1744)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1774)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1744)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1774)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1744)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1774)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1744)) & s1_executing_loads_2;
  wire        _GEN_98999 = _GEN_1809 & _GEN_1810;
  wire        _GEN_1811 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1775)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1745)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1775)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1745)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1775)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1745)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1775)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1745)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1775)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1745)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1775)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1745)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1775)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1745)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1775)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1745)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1775)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1745)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1775)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1745)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1775)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1745)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1775))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1745)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1775)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1745)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1775)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1745)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1775)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1745)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1775)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1745));
  wire        _GEN_1812 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1775)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1745)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1775)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1745)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1775)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1745)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1775)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1745)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1775)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1745)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1775)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1745)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1775)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1745)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1775)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1745)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1775)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1745)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1775)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1745)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1775)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1745)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1775)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1745))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1775)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1745)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1775)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1745)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1775)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1745)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1775)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1745)) & s1_executing_loads_3;
  wire        _GEN_99000 = _GEN_1811 & _GEN_1812;
  wire        _GEN_1813 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1776)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1746)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1776)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1746)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1776)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1746)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1776)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1746)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1776)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1746)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1776)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1746)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1776)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1746)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1776)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1746)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1776)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1746)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1776)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1746)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1776)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1746)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1776))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1746)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1776)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1746)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1776)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1746)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1776)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1746)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1776)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1746));
  wire        _GEN_1814 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1776)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1746)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1776)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1746)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1776)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1746)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1776)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1746)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1776)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1746)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1776)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1746)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1776)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1746)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1776)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1746)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1776)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1746)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1776)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1746)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1776)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1746)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1776)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1746))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1776)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1746)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1776)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1746)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1776)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1746)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1776)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1746)) & s1_executing_loads_4;
  wire        _GEN_99001 = _GEN_1813 & _GEN_1814;
  wire        _GEN_1815 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1777)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1747)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1777)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1747)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1777)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1747)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1777)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1747)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1777)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1747)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1777)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1747)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1777)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1747)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1777)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1747)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1777)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1747)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1777)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1747)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1777)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1747)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1777))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1747)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1777)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1747)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1777)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1747)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1777)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1747)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1777)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1747));
  wire        _GEN_1816 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1777)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1747)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1777)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1747)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1777)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1747)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1777)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1747)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1777)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1747)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1777)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1747)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1777)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1747)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1777)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1747)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1777)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1747)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1777)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1747)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1777)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1747)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1777)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1747))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1777)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1747)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1777)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1747)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1777)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1747)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1777)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1747)) & s1_executing_loads_5;
  wire        _GEN_99002 = _GEN_1815 & _GEN_1816;
  wire        _GEN_1817 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1778)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1748)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1778)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1748)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1778)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1748)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1778)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1748)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1778)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1748)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1778)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1748)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1778)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1748)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1778)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1748)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1778)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1748)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1778)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1748)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1778)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1748)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1778))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1748)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1778)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1748)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1778)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1748)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1778)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1748)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1778)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1748));
  wire        _GEN_1818 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1778)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1748)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1778)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1748)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1778)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1748)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1778)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1748)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1778)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1748)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1778)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1748)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1778)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1748)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1778)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1748)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1778)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1748)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1778)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1748)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1778)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1748)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1778)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1748))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1778)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1748)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1778)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1748)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1778)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1748)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1778)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1748)) & s1_executing_loads_6;
  wire        _GEN_99003 = _GEN_1817 & _GEN_1818;
  wire        _GEN_1819 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1779)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1749)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1779)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1749)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1779)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1749)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1779)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1749)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1779)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1749)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1779)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1749)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1779)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1749)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1779)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1749)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1779)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1749)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1779)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1749)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1779)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1749)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1779))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1749)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1779)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1749)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1779)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1749)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1779)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1749)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1779)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1749));
  wire        _GEN_1820 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1779)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1749)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1779)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1749)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1779)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1749)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1779)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1749)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1779)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1749)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1779)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1749)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1779)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1749)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1779)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1749)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1779)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1749)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1779)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1749)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1779)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1749)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1779)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1749))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1779)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1749)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1779)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1749)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1779)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1749)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1779)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1749)) & s1_executing_loads_7;
  wire        _GEN_99004 = _GEN_1819 & _GEN_1820;
  wire        _GEN_1821 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1780)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1750)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1780)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1750)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1780)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1750)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1780)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1750)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1780)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1750)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1780)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1750)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1780)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1750)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1780)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1750)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1780)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1750)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1780)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1750)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1780)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1750)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1780))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1750)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1780)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1750)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1780)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1750)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1780)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1750)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1780)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1750));
  wire        _GEN_1822 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1780)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1750)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1780)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1750)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1780)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1750)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1780)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1750)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1780)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1750)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1780)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1750)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1780)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1750)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1780)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1750)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1780)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1750)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1780)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1750)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1780)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1750)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1780)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1750))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1780)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1750)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1780)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1750)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1780)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1750)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1780)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1750)) & s1_executing_loads_8;
  wire        _GEN_99005 = _GEN_1821 & _GEN_1822;
  wire        _GEN_1823 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1781)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1751)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1781)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1751)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1781)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1751)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1781)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1751)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1781)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1751)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1781)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1751)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1781)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1751)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1781)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1751)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1781)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1751)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1781)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1751)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1781)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1751)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1781))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1751)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1781)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1751)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1781)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1751)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1781)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1751)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1781)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1751));
  wire        _GEN_1824 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1781)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1751)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1781)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1751)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1781)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1751)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1781)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1751)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1781)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1751)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1781)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1751)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1781)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1751)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1781)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1751)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1781)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1751)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1781)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1751)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1781)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1751)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1781)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1751))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1781)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1751)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1781)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1751)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1781)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1751)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1781)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1751)) & s1_executing_loads_9;
  wire        _GEN_99006 = _GEN_1823 & _GEN_1824;
  wire        _GEN_1825 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1782)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1752)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1782)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1752)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1782)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1752)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1782)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1752)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1782)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1752)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1782)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1752)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1782)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1752)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1782)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1752)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1782)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1752)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1782)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1752)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1782)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1752)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1782))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1752)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1782)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1752)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1782)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1752)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1782)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1752)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1782)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1752));
  wire        _GEN_1826 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1782)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1752)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1782)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1752)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1782)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1752)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1782)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1752)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1782)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1752)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1782)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1752)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1782)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1752)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1782)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1752)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1782)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1752)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1782)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1752)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1782)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1752)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1782)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1752))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1782)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1752)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1782)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1752)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1782)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1752)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1782)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1752)) & s1_executing_loads_10;
  wire        _GEN_99007 = _GEN_1825 & _GEN_1826;
  wire        _GEN_1827 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1783)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1753)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1783)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1753)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1783)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1753)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1783)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1753)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1783)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1753)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1783)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1753)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1783)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1753)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1783)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1753)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1783)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1753)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1783)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1753)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1783)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1753)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1783))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1753)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1783)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1753)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1783)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1753)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1783)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1753)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1783)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1753));
  wire        _GEN_1828 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1783)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1753)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1783)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1753)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1783)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1753)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1783)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1753)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1783)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1753)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1783)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1753)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1783)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1753)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1783)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1753)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1783)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1753)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1783)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1753)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1783)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1753)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1783)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1753))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1783)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1753)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1783)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1753)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1783)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1753)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1783)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1753)) & s1_executing_loads_11;
  wire        _GEN_99008 = _GEN_1827 & _GEN_1828;
  wire        _GEN_1829 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1784)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1754)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1784)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1754)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1784)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1754)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1784)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1754)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1784)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1754)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1784)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1754)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1784)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1754)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1784)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1754)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1784)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1754)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1784)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1754)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1784)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1754)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1784))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1754)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1784)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1754)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1784)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1754)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1784)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1754)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1784)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1754));
  wire        _GEN_1830 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1784)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1754)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1784)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1754)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1784)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1754)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1784)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1754)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1784)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1754)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1784)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1754)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1784)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1754)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1784)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1754)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1784)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1754)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1784)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1754)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1784)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1754)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1784)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1754))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1784)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1754)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1784)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1754)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1784)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1754)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1784)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1754)) & s1_executing_loads_12;
  wire        _GEN_99009 = _GEN_1829 & _GEN_1830;
  wire        _GEN_1831 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1785)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1755)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1785)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1755)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1785)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1755)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1785)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1755)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1785)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1755)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1785)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1755)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1785)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1755)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1785)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1755)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1785)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1755)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1785)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1755)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1785)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1755)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1785))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1755)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1785)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1755)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1785)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1755)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1785)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1755)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1785)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1755));
  wire        _GEN_1832 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1785)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1755)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1785)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1755)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1785)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1755)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1785)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1755)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1785)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1755)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1785)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1755)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1785)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1755)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1785)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1755)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1785)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1755)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1785)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1755)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1785)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1755)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1785)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1755))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1785)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1755)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1785)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1755)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1785)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1755)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1785)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1755)) & s1_executing_loads_13;
  wire        _GEN_99010 = _GEN_1831 & _GEN_1832;
  wire        _GEN_1833 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1786)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1756)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1786)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1756)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1786)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1756)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1786)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1756)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1786)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1756)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1786)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1756)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1786)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1756)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1786)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1756)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1786)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1756)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1786)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1756)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1786)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1756)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1786))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1756)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1786)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1756)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1786)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1756)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1786)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1756)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1786)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1756));
  wire        _GEN_1834 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1786)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1756)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1786)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1756)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1786)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1756)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1786)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1756)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1786)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1756)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1786)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1756)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1786)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1756)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1786)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1756)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1786)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1756)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1786)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1756)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1786)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1756)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1786)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1756))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1786)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1756)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1786)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1756)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1786)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1756)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1786)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1756)) & s1_executing_loads_14;
  wire        _GEN_99011 = _GEN_1833 & _GEN_1834;
  wire        _GEN_1835 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1787)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1757)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1787)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1757)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1787)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1757)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1787)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1757)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1787)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1757)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1787)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1757)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1787)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1757)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1787)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1757)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1787)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1757)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1787)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1757)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1787)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1757)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1787))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1757)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1787)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1757)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1787)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1757)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1787)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1757)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1787)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1757));
  wire        _GEN_1836 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1787)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1757)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1787)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1757)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1787)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1757)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1787)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1757)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1787)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1757)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1787)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1757)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1787)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1757)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1787)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1757)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1787)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1757)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1787)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1757)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1787)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1757)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1787)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1757))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1787)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1757)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1787)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1757)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1787)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1757)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1787)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1757)) & s1_executing_loads_15;
  wire        _GEN_99012 = _GEN_1835 & _GEN_1836;
  wire        _GEN_1837 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1788)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1758)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1788)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1758)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1788)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1758)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1788)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1758)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1788)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1758)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1788)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1758)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1788)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1758)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1788)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1758)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1788)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1758)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1788)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1758)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1788)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1758)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1788))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1758)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1788)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1758)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1788)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1758)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1788)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1758)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1788)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1758));
  wire        _GEN_1838 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1788)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1758)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1788)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1758)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1788)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1758)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1788)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1758)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1788)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1758)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1788)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1758)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1788)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1758)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1788)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1758)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1788)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1758)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1788)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1758)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1788)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1758)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1788)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1758))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1788)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1758)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1788)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1758)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1788)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1758)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1788)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1758)) & s1_executing_loads_16;
  wire        _GEN_99013 = _GEN_1837 & _GEN_1838;
  wire        _GEN_1839 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1789)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1759)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1789)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1759)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1789)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1759)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1789)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1759)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1789)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1759)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1789)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1759)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1789)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1759)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1789)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1759)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1789)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1759)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1789)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1759)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1789)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1759)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1789))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1759)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1789)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1759)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1789)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1759)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1789)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1759)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1789)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1759));
  wire        _GEN_1840 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1789)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1759)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1789)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1759)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1789)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1759)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1789)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1759)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1789)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1759)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1789)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1759)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1789)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1759)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1789)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1759)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1789)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1759)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1789)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1759)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1789)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1759)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1789)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1759))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1789)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1759)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1789)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1759)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1789)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1759)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1789)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1759)) & s1_executing_loads_17;
  wire        _GEN_99014 = _GEN_1839 & _GEN_1840;
  wire        _GEN_1841 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1790)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1760)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1790)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1760)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1790)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1760)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1790)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1760)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1790)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1760)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1790)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1760)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1790)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1760)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1790)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1760)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1790)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1760)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1790)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1760)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1790)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1760)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1790))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1760)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1790)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1760)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1790)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1760)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1790)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1760)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1790)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1760));
  wire        _GEN_1842 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1790)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1760)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1790)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1760)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1790)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1760)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1790)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1760)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1790)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1760)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1790)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1760)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1790)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1760)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1790)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1760)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1790)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1760)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1790)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1760)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1790)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1760)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1790)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1760))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1790)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1760)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1790)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1760)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1790)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1760)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1790)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1760)) & s1_executing_loads_18;
  wire        _GEN_99015 = _GEN_1841 & _GEN_1842;
  wire        _GEN_1843 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1791)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1761)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1791)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1761)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1791)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1761)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1791)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1761)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1791)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1761)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1791)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1761)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1791)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1761)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1791)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1761)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1791)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1761)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1791)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1761)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1791)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1761)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1791))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1761)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1791)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1761)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1791)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1761)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1791)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1761)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1791)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1761));
  wire        _GEN_1844 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1791)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1761)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1791)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1761)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1791)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1761)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1791)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1761)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1791)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1761)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1791)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1761)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1791)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1761)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1791)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1761)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1791)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1761)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1791)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1761)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1791)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1761)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1791)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1761))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1791)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1761)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1791)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1761)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1791)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1761)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1791)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1761)) & s1_executing_loads_19;
  wire        _GEN_99016 = _GEN_1843 & _GEN_1844;
  wire        _GEN_1845 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1792)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1762)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1792)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1762)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1792)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1762)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1792)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1762)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1792)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1762)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1792)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1762)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1792)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1762)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1792)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1762)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1792)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1762)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1792)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1762)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1792)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1762)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1792))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1762)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1792)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1762)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1792)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1762)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1792)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1762)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1792)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1762));
  wire        _GEN_1846 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1792)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1762)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1792)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1762)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1792)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1762)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1792)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1762)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1792)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1762)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1792)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1762)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1792)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1762)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1792)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1762)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1792)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1762)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1792)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1762)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1792)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1762)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1792)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1762))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1792)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1762)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1792)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1762)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1792)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1762)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1792)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1762)) & s1_executing_loads_20;
  wire        _GEN_99017 = _GEN_1845 & _GEN_1846;
  wire        _GEN_1847 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1793)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1763)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1793)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1763)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1793)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1763)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1793)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1763)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1793)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1763)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1793)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1763)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1793)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1763)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1793)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1763)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1793)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1763)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1793)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1763)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1793)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1763)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1793))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1763)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1793)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1763)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1793)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1763)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1793)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1763)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1793)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1763));
  wire        _GEN_1848 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1793)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1763)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1793)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1763)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1793)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1763)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1793)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1763)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1793)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1763)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1793)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1763)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1793)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1763)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1793)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1763)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1793)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1763)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1793)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1763)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1793)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1763)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1793)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1763))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1793)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1763)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1793)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1763)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1793)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1763)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1793)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1763)) & s1_executing_loads_21;
  wire        _GEN_99018 = _GEN_1847 & _GEN_1848;
  wire        _GEN_1849 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1794)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1764)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1794)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1764)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1794)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1764)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1794)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1764)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1794)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1764)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1794)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1764)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1794)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1764)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1794)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1764)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1794)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1764)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1794)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1764)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1794)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1764)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1794))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1764)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1794)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1764)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1794)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1764)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1794)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1764)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1794)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1764));
  wire        _GEN_1850 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1794)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1764)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1794)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1764)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1794)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1764)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1794)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1764)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1794)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1764)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1794)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1764)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1794)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1764)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1794)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1764)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1794)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1764)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1794)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1764)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1794)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1764)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1794)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1764))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1794)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1764)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1794)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1764)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1794)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1764)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1794)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1764)) & s1_executing_loads_22;
  wire        _GEN_99019 = _GEN_1849 & _GEN_1850;
  wire        _GEN_1851 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1795)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1765)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1795)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1765)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1795)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1765)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1795)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1765)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1795)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1765)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1795)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1765)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1795)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1765)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1795)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1765)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1795)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1765)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1795)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1765)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1795)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1765)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1795))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1765)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1795)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1765)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1795)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1765)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1795)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1765)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1795)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1765));
  wire        _GEN_1852 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1795)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1765)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1795)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1765)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1795)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1765)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1795)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1765)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1795)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1765)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1795)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1765)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1795)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1765)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1795)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1765)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1795)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1765)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1795)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1765)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1795)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1765)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1795)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1765))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1795)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1765)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1795)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1765)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1795)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1765)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1795)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1765)) & s1_executing_loads_23;
  wire        _GEN_99020 = _GEN_1851 & _GEN_1852;
  wire        _GEN_1853 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1796)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1766)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1796)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1766)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1796)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1766)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1796)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1766)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1796)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1766)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1796)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1766)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1796)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1766)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1796)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1766)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1796)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1766)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1796)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1766)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1796)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1766)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1796))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1766)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1796)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1766)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1796)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1766)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1796)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1766)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1796)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1766));
  wire        _GEN_1854 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1796)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1766)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1796)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1766)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1796)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1766)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1796)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1766)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1796)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1766)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1796)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1766)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1796)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1766)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1796)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1766)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1796)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1766)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1796)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1766)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1796)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1766)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1796)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1766))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1796)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1766)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1796)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1766)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1796)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1766)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1796)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1766)) & s1_executing_loads_24;
  wire        _GEN_99021 = _GEN_1853 & _GEN_1854;
  wire        _GEN_1855 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1797)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1767)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1797)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1767)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1797)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1767)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1797)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1767)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1797)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1767)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1797)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1767)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1797)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1767)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1797)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1767)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1797)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1767)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1797)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1767)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1797)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1767)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1797))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1767)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1797)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1767)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1797)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1767)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1797)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1767)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1797)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1767));
  wire        _GEN_1856 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1797)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1767)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1797)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1767)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1797)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1767)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1797)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1767)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1797)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1767)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1797)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1767)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1797)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1767)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1797)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1767)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1797)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1767)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1797)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1767)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1797)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1767)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1797)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1767))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1797)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1767)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1797)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1767)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1797)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1767)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1797)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1767)) & s1_executing_loads_25;
  wire        _GEN_99022 = _GEN_1855 & _GEN_1856;
  wire        _GEN_1857 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1798)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1768)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1798)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1768)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1798)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1768)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1798)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1768)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1798)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1768)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1798)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1768)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1798)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1768)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1798)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1768)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1798)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1768)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1798)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1768)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1798)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1768)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1798))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1768)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1798)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1768)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1798)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1768)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1798)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1768)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1798)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1768));
  wire        _GEN_1858 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1798)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1768)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1798)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1768)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1798)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1768)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1798)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1768)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1798)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1768)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1798)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1768)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1798)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1768)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1798)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1768)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1798)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1768)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1798)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1768)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1798)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1768)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1798)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1768))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1798)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1768)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1798)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1768)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1798)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1768)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1798)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1768)) & s1_executing_loads_26;
  wire        _GEN_99023 = _GEN_1857 & _GEN_1858;
  wire        _GEN_1859 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1799)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1769)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1799)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1769)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1799)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1769)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1799)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1769)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1799)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1769)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1799)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1769)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1799)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1769)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1799)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1769)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1799)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1769)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1799)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1769)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1799)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1769)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1799))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1769)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1799)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1769)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1799)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1769)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1799)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1769)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1799)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1769));
  wire        _GEN_1860 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1799)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1769)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1799)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1769)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1799)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1769)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1799)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1769)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1799)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1769)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1799)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1769)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1799)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1769)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1799)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1769)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1799)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1769)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1799)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1769)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1799)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1769)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1799)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1769))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1799)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1769)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1799)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1769)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1799)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1769)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1799)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1769)) & s1_executing_loads_27;
  wire        _GEN_99024 = _GEN_1859 & _GEN_1860;
  wire        _GEN_1861 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1800)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1770)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1800)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1770)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1800)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1770)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1800)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1770)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1800)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1770)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1800)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1770)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1800)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1770)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1800)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1770)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1800)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1770)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1800)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1770)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1800)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1770)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1800))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1770)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1800)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1770)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1800)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1770)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1800)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1770)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1800)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1770));
  wire        _GEN_1862 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1800)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1770)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1800)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1770)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1800)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1770)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1800)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1770)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1800)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1770)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1800)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1770)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1800)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1770)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1800)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1770)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1800)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1770)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1800)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1770)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1800)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1770)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1800)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1770))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1800)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1770)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1800)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1770)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1800)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1770)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1800)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1770)) & s1_executing_loads_28;
  wire        _GEN_99025 = _GEN_1861 & _GEN_1862;
  wire        _GEN_1863 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1801)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1771)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1801)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1771)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1801)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1771)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1801)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1771)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1801)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1771)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1801)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1771)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1801)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1771)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1801)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1771)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1801)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1771)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1801)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1771)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1801)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1771)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1801))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1771)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1801)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1771)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1801)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1771)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1801)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1771)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1801)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1771));
  wire        _GEN_1864 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1801)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1771)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1801)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1771)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1801)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1771)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1801)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1771)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1801)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1771)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1801)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1771)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1801)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1771)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1801)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1771)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1801)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1771)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1801)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1771)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1801)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1771)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1801)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1771))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1801)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1771)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1801)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1771)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1801)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1771)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1801)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1771)) & s1_executing_loads_29;
  wire        _GEN_99026 = _GEN_1863 & _GEN_1864;
  wire        _GEN_1865 =
    (_GEN_983 | ~_GEN_980 | searcher_is_older_63 | ~(~(&lcam_ldq_idx_1) & _GEN_981 & _GEN_1802)) & (_GEN_970 | ~_GEN_971 | searcher_is_older_62 | ~(~(&lcam_ldq_idx_0) & _GEN_974 & _GEN_1772)) & (_GEN_965 | ~_GEN_961 | searcher_is_older_61 | ~(_GEN_962 & _GEN_963 & _GEN_1802)) & (_GEN_950 | ~_GEN_951 | searcher_is_older_60 | ~(_GEN_953 & _GEN_955 & _GEN_1772)) & (_GEN_945 | ~_GEN_941 | searcher_is_older_59 | ~(_GEN_942 & _GEN_943 & _GEN_1802)) & (_GEN_930 | ~_GEN_931 | searcher_is_older_58 | ~(_GEN_933 & _GEN_935 & _GEN_1772)) & (_GEN_925 | ~_GEN_921 | searcher_is_older_57 | ~(_GEN_922 & _GEN_923 & _GEN_1802)) & (_GEN_910 | ~_GEN_911 | searcher_is_older_56 | ~(_GEN_913 & _GEN_915 & _GEN_1772)) & (_GEN_905 | ~_GEN_901 | searcher_is_older_55 | ~(_GEN_902 & _GEN_903 & _GEN_1802)) & (_GEN_890 | ~_GEN_891 | searcher_is_older_54 | ~(_GEN_893 & _GEN_895 & _GEN_1772)) & (_GEN_885 | ~_GEN_881 | searcher_is_older_53 | ~(_GEN_882 & _GEN_883 & _GEN_1802)) & (_GEN_870 | ~_GEN_871 | searcher_is_older_52 | ~(_GEN_873 & _GEN_875 & _GEN_1772)) & (_GEN_865 | ~_GEN_861 | searcher_is_older_51 | ~(_GEN_862 & _GEN_863 & _GEN_1802)) & (_GEN_850 | ~_GEN_851 | searcher_is_older_50 | ~(_GEN_853 & _GEN_855 & _GEN_1772)) & (_GEN_845 | ~_GEN_841 | searcher_is_older_49 | ~(_GEN_842 & _GEN_843 & _GEN_1802)) & (_GEN_830 | ~_GEN_831 | searcher_is_older_48 | ~(_GEN_833 & _GEN_835 & _GEN_1772)) & (_GEN_825 | ~_GEN_821 | searcher_is_older_47 | ~(_GEN_822 & _GEN_823 & _GEN_1802)) & (_GEN_810 | ~_GEN_811 | searcher_is_older_46 | ~(_GEN_813 & _GEN_815 & _GEN_1772)) & (_GEN_805 | ~_GEN_801 | searcher_is_older_45 | ~(_GEN_802 & _GEN_803 & _GEN_1802)) & (_GEN_790 | ~_GEN_791 | searcher_is_older_44 | ~(_GEN_793 & _GEN_795 & _GEN_1772)) & (_GEN_785 | ~_GEN_781 | searcher_is_older_43 | ~(_GEN_782 & _GEN_783 & _GEN_1802)) & (_GEN_770 | ~_GEN_771 | searcher_is_older_42 | ~(_GEN_773 & _GEN_775 & _GEN_1772)) & (_GEN_765 | ~_GEN_761 | searcher_is_older_41 | ~(_GEN_762 & _GEN_763 & _GEN_1802))
    & (_GEN_750 | ~_GEN_751 | searcher_is_older_40 | ~(_GEN_753 & _GEN_755 & _GEN_1772)) & (_GEN_745 | ~_GEN_741 | searcher_is_older_39 | ~(_GEN_742 & _GEN_743 & _GEN_1802)) & (_GEN_730 | ~_GEN_731 | searcher_is_older_38 | ~(_GEN_733 & _GEN_735 & _GEN_1772)) & (_GEN_725 | ~_GEN_721 | searcher_is_older_37 | ~(_GEN_722 & _GEN_723 & _GEN_1802)) & (_GEN_710 | ~_GEN_711 | searcher_is_older_36 | ~(_GEN_713 & _GEN_715 & _GEN_1772)) & (_GEN_705 | ~_GEN_701 | searcher_is_older_35 | ~(_GEN_702 & _GEN_703 & _GEN_1802)) & (_GEN_690 | ~_GEN_691 | searcher_is_older_34 | ~(_GEN_693 & _GEN_695 & _GEN_1772)) & (_GEN_685 | ~_GEN_681 | searcher_is_older_33 | ~(_GEN_682 & _GEN_683 & _GEN_1802)) & (_GEN_670 | ~_GEN_671 | searcher_is_older_32 | ~(_GEN_673 & _GEN_675 & _GEN_1772));
  wire        _GEN_1866 =
    (_GEN_665 | ~_GEN_661 | searcher_is_older_31 | ~(_GEN_662 & _GEN_663 & _GEN_1802)) & (_GEN_650 | ~_GEN_651 | searcher_is_older_30 | ~(_GEN_653 & _GEN_655 & _GEN_1772)) & (_GEN_645 | ~_GEN_641 | searcher_is_older_29 | ~(_GEN_642 & _GEN_643 & _GEN_1802)) & (_GEN_630 | ~_GEN_631 | searcher_is_older_28 | ~(_GEN_633 & _GEN_635 & _GEN_1772)) & (_GEN_625 | ~_GEN_621 | searcher_is_older_27 | ~(_GEN_622 & _GEN_623 & _GEN_1802)) & (_GEN_610 | ~_GEN_611 | searcher_is_older_26 | ~(_GEN_613 & _GEN_615 & _GEN_1772)) & (_GEN_605 | ~_GEN_601 | searcher_is_older_25 | ~(_GEN_602 & _GEN_603 & _GEN_1802)) & (_GEN_590 | ~_GEN_591 | searcher_is_older_24 | ~(_GEN_593 & _GEN_595 & _GEN_1772)) & (_GEN_585 | ~_GEN_581 | searcher_is_older_23 | ~(_GEN_582 & _GEN_583 & _GEN_1802)) & (_GEN_570 | ~_GEN_571 | searcher_is_older_22 | ~(_GEN_573 & _GEN_575 & _GEN_1772)) & (_GEN_565 | ~_GEN_561 | searcher_is_older_21 | ~(_GEN_562 & _GEN_563 & _GEN_1802)) & (_GEN_550 | ~_GEN_551 | searcher_is_older_20 | ~(_GEN_553 & _GEN_555 & _GEN_1772)) & (_GEN_545 | ~_GEN_541 | searcher_is_older_19 | ~(_GEN_542 & _GEN_543 & _GEN_1802)) & (_GEN_530 | ~_GEN_531 | searcher_is_older_18 | ~(_GEN_533 & _GEN_535 & _GEN_1772)) & (_GEN_525 | ~_GEN_521 | searcher_is_older_17 | ~(_GEN_522 & _GEN_523 & _GEN_1802)) & (_GEN_510 | ~_GEN_511 | searcher_is_older_16 | ~(_GEN_513 & _GEN_515 & _GEN_1772)) & (_GEN_505 | ~_GEN_501 | searcher_is_older_15 | ~(_GEN_502 & _GEN_503 & _GEN_1802)) & (_GEN_490 | ~_GEN_491 | searcher_is_older_14 | ~(_GEN_493 & _GEN_495 & _GEN_1772)) & (_GEN_485 | ~_GEN_481 | searcher_is_older_13 | ~(_GEN_482 & _GEN_483 & _GEN_1802)) & (_GEN_470 | ~_GEN_471 | searcher_is_older_12 | ~(_GEN_473 & _GEN_475 & _GEN_1772)) & (_GEN_465 | ~_GEN_461 | searcher_is_older_11 | ~(_GEN_462 & _GEN_463 & _GEN_1802)) & (_GEN_450 | ~_GEN_451 | searcher_is_older_10 | ~(_GEN_453 & _GEN_455 & _GEN_1772)) & (_GEN_445 | ~_GEN_441 | searcher_is_older_9 | ~(_GEN_442 & _GEN_443 & _GEN_1802)) & (_GEN_430 | ~_GEN_431 | searcher_is_older_8 | ~(_GEN_433 & _GEN_435 & _GEN_1772))
    & (_GEN_425 | ~_GEN_421 | searcher_is_older_7 | ~(_GEN_422 & _GEN_423 & _GEN_1802)) & (_GEN_410 | ~_GEN_411 | searcher_is_older_6 | ~(_GEN_413 & _GEN_415 & _GEN_1772)) & (_GEN_405 | ~_GEN_401 | searcher_is_older_5 | ~(_GEN_402 & _GEN_403 & _GEN_1802)) & (_GEN_390 | ~_GEN_391 | searcher_is_older_4 | ~(_GEN_393 & _GEN_395 & _GEN_1772)) & (_GEN_385 | ~_GEN_381 | searcher_is_older_3 | ~(_GEN_382 & _GEN_383 & _GEN_1802)) & (_GEN_370 | ~_GEN_371 | searcher_is_older_2 | ~(_GEN_373 & _GEN_375 & _GEN_1772)) & (_GEN_366 | ~_GEN_362 | searcher_is_older_1 | ~((|lcam_ldq_idx_1) & _GEN_363 & _GEN_1802)) & (_GEN_351 | ~_GEN_352 | searcher_is_older | ~((|lcam_ldq_idx_0) & _GEN_355 & _GEN_1772)) & s1_executing_loads_30;
  wire        _GEN_99027 = _GEN_1865 & _GEN_1866;
  wire        _GEN_99233 = _GEN_985 ? (_GEN_99196 ? (|lcam_ldq_idx_0) & _GEN_98997 : _GEN_987 ? (|lcam_ldq_idx_0) & _GEN_98997 : ~(_GEN_99361 & ~(|lcam_ldq_idx_0)) & _GEN_98997) : _GEN_98997;
  wire        _GEN_99234 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1743 & _GEN_98998 : _GEN_987 ? ~_GEN_1743 & _GEN_98998 : ~(_GEN_99361 & _GEN_1743) & _GEN_98998) : _GEN_98998;
  wire        _GEN_99235 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1744 & _GEN_98999 : _GEN_987 ? ~_GEN_1744 & _GEN_98999 : ~(_GEN_99361 & _GEN_1744) & _GEN_98999) : _GEN_98999;
  wire        _GEN_99236 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1745 & _GEN_99000 : _GEN_987 ? ~_GEN_1745 & _GEN_99000 : ~(_GEN_99361 & _GEN_1745) & _GEN_99000) : _GEN_99000;
  wire        _GEN_99237 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1746 & _GEN_99001 : _GEN_987 ? ~_GEN_1746 & _GEN_99001 : ~(_GEN_99361 & _GEN_1746) & _GEN_99001) : _GEN_99001;
  wire        _GEN_99238 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1747 & _GEN_99002 : _GEN_987 ? ~_GEN_1747 & _GEN_99002 : ~(_GEN_99361 & _GEN_1747) & _GEN_99002) : _GEN_99002;
  wire        _GEN_99239 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1748 & _GEN_99003 : _GEN_987 ? ~_GEN_1748 & _GEN_99003 : ~(_GEN_99361 & _GEN_1748) & _GEN_99003) : _GEN_99003;
  wire        _GEN_99240 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1749 & _GEN_99004 : _GEN_987 ? ~_GEN_1749 & _GEN_99004 : ~(_GEN_99361 & _GEN_1749) & _GEN_99004) : _GEN_99004;
  wire        _GEN_99241 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1750 & _GEN_99005 : _GEN_987 ? ~_GEN_1750 & _GEN_99005 : ~(_GEN_99361 & _GEN_1750) & _GEN_99005) : _GEN_99005;
  wire        _GEN_99242 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1751 & _GEN_99006 : _GEN_987 ? ~_GEN_1751 & _GEN_99006 : ~(_GEN_99361 & _GEN_1751) & _GEN_99006) : _GEN_99006;
  wire        _GEN_99243 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1752 & _GEN_99007 : _GEN_987 ? ~_GEN_1752 & _GEN_99007 : ~(_GEN_99361 & _GEN_1752) & _GEN_99007) : _GEN_99007;
  wire        _GEN_99244 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1753 & _GEN_99008 : _GEN_987 ? ~_GEN_1753 & _GEN_99008 : ~(_GEN_99361 & _GEN_1753) & _GEN_99008) : _GEN_99008;
  wire        _GEN_99245 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1754 & _GEN_99009 : _GEN_987 ? ~_GEN_1754 & _GEN_99009 : ~(_GEN_99361 & _GEN_1754) & _GEN_99009) : _GEN_99009;
  wire        _GEN_99246 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1755 & _GEN_99010 : _GEN_987 ? ~_GEN_1755 & _GEN_99010 : ~(_GEN_99361 & _GEN_1755) & _GEN_99010) : _GEN_99010;
  wire        _GEN_99247 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1756 & _GEN_99011 : _GEN_987 ? ~_GEN_1756 & _GEN_99011 : ~(_GEN_99361 & _GEN_1756) & _GEN_99011) : _GEN_99011;
  wire        _GEN_99248 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1757 & _GEN_99012 : _GEN_987 ? ~_GEN_1757 & _GEN_99012 : ~(_GEN_99361 & _GEN_1757) & _GEN_99012) : _GEN_99012;
  wire        _GEN_99249 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1758 & _GEN_99013 : _GEN_987 ? ~_GEN_1758 & _GEN_99013 : ~(_GEN_99361 & _GEN_1758) & _GEN_99013) : _GEN_99013;
  wire        _GEN_99250 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1759 & _GEN_99014 : _GEN_987 ? ~_GEN_1759 & _GEN_99014 : ~(_GEN_99361 & _GEN_1759) & _GEN_99014) : _GEN_99014;
  wire        _GEN_99251 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1760 & _GEN_99015 : _GEN_987 ? ~_GEN_1760 & _GEN_99015 : ~(_GEN_99361 & _GEN_1760) & _GEN_99015) : _GEN_99015;
  wire        _GEN_99252 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1761 & _GEN_99016 : _GEN_987 ? ~_GEN_1761 & _GEN_99016 : ~(_GEN_99361 & _GEN_1761) & _GEN_99016) : _GEN_99016;
  wire        _GEN_99253 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1762 & _GEN_99017 : _GEN_987 ? ~_GEN_1762 & _GEN_99017 : ~(_GEN_99361 & _GEN_1762) & _GEN_99017) : _GEN_99017;
  wire        _GEN_99254 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1763 & _GEN_99018 : _GEN_987 ? ~_GEN_1763 & _GEN_99018 : ~(_GEN_99361 & _GEN_1763) & _GEN_99018) : _GEN_99018;
  wire        _GEN_99255 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1764 & _GEN_99019 : _GEN_987 ? ~_GEN_1764 & _GEN_99019 : ~(_GEN_99361 & _GEN_1764) & _GEN_99019) : _GEN_99019;
  wire        _GEN_99256 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1765 & _GEN_99020 : _GEN_987 ? ~_GEN_1765 & _GEN_99020 : ~(_GEN_99361 & _GEN_1765) & _GEN_99020) : _GEN_99020;
  wire        _GEN_99257 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1766 & _GEN_99021 : _GEN_987 ? ~_GEN_1766 & _GEN_99021 : ~(_GEN_99361 & _GEN_1766) & _GEN_99021) : _GEN_99021;
  wire        _GEN_99258 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1767 & _GEN_99022 : _GEN_987 ? ~_GEN_1767 & _GEN_99022 : ~(_GEN_99361 & _GEN_1767) & _GEN_99022) : _GEN_99022;
  wire        _GEN_99259 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1768 & _GEN_99023 : _GEN_987 ? ~_GEN_1768 & _GEN_99023 : ~(_GEN_99361 & _GEN_1768) & _GEN_99023) : _GEN_99023;
  wire        _GEN_99260 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1769 & _GEN_99024 : _GEN_987 ? ~_GEN_1769 & _GEN_99024 : ~(_GEN_99361 & _GEN_1769) & _GEN_99024) : _GEN_99024;
  wire        _GEN_99261 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1770 & _GEN_99025 : _GEN_987 ? ~_GEN_1770 & _GEN_99025 : ~(_GEN_99361 & _GEN_1770) & _GEN_99025) : _GEN_99025;
  wire        _GEN_99262 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1771 & _GEN_99026 : _GEN_987 ? ~_GEN_1771 & _GEN_99026 : ~(_GEN_99361 & _GEN_1771) & _GEN_99026) : _GEN_99026;
  wire        _GEN_99263 = _GEN_985 ? (_GEN_99196 ? ~_GEN_1772 & _GEN_99027 : _GEN_987 ? ~_GEN_1772 & _GEN_99027 : ~(_GEN_99361 & _GEN_1772) & _GEN_99027) : _GEN_99027;
  wire        _GEN_99264 = _GEN_985 ? (_GEN_99196 ? ~(&lcam_ldq_idx_0) & _GEN_98530 : _GEN_987 ? ~(&lcam_ldq_idx_0) & _GEN_98530 : ~(_GEN_99361 & (&lcam_ldq_idx_0)) & _GEN_98530) : _GEN_98530;
  wire        _GEN_99467 = _GEN_988 ? (_GEN_99430 ? (|lcam_ldq_idx_1) & _GEN_99233 : _GEN_990 ? (|lcam_ldq_idx_1) & _GEN_99233 : ~(_GEN_99361 & ~(|lcam_ldq_idx_1)) & _GEN_99233) : _GEN_99233;
  wire        _GEN_99468 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1773 & _GEN_99234 : _GEN_990 ? ~_GEN_1773 & _GEN_99234 : ~(_GEN_99361 & _GEN_1773) & _GEN_99234) : _GEN_99234;
  wire        _GEN_99469 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1774 & _GEN_99235 : _GEN_990 ? ~_GEN_1774 & _GEN_99235 : ~(_GEN_99361 & _GEN_1774) & _GEN_99235) : _GEN_99235;
  wire        _GEN_99470 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1775 & _GEN_99236 : _GEN_990 ? ~_GEN_1775 & _GEN_99236 : ~(_GEN_99361 & _GEN_1775) & _GEN_99236) : _GEN_99236;
  wire        _GEN_99471 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1776 & _GEN_99237 : _GEN_990 ? ~_GEN_1776 & _GEN_99237 : ~(_GEN_99361 & _GEN_1776) & _GEN_99237) : _GEN_99237;
  wire        _GEN_99472 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1777 & _GEN_99238 : _GEN_990 ? ~_GEN_1777 & _GEN_99238 : ~(_GEN_99361 & _GEN_1777) & _GEN_99238) : _GEN_99238;
  wire        _GEN_99473 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1778 & _GEN_99239 : _GEN_990 ? ~_GEN_1778 & _GEN_99239 : ~(_GEN_99361 & _GEN_1778) & _GEN_99239) : _GEN_99239;
  wire        _GEN_99474 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1779 & _GEN_99240 : _GEN_990 ? ~_GEN_1779 & _GEN_99240 : ~(_GEN_99361 & _GEN_1779) & _GEN_99240) : _GEN_99240;
  wire        _GEN_99475 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1780 & _GEN_99241 : _GEN_990 ? ~_GEN_1780 & _GEN_99241 : ~(_GEN_99361 & _GEN_1780) & _GEN_99241) : _GEN_99241;
  wire        _GEN_99476 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1781 & _GEN_99242 : _GEN_990 ? ~_GEN_1781 & _GEN_99242 : ~(_GEN_99361 & _GEN_1781) & _GEN_99242) : _GEN_99242;
  wire        _GEN_99477 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1782 & _GEN_99243 : _GEN_990 ? ~_GEN_1782 & _GEN_99243 : ~(_GEN_99361 & _GEN_1782) & _GEN_99243) : _GEN_99243;
  wire        _GEN_99478 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1783 & _GEN_99244 : _GEN_990 ? ~_GEN_1783 & _GEN_99244 : ~(_GEN_99361 & _GEN_1783) & _GEN_99244) : _GEN_99244;
  wire        _GEN_99479 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1784 & _GEN_99245 : _GEN_990 ? ~_GEN_1784 & _GEN_99245 : ~(_GEN_99361 & _GEN_1784) & _GEN_99245) : _GEN_99245;
  wire        _GEN_99480 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1785 & _GEN_99246 : _GEN_990 ? ~_GEN_1785 & _GEN_99246 : ~(_GEN_99361 & _GEN_1785) & _GEN_99246) : _GEN_99246;
  wire        _GEN_99481 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1786 & _GEN_99247 : _GEN_990 ? ~_GEN_1786 & _GEN_99247 : ~(_GEN_99361 & _GEN_1786) & _GEN_99247) : _GEN_99247;
  wire        _GEN_99482 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1787 & _GEN_99248 : _GEN_990 ? ~_GEN_1787 & _GEN_99248 : ~(_GEN_99361 & _GEN_1787) & _GEN_99248) : _GEN_99248;
  wire        _GEN_99483 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1788 & _GEN_99249 : _GEN_990 ? ~_GEN_1788 & _GEN_99249 : ~(_GEN_99361 & _GEN_1788) & _GEN_99249) : _GEN_99249;
  wire        _GEN_99484 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1789 & _GEN_99250 : _GEN_990 ? ~_GEN_1789 & _GEN_99250 : ~(_GEN_99361 & _GEN_1789) & _GEN_99250) : _GEN_99250;
  wire        _GEN_99485 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1790 & _GEN_99251 : _GEN_990 ? ~_GEN_1790 & _GEN_99251 : ~(_GEN_99361 & _GEN_1790) & _GEN_99251) : _GEN_99251;
  wire        _GEN_99486 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1791 & _GEN_99252 : _GEN_990 ? ~_GEN_1791 & _GEN_99252 : ~(_GEN_99361 & _GEN_1791) & _GEN_99252) : _GEN_99252;
  wire        _GEN_99487 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1792 & _GEN_99253 : _GEN_990 ? ~_GEN_1792 & _GEN_99253 : ~(_GEN_99361 & _GEN_1792) & _GEN_99253) : _GEN_99253;
  wire        _GEN_99488 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1793 & _GEN_99254 : _GEN_990 ? ~_GEN_1793 & _GEN_99254 : ~(_GEN_99361 & _GEN_1793) & _GEN_99254) : _GEN_99254;
  wire        _GEN_99489 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1794 & _GEN_99255 : _GEN_990 ? ~_GEN_1794 & _GEN_99255 : ~(_GEN_99361 & _GEN_1794) & _GEN_99255) : _GEN_99255;
  wire        _GEN_99490 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1795 & _GEN_99256 : _GEN_990 ? ~_GEN_1795 & _GEN_99256 : ~(_GEN_99361 & _GEN_1795) & _GEN_99256) : _GEN_99256;
  wire        _GEN_99491 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1796 & _GEN_99257 : _GEN_990 ? ~_GEN_1796 & _GEN_99257 : ~(_GEN_99361 & _GEN_1796) & _GEN_99257) : _GEN_99257;
  wire        _GEN_99492 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1797 & _GEN_99258 : _GEN_990 ? ~_GEN_1797 & _GEN_99258 : ~(_GEN_99361 & _GEN_1797) & _GEN_99258) : _GEN_99258;
  wire        _GEN_99493 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1798 & _GEN_99259 : _GEN_990 ? ~_GEN_1798 & _GEN_99259 : ~(_GEN_99361 & _GEN_1798) & _GEN_99259) : _GEN_99259;
  wire        _GEN_99494 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1799 & _GEN_99260 : _GEN_990 ? ~_GEN_1799 & _GEN_99260 : ~(_GEN_99361 & _GEN_1799) & _GEN_99260) : _GEN_99260;
  wire        _GEN_99495 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1800 & _GEN_99261 : _GEN_990 ? ~_GEN_1800 & _GEN_99261 : ~(_GEN_99361 & _GEN_1800) & _GEN_99261) : _GEN_99261;
  wire        _GEN_99496 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1801 & _GEN_99262 : _GEN_990 ? ~_GEN_1801 & _GEN_99262 : ~(_GEN_99361 & _GEN_1801) & _GEN_99262) : _GEN_99262;
  wire        _GEN_99497 = _GEN_988 ? (_GEN_99430 ? ~_GEN_1802 & _GEN_99263 : _GEN_990 ? ~_GEN_1802 & _GEN_99263 : ~(_GEN_99361 & _GEN_1802) & _GEN_99263) : _GEN_99263;
  wire        _GEN_99498 = _GEN_988 ? (_GEN_99430 ? ~(&lcam_ldq_idx_1) & _GEN_99264 : _GEN_990 ? ~(&lcam_ldq_idx_1) & _GEN_99264 : ~(_GEN_99361 & (&lcam_ldq_idx_1)) & _GEN_99264) : _GEN_99264;
  wire        _GEN_99701 = _GEN_991 ? (_GEN_99664 ? (|lcam_ldq_idx_0) & _GEN_99467 : _GEN_993 ? (|lcam_ldq_idx_0) & _GEN_99467 : ~(_GEN_99829 & ~(|lcam_ldq_idx_0)) & _GEN_99467) : _GEN_99467;
  wire        _GEN_99702 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1743 & _GEN_99468 : _GEN_993 ? ~_GEN_1743 & _GEN_99468 : ~(_GEN_99829 & _GEN_1743) & _GEN_99468) : _GEN_99468;
  wire        _GEN_99703 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1744 & _GEN_99469 : _GEN_993 ? ~_GEN_1744 & _GEN_99469 : ~(_GEN_99829 & _GEN_1744) & _GEN_99469) : _GEN_99469;
  wire        _GEN_99704 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1745 & _GEN_99470 : _GEN_993 ? ~_GEN_1745 & _GEN_99470 : ~(_GEN_99829 & _GEN_1745) & _GEN_99470) : _GEN_99470;
  wire        _GEN_99705 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1746 & _GEN_99471 : _GEN_993 ? ~_GEN_1746 & _GEN_99471 : ~(_GEN_99829 & _GEN_1746) & _GEN_99471) : _GEN_99471;
  wire        _GEN_99706 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1747 & _GEN_99472 : _GEN_993 ? ~_GEN_1747 & _GEN_99472 : ~(_GEN_99829 & _GEN_1747) & _GEN_99472) : _GEN_99472;
  wire        _GEN_99707 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1748 & _GEN_99473 : _GEN_993 ? ~_GEN_1748 & _GEN_99473 : ~(_GEN_99829 & _GEN_1748) & _GEN_99473) : _GEN_99473;
  wire        _GEN_99708 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1749 & _GEN_99474 : _GEN_993 ? ~_GEN_1749 & _GEN_99474 : ~(_GEN_99829 & _GEN_1749) & _GEN_99474) : _GEN_99474;
  wire        _GEN_99709 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1750 & _GEN_99475 : _GEN_993 ? ~_GEN_1750 & _GEN_99475 : ~(_GEN_99829 & _GEN_1750) & _GEN_99475) : _GEN_99475;
  wire        _GEN_99710 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1751 & _GEN_99476 : _GEN_993 ? ~_GEN_1751 & _GEN_99476 : ~(_GEN_99829 & _GEN_1751) & _GEN_99476) : _GEN_99476;
  wire        _GEN_99711 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1752 & _GEN_99477 : _GEN_993 ? ~_GEN_1752 & _GEN_99477 : ~(_GEN_99829 & _GEN_1752) & _GEN_99477) : _GEN_99477;
  wire        _GEN_99712 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1753 & _GEN_99478 : _GEN_993 ? ~_GEN_1753 & _GEN_99478 : ~(_GEN_99829 & _GEN_1753) & _GEN_99478) : _GEN_99478;
  wire        _GEN_99713 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1754 & _GEN_99479 : _GEN_993 ? ~_GEN_1754 & _GEN_99479 : ~(_GEN_99829 & _GEN_1754) & _GEN_99479) : _GEN_99479;
  wire        _GEN_99714 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1755 & _GEN_99480 : _GEN_993 ? ~_GEN_1755 & _GEN_99480 : ~(_GEN_99829 & _GEN_1755) & _GEN_99480) : _GEN_99480;
  wire        _GEN_99715 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1756 & _GEN_99481 : _GEN_993 ? ~_GEN_1756 & _GEN_99481 : ~(_GEN_99829 & _GEN_1756) & _GEN_99481) : _GEN_99481;
  wire        _GEN_99716 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1757 & _GEN_99482 : _GEN_993 ? ~_GEN_1757 & _GEN_99482 : ~(_GEN_99829 & _GEN_1757) & _GEN_99482) : _GEN_99482;
  wire        _GEN_99717 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1758 & _GEN_99483 : _GEN_993 ? ~_GEN_1758 & _GEN_99483 : ~(_GEN_99829 & _GEN_1758) & _GEN_99483) : _GEN_99483;
  wire        _GEN_99718 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1759 & _GEN_99484 : _GEN_993 ? ~_GEN_1759 & _GEN_99484 : ~(_GEN_99829 & _GEN_1759) & _GEN_99484) : _GEN_99484;
  wire        _GEN_99719 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1760 & _GEN_99485 : _GEN_993 ? ~_GEN_1760 & _GEN_99485 : ~(_GEN_99829 & _GEN_1760) & _GEN_99485) : _GEN_99485;
  wire        _GEN_99720 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1761 & _GEN_99486 : _GEN_993 ? ~_GEN_1761 & _GEN_99486 : ~(_GEN_99829 & _GEN_1761) & _GEN_99486) : _GEN_99486;
  wire        _GEN_99721 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1762 & _GEN_99487 : _GEN_993 ? ~_GEN_1762 & _GEN_99487 : ~(_GEN_99829 & _GEN_1762) & _GEN_99487) : _GEN_99487;
  wire        _GEN_99722 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1763 & _GEN_99488 : _GEN_993 ? ~_GEN_1763 & _GEN_99488 : ~(_GEN_99829 & _GEN_1763) & _GEN_99488) : _GEN_99488;
  wire        _GEN_99723 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1764 & _GEN_99489 : _GEN_993 ? ~_GEN_1764 & _GEN_99489 : ~(_GEN_99829 & _GEN_1764) & _GEN_99489) : _GEN_99489;
  wire        _GEN_99724 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1765 & _GEN_99490 : _GEN_993 ? ~_GEN_1765 & _GEN_99490 : ~(_GEN_99829 & _GEN_1765) & _GEN_99490) : _GEN_99490;
  wire        _GEN_99725 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1766 & _GEN_99491 : _GEN_993 ? ~_GEN_1766 & _GEN_99491 : ~(_GEN_99829 & _GEN_1766) & _GEN_99491) : _GEN_99491;
  wire        _GEN_99726 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1767 & _GEN_99492 : _GEN_993 ? ~_GEN_1767 & _GEN_99492 : ~(_GEN_99829 & _GEN_1767) & _GEN_99492) : _GEN_99492;
  wire        _GEN_99727 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1768 & _GEN_99493 : _GEN_993 ? ~_GEN_1768 & _GEN_99493 : ~(_GEN_99829 & _GEN_1768) & _GEN_99493) : _GEN_99493;
  wire        _GEN_99728 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1769 & _GEN_99494 : _GEN_993 ? ~_GEN_1769 & _GEN_99494 : ~(_GEN_99829 & _GEN_1769) & _GEN_99494) : _GEN_99494;
  wire        _GEN_99729 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1770 & _GEN_99495 : _GEN_993 ? ~_GEN_1770 & _GEN_99495 : ~(_GEN_99829 & _GEN_1770) & _GEN_99495) : _GEN_99495;
  wire        _GEN_99730 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1771 & _GEN_99496 : _GEN_993 ? ~_GEN_1771 & _GEN_99496 : ~(_GEN_99829 & _GEN_1771) & _GEN_99496) : _GEN_99496;
  wire        _GEN_99731 = _GEN_991 ? (_GEN_99664 ? ~_GEN_1772 & _GEN_99497 : _GEN_993 ? ~_GEN_1772 & _GEN_99497 : ~(_GEN_99829 & _GEN_1772) & _GEN_99497) : _GEN_99497;
  wire        _GEN_99732 = _GEN_991 ? (_GEN_99664 ? ~(&lcam_ldq_idx_0) & _GEN_99498 : _GEN_993 ? ~(&lcam_ldq_idx_0) & _GEN_99498 : ~(_GEN_99829 & (&lcam_ldq_idx_0)) & _GEN_99498) : _GEN_99498;
  wire        _GEN_99935 = _GEN_994 ? (_GEN_99898 ? (|lcam_ldq_idx_1) & _GEN_99701 : _GEN_996 ? (|lcam_ldq_idx_1) & _GEN_99701 : ~(_GEN_99829 & ~(|lcam_ldq_idx_1)) & _GEN_99701) : _GEN_99701;
  wire        _GEN_99936 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1773 & _GEN_99702 : _GEN_996 ? ~_GEN_1773 & _GEN_99702 : ~(_GEN_99829 & _GEN_1773) & _GEN_99702) : _GEN_99702;
  wire        _GEN_99937 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1774 & _GEN_99703 : _GEN_996 ? ~_GEN_1774 & _GEN_99703 : ~(_GEN_99829 & _GEN_1774) & _GEN_99703) : _GEN_99703;
  wire        _GEN_99938 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1775 & _GEN_99704 : _GEN_996 ? ~_GEN_1775 & _GEN_99704 : ~(_GEN_99829 & _GEN_1775) & _GEN_99704) : _GEN_99704;
  wire        _GEN_99939 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1776 & _GEN_99705 : _GEN_996 ? ~_GEN_1776 & _GEN_99705 : ~(_GEN_99829 & _GEN_1776) & _GEN_99705) : _GEN_99705;
  wire        _GEN_99940 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1777 & _GEN_99706 : _GEN_996 ? ~_GEN_1777 & _GEN_99706 : ~(_GEN_99829 & _GEN_1777) & _GEN_99706) : _GEN_99706;
  wire        _GEN_99941 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1778 & _GEN_99707 : _GEN_996 ? ~_GEN_1778 & _GEN_99707 : ~(_GEN_99829 & _GEN_1778) & _GEN_99707) : _GEN_99707;
  wire        _GEN_99942 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1779 & _GEN_99708 : _GEN_996 ? ~_GEN_1779 & _GEN_99708 : ~(_GEN_99829 & _GEN_1779) & _GEN_99708) : _GEN_99708;
  wire        _GEN_99943 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1780 & _GEN_99709 : _GEN_996 ? ~_GEN_1780 & _GEN_99709 : ~(_GEN_99829 & _GEN_1780) & _GEN_99709) : _GEN_99709;
  wire        _GEN_99944 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1781 & _GEN_99710 : _GEN_996 ? ~_GEN_1781 & _GEN_99710 : ~(_GEN_99829 & _GEN_1781) & _GEN_99710) : _GEN_99710;
  wire        _GEN_99945 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1782 & _GEN_99711 : _GEN_996 ? ~_GEN_1782 & _GEN_99711 : ~(_GEN_99829 & _GEN_1782) & _GEN_99711) : _GEN_99711;
  wire        _GEN_99946 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1783 & _GEN_99712 : _GEN_996 ? ~_GEN_1783 & _GEN_99712 : ~(_GEN_99829 & _GEN_1783) & _GEN_99712) : _GEN_99712;
  wire        _GEN_99947 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1784 & _GEN_99713 : _GEN_996 ? ~_GEN_1784 & _GEN_99713 : ~(_GEN_99829 & _GEN_1784) & _GEN_99713) : _GEN_99713;
  wire        _GEN_99948 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1785 & _GEN_99714 : _GEN_996 ? ~_GEN_1785 & _GEN_99714 : ~(_GEN_99829 & _GEN_1785) & _GEN_99714) : _GEN_99714;
  wire        _GEN_99949 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1786 & _GEN_99715 : _GEN_996 ? ~_GEN_1786 & _GEN_99715 : ~(_GEN_99829 & _GEN_1786) & _GEN_99715) : _GEN_99715;
  wire        _GEN_99950 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1787 & _GEN_99716 : _GEN_996 ? ~_GEN_1787 & _GEN_99716 : ~(_GEN_99829 & _GEN_1787) & _GEN_99716) : _GEN_99716;
  wire        _GEN_99951 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1788 & _GEN_99717 : _GEN_996 ? ~_GEN_1788 & _GEN_99717 : ~(_GEN_99829 & _GEN_1788) & _GEN_99717) : _GEN_99717;
  wire        _GEN_99952 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1789 & _GEN_99718 : _GEN_996 ? ~_GEN_1789 & _GEN_99718 : ~(_GEN_99829 & _GEN_1789) & _GEN_99718) : _GEN_99718;
  wire        _GEN_99953 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1790 & _GEN_99719 : _GEN_996 ? ~_GEN_1790 & _GEN_99719 : ~(_GEN_99829 & _GEN_1790) & _GEN_99719) : _GEN_99719;
  wire        _GEN_99954 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1791 & _GEN_99720 : _GEN_996 ? ~_GEN_1791 & _GEN_99720 : ~(_GEN_99829 & _GEN_1791) & _GEN_99720) : _GEN_99720;
  wire        _GEN_99955 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1792 & _GEN_99721 : _GEN_996 ? ~_GEN_1792 & _GEN_99721 : ~(_GEN_99829 & _GEN_1792) & _GEN_99721) : _GEN_99721;
  wire        _GEN_99956 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1793 & _GEN_99722 : _GEN_996 ? ~_GEN_1793 & _GEN_99722 : ~(_GEN_99829 & _GEN_1793) & _GEN_99722) : _GEN_99722;
  wire        _GEN_99957 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1794 & _GEN_99723 : _GEN_996 ? ~_GEN_1794 & _GEN_99723 : ~(_GEN_99829 & _GEN_1794) & _GEN_99723) : _GEN_99723;
  wire        _GEN_99958 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1795 & _GEN_99724 : _GEN_996 ? ~_GEN_1795 & _GEN_99724 : ~(_GEN_99829 & _GEN_1795) & _GEN_99724) : _GEN_99724;
  wire        _GEN_99959 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1796 & _GEN_99725 : _GEN_996 ? ~_GEN_1796 & _GEN_99725 : ~(_GEN_99829 & _GEN_1796) & _GEN_99725) : _GEN_99725;
  wire        _GEN_99960 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1797 & _GEN_99726 : _GEN_996 ? ~_GEN_1797 & _GEN_99726 : ~(_GEN_99829 & _GEN_1797) & _GEN_99726) : _GEN_99726;
  wire        _GEN_99961 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1798 & _GEN_99727 : _GEN_996 ? ~_GEN_1798 & _GEN_99727 : ~(_GEN_99829 & _GEN_1798) & _GEN_99727) : _GEN_99727;
  wire        _GEN_99962 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1799 & _GEN_99728 : _GEN_996 ? ~_GEN_1799 & _GEN_99728 : ~(_GEN_99829 & _GEN_1799) & _GEN_99728) : _GEN_99728;
  wire        _GEN_99963 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1800 & _GEN_99729 : _GEN_996 ? ~_GEN_1800 & _GEN_99729 : ~(_GEN_99829 & _GEN_1800) & _GEN_99729) : _GEN_99729;
  wire        _GEN_99964 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1801 & _GEN_99730 : _GEN_996 ? ~_GEN_1801 & _GEN_99730 : ~(_GEN_99829 & _GEN_1801) & _GEN_99730) : _GEN_99730;
  wire        _GEN_99965 = _GEN_994 ? (_GEN_99898 ? ~_GEN_1802 & _GEN_99731 : _GEN_996 ? ~_GEN_1802 & _GEN_99731 : ~(_GEN_99829 & _GEN_1802) & _GEN_99731) : _GEN_99731;
  wire        _GEN_99966 = _GEN_994 ? (_GEN_99898 ? ~(&lcam_ldq_idx_1) & _GEN_99732 : _GEN_996 ? ~(&lcam_ldq_idx_1) & _GEN_99732 : ~(_GEN_99829 & (&lcam_ldq_idx_1)) & _GEN_99732) : _GEN_99732;
  wire        _GEN_100169 = _GEN_997 ? (_GEN_100132 ? (|lcam_ldq_idx_0) & _GEN_99935 : _GEN_999 ? (|lcam_ldq_idx_0) & _GEN_99935 : ~(_GEN_100297 & ~(|lcam_ldq_idx_0)) & _GEN_99935) : _GEN_99935;
  wire        _GEN_100170 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1743 & _GEN_99936 : _GEN_999 ? ~_GEN_1743 & _GEN_99936 : ~(_GEN_100297 & _GEN_1743) & _GEN_99936) : _GEN_99936;
  wire        _GEN_100171 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1744 & _GEN_99937 : _GEN_999 ? ~_GEN_1744 & _GEN_99937 : ~(_GEN_100297 & _GEN_1744) & _GEN_99937) : _GEN_99937;
  wire        _GEN_100172 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1745 & _GEN_99938 : _GEN_999 ? ~_GEN_1745 & _GEN_99938 : ~(_GEN_100297 & _GEN_1745) & _GEN_99938) : _GEN_99938;
  wire        _GEN_100173 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1746 & _GEN_99939 : _GEN_999 ? ~_GEN_1746 & _GEN_99939 : ~(_GEN_100297 & _GEN_1746) & _GEN_99939) : _GEN_99939;
  wire        _GEN_100174 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1747 & _GEN_99940 : _GEN_999 ? ~_GEN_1747 & _GEN_99940 : ~(_GEN_100297 & _GEN_1747) & _GEN_99940) : _GEN_99940;
  wire        _GEN_100175 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1748 & _GEN_99941 : _GEN_999 ? ~_GEN_1748 & _GEN_99941 : ~(_GEN_100297 & _GEN_1748) & _GEN_99941) : _GEN_99941;
  wire        _GEN_100176 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1749 & _GEN_99942 : _GEN_999 ? ~_GEN_1749 & _GEN_99942 : ~(_GEN_100297 & _GEN_1749) & _GEN_99942) : _GEN_99942;
  wire        _GEN_100177 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1750 & _GEN_99943 : _GEN_999 ? ~_GEN_1750 & _GEN_99943 : ~(_GEN_100297 & _GEN_1750) & _GEN_99943) : _GEN_99943;
  wire        _GEN_100178 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1751 & _GEN_99944 : _GEN_999 ? ~_GEN_1751 & _GEN_99944 : ~(_GEN_100297 & _GEN_1751) & _GEN_99944) : _GEN_99944;
  wire        _GEN_100179 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1752 & _GEN_99945 : _GEN_999 ? ~_GEN_1752 & _GEN_99945 : ~(_GEN_100297 & _GEN_1752) & _GEN_99945) : _GEN_99945;
  wire        _GEN_100180 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1753 & _GEN_99946 : _GEN_999 ? ~_GEN_1753 & _GEN_99946 : ~(_GEN_100297 & _GEN_1753) & _GEN_99946) : _GEN_99946;
  wire        _GEN_100181 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1754 & _GEN_99947 : _GEN_999 ? ~_GEN_1754 & _GEN_99947 : ~(_GEN_100297 & _GEN_1754) & _GEN_99947) : _GEN_99947;
  wire        _GEN_100182 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1755 & _GEN_99948 : _GEN_999 ? ~_GEN_1755 & _GEN_99948 : ~(_GEN_100297 & _GEN_1755) & _GEN_99948) : _GEN_99948;
  wire        _GEN_100183 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1756 & _GEN_99949 : _GEN_999 ? ~_GEN_1756 & _GEN_99949 : ~(_GEN_100297 & _GEN_1756) & _GEN_99949) : _GEN_99949;
  wire        _GEN_100184 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1757 & _GEN_99950 : _GEN_999 ? ~_GEN_1757 & _GEN_99950 : ~(_GEN_100297 & _GEN_1757) & _GEN_99950) : _GEN_99950;
  wire        _GEN_100185 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1758 & _GEN_99951 : _GEN_999 ? ~_GEN_1758 & _GEN_99951 : ~(_GEN_100297 & _GEN_1758) & _GEN_99951) : _GEN_99951;
  wire        _GEN_100186 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1759 & _GEN_99952 : _GEN_999 ? ~_GEN_1759 & _GEN_99952 : ~(_GEN_100297 & _GEN_1759) & _GEN_99952) : _GEN_99952;
  wire        _GEN_100187 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1760 & _GEN_99953 : _GEN_999 ? ~_GEN_1760 & _GEN_99953 : ~(_GEN_100297 & _GEN_1760) & _GEN_99953) : _GEN_99953;
  wire        _GEN_100188 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1761 & _GEN_99954 : _GEN_999 ? ~_GEN_1761 & _GEN_99954 : ~(_GEN_100297 & _GEN_1761) & _GEN_99954) : _GEN_99954;
  wire        _GEN_100189 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1762 & _GEN_99955 : _GEN_999 ? ~_GEN_1762 & _GEN_99955 : ~(_GEN_100297 & _GEN_1762) & _GEN_99955) : _GEN_99955;
  wire        _GEN_100190 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1763 & _GEN_99956 : _GEN_999 ? ~_GEN_1763 & _GEN_99956 : ~(_GEN_100297 & _GEN_1763) & _GEN_99956) : _GEN_99956;
  wire        _GEN_100191 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1764 & _GEN_99957 : _GEN_999 ? ~_GEN_1764 & _GEN_99957 : ~(_GEN_100297 & _GEN_1764) & _GEN_99957) : _GEN_99957;
  wire        _GEN_100192 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1765 & _GEN_99958 : _GEN_999 ? ~_GEN_1765 & _GEN_99958 : ~(_GEN_100297 & _GEN_1765) & _GEN_99958) : _GEN_99958;
  wire        _GEN_100193 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1766 & _GEN_99959 : _GEN_999 ? ~_GEN_1766 & _GEN_99959 : ~(_GEN_100297 & _GEN_1766) & _GEN_99959) : _GEN_99959;
  wire        _GEN_100194 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1767 & _GEN_99960 : _GEN_999 ? ~_GEN_1767 & _GEN_99960 : ~(_GEN_100297 & _GEN_1767) & _GEN_99960) : _GEN_99960;
  wire        _GEN_100195 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1768 & _GEN_99961 : _GEN_999 ? ~_GEN_1768 & _GEN_99961 : ~(_GEN_100297 & _GEN_1768) & _GEN_99961) : _GEN_99961;
  wire        _GEN_100196 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1769 & _GEN_99962 : _GEN_999 ? ~_GEN_1769 & _GEN_99962 : ~(_GEN_100297 & _GEN_1769) & _GEN_99962) : _GEN_99962;
  wire        _GEN_100197 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1770 & _GEN_99963 : _GEN_999 ? ~_GEN_1770 & _GEN_99963 : ~(_GEN_100297 & _GEN_1770) & _GEN_99963) : _GEN_99963;
  wire        _GEN_100198 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1771 & _GEN_99964 : _GEN_999 ? ~_GEN_1771 & _GEN_99964 : ~(_GEN_100297 & _GEN_1771) & _GEN_99964) : _GEN_99964;
  wire        _GEN_100199 = _GEN_997 ? (_GEN_100132 ? ~_GEN_1772 & _GEN_99965 : _GEN_999 ? ~_GEN_1772 & _GEN_99965 : ~(_GEN_100297 & _GEN_1772) & _GEN_99965) : _GEN_99965;
  wire        _GEN_100200 = _GEN_997 ? (_GEN_100132 ? ~(&lcam_ldq_idx_0) & _GEN_99966 : _GEN_999 ? ~(&lcam_ldq_idx_0) & _GEN_99966 : ~(_GEN_100297 & (&lcam_ldq_idx_0)) & _GEN_99966) : _GEN_99966;
  wire        _GEN_100403 = _GEN_1000 ? (_GEN_100366 ? (|lcam_ldq_idx_1) & _GEN_100169 : _GEN_1002 ? (|lcam_ldq_idx_1) & _GEN_100169 : ~(_GEN_100297 & ~(|lcam_ldq_idx_1)) & _GEN_100169) : _GEN_100169;
  wire        _GEN_100404 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1773 & _GEN_100170 : _GEN_1002 ? ~_GEN_1773 & _GEN_100170 : ~(_GEN_100297 & _GEN_1773) & _GEN_100170) : _GEN_100170;
  wire        _GEN_100405 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1774 & _GEN_100171 : _GEN_1002 ? ~_GEN_1774 & _GEN_100171 : ~(_GEN_100297 & _GEN_1774) & _GEN_100171) : _GEN_100171;
  wire        _GEN_100406 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1775 & _GEN_100172 : _GEN_1002 ? ~_GEN_1775 & _GEN_100172 : ~(_GEN_100297 & _GEN_1775) & _GEN_100172) : _GEN_100172;
  wire        _GEN_100407 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1776 & _GEN_100173 : _GEN_1002 ? ~_GEN_1776 & _GEN_100173 : ~(_GEN_100297 & _GEN_1776) & _GEN_100173) : _GEN_100173;
  wire        _GEN_100408 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1777 & _GEN_100174 : _GEN_1002 ? ~_GEN_1777 & _GEN_100174 : ~(_GEN_100297 & _GEN_1777) & _GEN_100174) : _GEN_100174;
  wire        _GEN_100409 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1778 & _GEN_100175 : _GEN_1002 ? ~_GEN_1778 & _GEN_100175 : ~(_GEN_100297 & _GEN_1778) & _GEN_100175) : _GEN_100175;
  wire        _GEN_100410 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1779 & _GEN_100176 : _GEN_1002 ? ~_GEN_1779 & _GEN_100176 : ~(_GEN_100297 & _GEN_1779) & _GEN_100176) : _GEN_100176;
  wire        _GEN_100411 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1780 & _GEN_100177 : _GEN_1002 ? ~_GEN_1780 & _GEN_100177 : ~(_GEN_100297 & _GEN_1780) & _GEN_100177) : _GEN_100177;
  wire        _GEN_100412 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1781 & _GEN_100178 : _GEN_1002 ? ~_GEN_1781 & _GEN_100178 : ~(_GEN_100297 & _GEN_1781) & _GEN_100178) : _GEN_100178;
  wire        _GEN_100413 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1782 & _GEN_100179 : _GEN_1002 ? ~_GEN_1782 & _GEN_100179 : ~(_GEN_100297 & _GEN_1782) & _GEN_100179) : _GEN_100179;
  wire        _GEN_100414 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1783 & _GEN_100180 : _GEN_1002 ? ~_GEN_1783 & _GEN_100180 : ~(_GEN_100297 & _GEN_1783) & _GEN_100180) : _GEN_100180;
  wire        _GEN_100415 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1784 & _GEN_100181 : _GEN_1002 ? ~_GEN_1784 & _GEN_100181 : ~(_GEN_100297 & _GEN_1784) & _GEN_100181) : _GEN_100181;
  wire        _GEN_100416 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1785 & _GEN_100182 : _GEN_1002 ? ~_GEN_1785 & _GEN_100182 : ~(_GEN_100297 & _GEN_1785) & _GEN_100182) : _GEN_100182;
  wire        _GEN_100417 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1786 & _GEN_100183 : _GEN_1002 ? ~_GEN_1786 & _GEN_100183 : ~(_GEN_100297 & _GEN_1786) & _GEN_100183) : _GEN_100183;
  wire        _GEN_100418 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1787 & _GEN_100184 : _GEN_1002 ? ~_GEN_1787 & _GEN_100184 : ~(_GEN_100297 & _GEN_1787) & _GEN_100184) : _GEN_100184;
  wire        _GEN_100419 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1788 & _GEN_100185 : _GEN_1002 ? ~_GEN_1788 & _GEN_100185 : ~(_GEN_100297 & _GEN_1788) & _GEN_100185) : _GEN_100185;
  wire        _GEN_100420 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1789 & _GEN_100186 : _GEN_1002 ? ~_GEN_1789 & _GEN_100186 : ~(_GEN_100297 & _GEN_1789) & _GEN_100186) : _GEN_100186;
  wire        _GEN_100421 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1790 & _GEN_100187 : _GEN_1002 ? ~_GEN_1790 & _GEN_100187 : ~(_GEN_100297 & _GEN_1790) & _GEN_100187) : _GEN_100187;
  wire        _GEN_100422 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1791 & _GEN_100188 : _GEN_1002 ? ~_GEN_1791 & _GEN_100188 : ~(_GEN_100297 & _GEN_1791) & _GEN_100188) : _GEN_100188;
  wire        _GEN_100423 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1792 & _GEN_100189 : _GEN_1002 ? ~_GEN_1792 & _GEN_100189 : ~(_GEN_100297 & _GEN_1792) & _GEN_100189) : _GEN_100189;
  wire        _GEN_100424 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1793 & _GEN_100190 : _GEN_1002 ? ~_GEN_1793 & _GEN_100190 : ~(_GEN_100297 & _GEN_1793) & _GEN_100190) : _GEN_100190;
  wire        _GEN_100425 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1794 & _GEN_100191 : _GEN_1002 ? ~_GEN_1794 & _GEN_100191 : ~(_GEN_100297 & _GEN_1794) & _GEN_100191) : _GEN_100191;
  wire        _GEN_100426 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1795 & _GEN_100192 : _GEN_1002 ? ~_GEN_1795 & _GEN_100192 : ~(_GEN_100297 & _GEN_1795) & _GEN_100192) : _GEN_100192;
  wire        _GEN_100427 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1796 & _GEN_100193 : _GEN_1002 ? ~_GEN_1796 & _GEN_100193 : ~(_GEN_100297 & _GEN_1796) & _GEN_100193) : _GEN_100193;
  wire        _GEN_100428 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1797 & _GEN_100194 : _GEN_1002 ? ~_GEN_1797 & _GEN_100194 : ~(_GEN_100297 & _GEN_1797) & _GEN_100194) : _GEN_100194;
  wire        _GEN_100429 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1798 & _GEN_100195 : _GEN_1002 ? ~_GEN_1798 & _GEN_100195 : ~(_GEN_100297 & _GEN_1798) & _GEN_100195) : _GEN_100195;
  wire        _GEN_100430 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1799 & _GEN_100196 : _GEN_1002 ? ~_GEN_1799 & _GEN_100196 : ~(_GEN_100297 & _GEN_1799) & _GEN_100196) : _GEN_100196;
  wire        _GEN_100431 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1800 & _GEN_100197 : _GEN_1002 ? ~_GEN_1800 & _GEN_100197 : ~(_GEN_100297 & _GEN_1800) & _GEN_100197) : _GEN_100197;
  wire        _GEN_100432 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1801 & _GEN_100198 : _GEN_1002 ? ~_GEN_1801 & _GEN_100198 : ~(_GEN_100297 & _GEN_1801) & _GEN_100198) : _GEN_100198;
  wire        _GEN_100433 = _GEN_1000 ? (_GEN_100366 ? ~_GEN_1802 & _GEN_100199 : _GEN_1002 ? ~_GEN_1802 & _GEN_100199 : ~(_GEN_100297 & _GEN_1802) & _GEN_100199) : _GEN_100199;
  wire        _GEN_100434 = _GEN_1000 ? (_GEN_100366 ? ~(&lcam_ldq_idx_1) & _GEN_100200 : _GEN_1002 ? ~(&lcam_ldq_idx_1) & _GEN_100200 : ~(_GEN_100297 & (&lcam_ldq_idx_1)) & _GEN_100200) : _GEN_100200;
  wire        _GEN_100637 = _GEN_1003 ? (_GEN_100600 ? (|lcam_ldq_idx_0) & _GEN_100403 : _GEN_1005 ? (|lcam_ldq_idx_0) & _GEN_100403 : ~(_GEN_100765 & ~(|lcam_ldq_idx_0)) & _GEN_100403) : _GEN_100403;
  wire        _GEN_100638 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1743 & _GEN_100404 : _GEN_1005 ? ~_GEN_1743 & _GEN_100404 : ~(_GEN_100765 & _GEN_1743) & _GEN_100404) : _GEN_100404;
  wire        _GEN_100639 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1744 & _GEN_100405 : _GEN_1005 ? ~_GEN_1744 & _GEN_100405 : ~(_GEN_100765 & _GEN_1744) & _GEN_100405) : _GEN_100405;
  wire        _GEN_100640 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1745 & _GEN_100406 : _GEN_1005 ? ~_GEN_1745 & _GEN_100406 : ~(_GEN_100765 & _GEN_1745) & _GEN_100406) : _GEN_100406;
  wire        _GEN_100641 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1746 & _GEN_100407 : _GEN_1005 ? ~_GEN_1746 & _GEN_100407 : ~(_GEN_100765 & _GEN_1746) & _GEN_100407) : _GEN_100407;
  wire        _GEN_100642 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1747 & _GEN_100408 : _GEN_1005 ? ~_GEN_1747 & _GEN_100408 : ~(_GEN_100765 & _GEN_1747) & _GEN_100408) : _GEN_100408;
  wire        _GEN_100643 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1748 & _GEN_100409 : _GEN_1005 ? ~_GEN_1748 & _GEN_100409 : ~(_GEN_100765 & _GEN_1748) & _GEN_100409) : _GEN_100409;
  wire        _GEN_100644 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1749 & _GEN_100410 : _GEN_1005 ? ~_GEN_1749 & _GEN_100410 : ~(_GEN_100765 & _GEN_1749) & _GEN_100410) : _GEN_100410;
  wire        _GEN_100645 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1750 & _GEN_100411 : _GEN_1005 ? ~_GEN_1750 & _GEN_100411 : ~(_GEN_100765 & _GEN_1750) & _GEN_100411) : _GEN_100411;
  wire        _GEN_100646 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1751 & _GEN_100412 : _GEN_1005 ? ~_GEN_1751 & _GEN_100412 : ~(_GEN_100765 & _GEN_1751) & _GEN_100412) : _GEN_100412;
  wire        _GEN_100647 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1752 & _GEN_100413 : _GEN_1005 ? ~_GEN_1752 & _GEN_100413 : ~(_GEN_100765 & _GEN_1752) & _GEN_100413) : _GEN_100413;
  wire        _GEN_100648 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1753 & _GEN_100414 : _GEN_1005 ? ~_GEN_1753 & _GEN_100414 : ~(_GEN_100765 & _GEN_1753) & _GEN_100414) : _GEN_100414;
  wire        _GEN_100649 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1754 & _GEN_100415 : _GEN_1005 ? ~_GEN_1754 & _GEN_100415 : ~(_GEN_100765 & _GEN_1754) & _GEN_100415) : _GEN_100415;
  wire        _GEN_100650 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1755 & _GEN_100416 : _GEN_1005 ? ~_GEN_1755 & _GEN_100416 : ~(_GEN_100765 & _GEN_1755) & _GEN_100416) : _GEN_100416;
  wire        _GEN_100651 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1756 & _GEN_100417 : _GEN_1005 ? ~_GEN_1756 & _GEN_100417 : ~(_GEN_100765 & _GEN_1756) & _GEN_100417) : _GEN_100417;
  wire        _GEN_100652 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1757 & _GEN_100418 : _GEN_1005 ? ~_GEN_1757 & _GEN_100418 : ~(_GEN_100765 & _GEN_1757) & _GEN_100418) : _GEN_100418;
  wire        _GEN_100653 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1758 & _GEN_100419 : _GEN_1005 ? ~_GEN_1758 & _GEN_100419 : ~(_GEN_100765 & _GEN_1758) & _GEN_100419) : _GEN_100419;
  wire        _GEN_100654 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1759 & _GEN_100420 : _GEN_1005 ? ~_GEN_1759 & _GEN_100420 : ~(_GEN_100765 & _GEN_1759) & _GEN_100420) : _GEN_100420;
  wire        _GEN_100655 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1760 & _GEN_100421 : _GEN_1005 ? ~_GEN_1760 & _GEN_100421 : ~(_GEN_100765 & _GEN_1760) & _GEN_100421) : _GEN_100421;
  wire        _GEN_100656 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1761 & _GEN_100422 : _GEN_1005 ? ~_GEN_1761 & _GEN_100422 : ~(_GEN_100765 & _GEN_1761) & _GEN_100422) : _GEN_100422;
  wire        _GEN_100657 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1762 & _GEN_100423 : _GEN_1005 ? ~_GEN_1762 & _GEN_100423 : ~(_GEN_100765 & _GEN_1762) & _GEN_100423) : _GEN_100423;
  wire        _GEN_100658 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1763 & _GEN_100424 : _GEN_1005 ? ~_GEN_1763 & _GEN_100424 : ~(_GEN_100765 & _GEN_1763) & _GEN_100424) : _GEN_100424;
  wire        _GEN_100659 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1764 & _GEN_100425 : _GEN_1005 ? ~_GEN_1764 & _GEN_100425 : ~(_GEN_100765 & _GEN_1764) & _GEN_100425) : _GEN_100425;
  wire        _GEN_100660 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1765 & _GEN_100426 : _GEN_1005 ? ~_GEN_1765 & _GEN_100426 : ~(_GEN_100765 & _GEN_1765) & _GEN_100426) : _GEN_100426;
  wire        _GEN_100661 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1766 & _GEN_100427 : _GEN_1005 ? ~_GEN_1766 & _GEN_100427 : ~(_GEN_100765 & _GEN_1766) & _GEN_100427) : _GEN_100427;
  wire        _GEN_100662 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1767 & _GEN_100428 : _GEN_1005 ? ~_GEN_1767 & _GEN_100428 : ~(_GEN_100765 & _GEN_1767) & _GEN_100428) : _GEN_100428;
  wire        _GEN_100663 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1768 & _GEN_100429 : _GEN_1005 ? ~_GEN_1768 & _GEN_100429 : ~(_GEN_100765 & _GEN_1768) & _GEN_100429) : _GEN_100429;
  wire        _GEN_100664 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1769 & _GEN_100430 : _GEN_1005 ? ~_GEN_1769 & _GEN_100430 : ~(_GEN_100765 & _GEN_1769) & _GEN_100430) : _GEN_100430;
  wire        _GEN_100665 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1770 & _GEN_100431 : _GEN_1005 ? ~_GEN_1770 & _GEN_100431 : ~(_GEN_100765 & _GEN_1770) & _GEN_100431) : _GEN_100431;
  wire        _GEN_100666 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1771 & _GEN_100432 : _GEN_1005 ? ~_GEN_1771 & _GEN_100432 : ~(_GEN_100765 & _GEN_1771) & _GEN_100432) : _GEN_100432;
  wire        _GEN_100667 = _GEN_1003 ? (_GEN_100600 ? ~_GEN_1772 & _GEN_100433 : _GEN_1005 ? ~_GEN_1772 & _GEN_100433 : ~(_GEN_100765 & _GEN_1772) & _GEN_100433) : _GEN_100433;
  wire        _GEN_100668 = _GEN_1003 ? (_GEN_100600 ? ~(&lcam_ldq_idx_0) & _GEN_100434 : _GEN_1005 ? ~(&lcam_ldq_idx_0) & _GEN_100434 : ~(_GEN_100765 & (&lcam_ldq_idx_0)) & _GEN_100434) : _GEN_100434;
  wire        _GEN_100871 = _GEN_1006 ? (_GEN_100834 ? (|lcam_ldq_idx_1) & _GEN_100637 : _GEN_1008 ? (|lcam_ldq_idx_1) & _GEN_100637 : ~(_GEN_100765 & ~(|lcam_ldq_idx_1)) & _GEN_100637) : _GEN_100637;
  wire        _GEN_100872 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1773 & _GEN_100638 : _GEN_1008 ? ~_GEN_1773 & _GEN_100638 : ~(_GEN_100765 & _GEN_1773) & _GEN_100638) : _GEN_100638;
  wire        _GEN_100873 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1774 & _GEN_100639 : _GEN_1008 ? ~_GEN_1774 & _GEN_100639 : ~(_GEN_100765 & _GEN_1774) & _GEN_100639) : _GEN_100639;
  wire        _GEN_100874 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1775 & _GEN_100640 : _GEN_1008 ? ~_GEN_1775 & _GEN_100640 : ~(_GEN_100765 & _GEN_1775) & _GEN_100640) : _GEN_100640;
  wire        _GEN_100875 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1776 & _GEN_100641 : _GEN_1008 ? ~_GEN_1776 & _GEN_100641 : ~(_GEN_100765 & _GEN_1776) & _GEN_100641) : _GEN_100641;
  wire        _GEN_100876 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1777 & _GEN_100642 : _GEN_1008 ? ~_GEN_1777 & _GEN_100642 : ~(_GEN_100765 & _GEN_1777) & _GEN_100642) : _GEN_100642;
  wire        _GEN_100877 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1778 & _GEN_100643 : _GEN_1008 ? ~_GEN_1778 & _GEN_100643 : ~(_GEN_100765 & _GEN_1778) & _GEN_100643) : _GEN_100643;
  wire        _GEN_100878 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1779 & _GEN_100644 : _GEN_1008 ? ~_GEN_1779 & _GEN_100644 : ~(_GEN_100765 & _GEN_1779) & _GEN_100644) : _GEN_100644;
  wire        _GEN_100879 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1780 & _GEN_100645 : _GEN_1008 ? ~_GEN_1780 & _GEN_100645 : ~(_GEN_100765 & _GEN_1780) & _GEN_100645) : _GEN_100645;
  wire        _GEN_100880 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1781 & _GEN_100646 : _GEN_1008 ? ~_GEN_1781 & _GEN_100646 : ~(_GEN_100765 & _GEN_1781) & _GEN_100646) : _GEN_100646;
  wire        _GEN_100881 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1782 & _GEN_100647 : _GEN_1008 ? ~_GEN_1782 & _GEN_100647 : ~(_GEN_100765 & _GEN_1782) & _GEN_100647) : _GEN_100647;
  wire        _GEN_100882 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1783 & _GEN_100648 : _GEN_1008 ? ~_GEN_1783 & _GEN_100648 : ~(_GEN_100765 & _GEN_1783) & _GEN_100648) : _GEN_100648;
  wire        _GEN_100883 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1784 & _GEN_100649 : _GEN_1008 ? ~_GEN_1784 & _GEN_100649 : ~(_GEN_100765 & _GEN_1784) & _GEN_100649) : _GEN_100649;
  wire        _GEN_100884 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1785 & _GEN_100650 : _GEN_1008 ? ~_GEN_1785 & _GEN_100650 : ~(_GEN_100765 & _GEN_1785) & _GEN_100650) : _GEN_100650;
  wire        _GEN_100885 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1786 & _GEN_100651 : _GEN_1008 ? ~_GEN_1786 & _GEN_100651 : ~(_GEN_100765 & _GEN_1786) & _GEN_100651) : _GEN_100651;
  wire        _GEN_100886 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1787 & _GEN_100652 : _GEN_1008 ? ~_GEN_1787 & _GEN_100652 : ~(_GEN_100765 & _GEN_1787) & _GEN_100652) : _GEN_100652;
  wire        _GEN_100887 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1788 & _GEN_100653 : _GEN_1008 ? ~_GEN_1788 & _GEN_100653 : ~(_GEN_100765 & _GEN_1788) & _GEN_100653) : _GEN_100653;
  wire        _GEN_100888 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1789 & _GEN_100654 : _GEN_1008 ? ~_GEN_1789 & _GEN_100654 : ~(_GEN_100765 & _GEN_1789) & _GEN_100654) : _GEN_100654;
  wire        _GEN_100889 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1790 & _GEN_100655 : _GEN_1008 ? ~_GEN_1790 & _GEN_100655 : ~(_GEN_100765 & _GEN_1790) & _GEN_100655) : _GEN_100655;
  wire        _GEN_100890 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1791 & _GEN_100656 : _GEN_1008 ? ~_GEN_1791 & _GEN_100656 : ~(_GEN_100765 & _GEN_1791) & _GEN_100656) : _GEN_100656;
  wire        _GEN_100891 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1792 & _GEN_100657 : _GEN_1008 ? ~_GEN_1792 & _GEN_100657 : ~(_GEN_100765 & _GEN_1792) & _GEN_100657) : _GEN_100657;
  wire        _GEN_100892 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1793 & _GEN_100658 : _GEN_1008 ? ~_GEN_1793 & _GEN_100658 : ~(_GEN_100765 & _GEN_1793) & _GEN_100658) : _GEN_100658;
  wire        _GEN_100893 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1794 & _GEN_100659 : _GEN_1008 ? ~_GEN_1794 & _GEN_100659 : ~(_GEN_100765 & _GEN_1794) & _GEN_100659) : _GEN_100659;
  wire        _GEN_100894 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1795 & _GEN_100660 : _GEN_1008 ? ~_GEN_1795 & _GEN_100660 : ~(_GEN_100765 & _GEN_1795) & _GEN_100660) : _GEN_100660;
  wire        _GEN_100895 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1796 & _GEN_100661 : _GEN_1008 ? ~_GEN_1796 & _GEN_100661 : ~(_GEN_100765 & _GEN_1796) & _GEN_100661) : _GEN_100661;
  wire        _GEN_100896 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1797 & _GEN_100662 : _GEN_1008 ? ~_GEN_1797 & _GEN_100662 : ~(_GEN_100765 & _GEN_1797) & _GEN_100662) : _GEN_100662;
  wire        _GEN_100897 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1798 & _GEN_100663 : _GEN_1008 ? ~_GEN_1798 & _GEN_100663 : ~(_GEN_100765 & _GEN_1798) & _GEN_100663) : _GEN_100663;
  wire        _GEN_100898 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1799 & _GEN_100664 : _GEN_1008 ? ~_GEN_1799 & _GEN_100664 : ~(_GEN_100765 & _GEN_1799) & _GEN_100664) : _GEN_100664;
  wire        _GEN_100899 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1800 & _GEN_100665 : _GEN_1008 ? ~_GEN_1800 & _GEN_100665 : ~(_GEN_100765 & _GEN_1800) & _GEN_100665) : _GEN_100665;
  wire        _GEN_100900 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1801 & _GEN_100666 : _GEN_1008 ? ~_GEN_1801 & _GEN_100666 : ~(_GEN_100765 & _GEN_1801) & _GEN_100666) : _GEN_100666;
  wire        _GEN_100901 = _GEN_1006 ? (_GEN_100834 ? ~_GEN_1802 & _GEN_100667 : _GEN_1008 ? ~_GEN_1802 & _GEN_100667 : ~(_GEN_100765 & _GEN_1802) & _GEN_100667) : _GEN_100667;
  wire        _GEN_100902 = _GEN_1006 ? (_GEN_100834 ? ~(&lcam_ldq_idx_1) & _GEN_100668 : _GEN_1008 ? ~(&lcam_ldq_idx_1) & _GEN_100668 : ~(_GEN_100765 & (&lcam_ldq_idx_1)) & _GEN_100668) : _GEN_100668;
  wire        _GEN_101105 = _GEN_1009 ? (_GEN_101068 ? (|lcam_ldq_idx_0) & _GEN_100871 : _GEN_1011 ? (|lcam_ldq_idx_0) & _GEN_100871 : ~(_GEN_101233 & ~(|lcam_ldq_idx_0)) & _GEN_100871) : _GEN_100871;
  wire        _GEN_101106 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1743 & _GEN_100872 : _GEN_1011 ? ~_GEN_1743 & _GEN_100872 : ~(_GEN_101233 & _GEN_1743) & _GEN_100872) : _GEN_100872;
  wire        _GEN_101107 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1744 & _GEN_100873 : _GEN_1011 ? ~_GEN_1744 & _GEN_100873 : ~(_GEN_101233 & _GEN_1744) & _GEN_100873) : _GEN_100873;
  wire        _GEN_101108 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1745 & _GEN_100874 : _GEN_1011 ? ~_GEN_1745 & _GEN_100874 : ~(_GEN_101233 & _GEN_1745) & _GEN_100874) : _GEN_100874;
  wire        _GEN_101109 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1746 & _GEN_100875 : _GEN_1011 ? ~_GEN_1746 & _GEN_100875 : ~(_GEN_101233 & _GEN_1746) & _GEN_100875) : _GEN_100875;
  wire        _GEN_101110 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1747 & _GEN_100876 : _GEN_1011 ? ~_GEN_1747 & _GEN_100876 : ~(_GEN_101233 & _GEN_1747) & _GEN_100876) : _GEN_100876;
  wire        _GEN_101111 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1748 & _GEN_100877 : _GEN_1011 ? ~_GEN_1748 & _GEN_100877 : ~(_GEN_101233 & _GEN_1748) & _GEN_100877) : _GEN_100877;
  wire        _GEN_101112 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1749 & _GEN_100878 : _GEN_1011 ? ~_GEN_1749 & _GEN_100878 : ~(_GEN_101233 & _GEN_1749) & _GEN_100878) : _GEN_100878;
  wire        _GEN_101113 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1750 & _GEN_100879 : _GEN_1011 ? ~_GEN_1750 & _GEN_100879 : ~(_GEN_101233 & _GEN_1750) & _GEN_100879) : _GEN_100879;
  wire        _GEN_101114 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1751 & _GEN_100880 : _GEN_1011 ? ~_GEN_1751 & _GEN_100880 : ~(_GEN_101233 & _GEN_1751) & _GEN_100880) : _GEN_100880;
  wire        _GEN_101115 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1752 & _GEN_100881 : _GEN_1011 ? ~_GEN_1752 & _GEN_100881 : ~(_GEN_101233 & _GEN_1752) & _GEN_100881) : _GEN_100881;
  wire        _GEN_101116 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1753 & _GEN_100882 : _GEN_1011 ? ~_GEN_1753 & _GEN_100882 : ~(_GEN_101233 & _GEN_1753) & _GEN_100882) : _GEN_100882;
  wire        _GEN_101117 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1754 & _GEN_100883 : _GEN_1011 ? ~_GEN_1754 & _GEN_100883 : ~(_GEN_101233 & _GEN_1754) & _GEN_100883) : _GEN_100883;
  wire        _GEN_101118 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1755 & _GEN_100884 : _GEN_1011 ? ~_GEN_1755 & _GEN_100884 : ~(_GEN_101233 & _GEN_1755) & _GEN_100884) : _GEN_100884;
  wire        _GEN_101119 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1756 & _GEN_100885 : _GEN_1011 ? ~_GEN_1756 & _GEN_100885 : ~(_GEN_101233 & _GEN_1756) & _GEN_100885) : _GEN_100885;
  wire        _GEN_101120 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1757 & _GEN_100886 : _GEN_1011 ? ~_GEN_1757 & _GEN_100886 : ~(_GEN_101233 & _GEN_1757) & _GEN_100886) : _GEN_100886;
  wire        _GEN_101121 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1758 & _GEN_100887 : _GEN_1011 ? ~_GEN_1758 & _GEN_100887 : ~(_GEN_101233 & _GEN_1758) & _GEN_100887) : _GEN_100887;
  wire        _GEN_101122 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1759 & _GEN_100888 : _GEN_1011 ? ~_GEN_1759 & _GEN_100888 : ~(_GEN_101233 & _GEN_1759) & _GEN_100888) : _GEN_100888;
  wire        _GEN_101123 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1760 & _GEN_100889 : _GEN_1011 ? ~_GEN_1760 & _GEN_100889 : ~(_GEN_101233 & _GEN_1760) & _GEN_100889) : _GEN_100889;
  wire        _GEN_101124 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1761 & _GEN_100890 : _GEN_1011 ? ~_GEN_1761 & _GEN_100890 : ~(_GEN_101233 & _GEN_1761) & _GEN_100890) : _GEN_100890;
  wire        _GEN_101125 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1762 & _GEN_100891 : _GEN_1011 ? ~_GEN_1762 & _GEN_100891 : ~(_GEN_101233 & _GEN_1762) & _GEN_100891) : _GEN_100891;
  wire        _GEN_101126 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1763 & _GEN_100892 : _GEN_1011 ? ~_GEN_1763 & _GEN_100892 : ~(_GEN_101233 & _GEN_1763) & _GEN_100892) : _GEN_100892;
  wire        _GEN_101127 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1764 & _GEN_100893 : _GEN_1011 ? ~_GEN_1764 & _GEN_100893 : ~(_GEN_101233 & _GEN_1764) & _GEN_100893) : _GEN_100893;
  wire        _GEN_101128 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1765 & _GEN_100894 : _GEN_1011 ? ~_GEN_1765 & _GEN_100894 : ~(_GEN_101233 & _GEN_1765) & _GEN_100894) : _GEN_100894;
  wire        _GEN_101129 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1766 & _GEN_100895 : _GEN_1011 ? ~_GEN_1766 & _GEN_100895 : ~(_GEN_101233 & _GEN_1766) & _GEN_100895) : _GEN_100895;
  wire        _GEN_101130 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1767 & _GEN_100896 : _GEN_1011 ? ~_GEN_1767 & _GEN_100896 : ~(_GEN_101233 & _GEN_1767) & _GEN_100896) : _GEN_100896;
  wire        _GEN_101131 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1768 & _GEN_100897 : _GEN_1011 ? ~_GEN_1768 & _GEN_100897 : ~(_GEN_101233 & _GEN_1768) & _GEN_100897) : _GEN_100897;
  wire        _GEN_101132 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1769 & _GEN_100898 : _GEN_1011 ? ~_GEN_1769 & _GEN_100898 : ~(_GEN_101233 & _GEN_1769) & _GEN_100898) : _GEN_100898;
  wire        _GEN_101133 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1770 & _GEN_100899 : _GEN_1011 ? ~_GEN_1770 & _GEN_100899 : ~(_GEN_101233 & _GEN_1770) & _GEN_100899) : _GEN_100899;
  wire        _GEN_101134 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1771 & _GEN_100900 : _GEN_1011 ? ~_GEN_1771 & _GEN_100900 : ~(_GEN_101233 & _GEN_1771) & _GEN_100900) : _GEN_100900;
  wire        _GEN_101135 = _GEN_1009 ? (_GEN_101068 ? ~_GEN_1772 & _GEN_100901 : _GEN_1011 ? ~_GEN_1772 & _GEN_100901 : ~(_GEN_101233 & _GEN_1772) & _GEN_100901) : _GEN_100901;
  wire        _GEN_101136 = _GEN_1009 ? (_GEN_101068 ? ~(&lcam_ldq_idx_0) & _GEN_100902 : _GEN_1011 ? ~(&lcam_ldq_idx_0) & _GEN_100902 : ~(_GEN_101233 & (&lcam_ldq_idx_0)) & _GEN_100902) : _GEN_100902;
  wire        _GEN_101339 = _GEN_1012 ? (_GEN_101302 ? (|lcam_ldq_idx_1) & _GEN_101105 : _GEN_1014 ? (|lcam_ldq_idx_1) & _GEN_101105 : ~(_GEN_101233 & ~(|lcam_ldq_idx_1)) & _GEN_101105) : _GEN_101105;
  wire        _GEN_101340 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1773 & _GEN_101106 : _GEN_1014 ? ~_GEN_1773 & _GEN_101106 : ~(_GEN_101233 & _GEN_1773) & _GEN_101106) : _GEN_101106;
  wire        _GEN_101341 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1774 & _GEN_101107 : _GEN_1014 ? ~_GEN_1774 & _GEN_101107 : ~(_GEN_101233 & _GEN_1774) & _GEN_101107) : _GEN_101107;
  wire        _GEN_101342 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1775 & _GEN_101108 : _GEN_1014 ? ~_GEN_1775 & _GEN_101108 : ~(_GEN_101233 & _GEN_1775) & _GEN_101108) : _GEN_101108;
  wire        _GEN_101343 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1776 & _GEN_101109 : _GEN_1014 ? ~_GEN_1776 & _GEN_101109 : ~(_GEN_101233 & _GEN_1776) & _GEN_101109) : _GEN_101109;
  wire        _GEN_101344 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1777 & _GEN_101110 : _GEN_1014 ? ~_GEN_1777 & _GEN_101110 : ~(_GEN_101233 & _GEN_1777) & _GEN_101110) : _GEN_101110;
  wire        _GEN_101345 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1778 & _GEN_101111 : _GEN_1014 ? ~_GEN_1778 & _GEN_101111 : ~(_GEN_101233 & _GEN_1778) & _GEN_101111) : _GEN_101111;
  wire        _GEN_101346 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1779 & _GEN_101112 : _GEN_1014 ? ~_GEN_1779 & _GEN_101112 : ~(_GEN_101233 & _GEN_1779) & _GEN_101112) : _GEN_101112;
  wire        _GEN_101347 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1780 & _GEN_101113 : _GEN_1014 ? ~_GEN_1780 & _GEN_101113 : ~(_GEN_101233 & _GEN_1780) & _GEN_101113) : _GEN_101113;
  wire        _GEN_101348 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1781 & _GEN_101114 : _GEN_1014 ? ~_GEN_1781 & _GEN_101114 : ~(_GEN_101233 & _GEN_1781) & _GEN_101114) : _GEN_101114;
  wire        _GEN_101349 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1782 & _GEN_101115 : _GEN_1014 ? ~_GEN_1782 & _GEN_101115 : ~(_GEN_101233 & _GEN_1782) & _GEN_101115) : _GEN_101115;
  wire        _GEN_101350 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1783 & _GEN_101116 : _GEN_1014 ? ~_GEN_1783 & _GEN_101116 : ~(_GEN_101233 & _GEN_1783) & _GEN_101116) : _GEN_101116;
  wire        _GEN_101351 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1784 & _GEN_101117 : _GEN_1014 ? ~_GEN_1784 & _GEN_101117 : ~(_GEN_101233 & _GEN_1784) & _GEN_101117) : _GEN_101117;
  wire        _GEN_101352 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1785 & _GEN_101118 : _GEN_1014 ? ~_GEN_1785 & _GEN_101118 : ~(_GEN_101233 & _GEN_1785) & _GEN_101118) : _GEN_101118;
  wire        _GEN_101353 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1786 & _GEN_101119 : _GEN_1014 ? ~_GEN_1786 & _GEN_101119 : ~(_GEN_101233 & _GEN_1786) & _GEN_101119) : _GEN_101119;
  wire        _GEN_101354 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1787 & _GEN_101120 : _GEN_1014 ? ~_GEN_1787 & _GEN_101120 : ~(_GEN_101233 & _GEN_1787) & _GEN_101120) : _GEN_101120;
  wire        _GEN_101355 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1788 & _GEN_101121 : _GEN_1014 ? ~_GEN_1788 & _GEN_101121 : ~(_GEN_101233 & _GEN_1788) & _GEN_101121) : _GEN_101121;
  wire        _GEN_101356 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1789 & _GEN_101122 : _GEN_1014 ? ~_GEN_1789 & _GEN_101122 : ~(_GEN_101233 & _GEN_1789) & _GEN_101122) : _GEN_101122;
  wire        _GEN_101357 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1790 & _GEN_101123 : _GEN_1014 ? ~_GEN_1790 & _GEN_101123 : ~(_GEN_101233 & _GEN_1790) & _GEN_101123) : _GEN_101123;
  wire        _GEN_101358 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1791 & _GEN_101124 : _GEN_1014 ? ~_GEN_1791 & _GEN_101124 : ~(_GEN_101233 & _GEN_1791) & _GEN_101124) : _GEN_101124;
  wire        _GEN_101359 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1792 & _GEN_101125 : _GEN_1014 ? ~_GEN_1792 & _GEN_101125 : ~(_GEN_101233 & _GEN_1792) & _GEN_101125) : _GEN_101125;
  wire        _GEN_101360 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1793 & _GEN_101126 : _GEN_1014 ? ~_GEN_1793 & _GEN_101126 : ~(_GEN_101233 & _GEN_1793) & _GEN_101126) : _GEN_101126;
  wire        _GEN_101361 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1794 & _GEN_101127 : _GEN_1014 ? ~_GEN_1794 & _GEN_101127 : ~(_GEN_101233 & _GEN_1794) & _GEN_101127) : _GEN_101127;
  wire        _GEN_101362 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1795 & _GEN_101128 : _GEN_1014 ? ~_GEN_1795 & _GEN_101128 : ~(_GEN_101233 & _GEN_1795) & _GEN_101128) : _GEN_101128;
  wire        _GEN_101363 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1796 & _GEN_101129 : _GEN_1014 ? ~_GEN_1796 & _GEN_101129 : ~(_GEN_101233 & _GEN_1796) & _GEN_101129) : _GEN_101129;
  wire        _GEN_101364 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1797 & _GEN_101130 : _GEN_1014 ? ~_GEN_1797 & _GEN_101130 : ~(_GEN_101233 & _GEN_1797) & _GEN_101130) : _GEN_101130;
  wire        _GEN_101365 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1798 & _GEN_101131 : _GEN_1014 ? ~_GEN_1798 & _GEN_101131 : ~(_GEN_101233 & _GEN_1798) & _GEN_101131) : _GEN_101131;
  wire        _GEN_101366 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1799 & _GEN_101132 : _GEN_1014 ? ~_GEN_1799 & _GEN_101132 : ~(_GEN_101233 & _GEN_1799) & _GEN_101132) : _GEN_101132;
  wire        _GEN_101367 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1800 & _GEN_101133 : _GEN_1014 ? ~_GEN_1800 & _GEN_101133 : ~(_GEN_101233 & _GEN_1800) & _GEN_101133) : _GEN_101133;
  wire        _GEN_101368 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1801 & _GEN_101134 : _GEN_1014 ? ~_GEN_1801 & _GEN_101134 : ~(_GEN_101233 & _GEN_1801) & _GEN_101134) : _GEN_101134;
  wire        _GEN_101369 = _GEN_1012 ? (_GEN_101302 ? ~_GEN_1802 & _GEN_101135 : _GEN_1014 ? ~_GEN_1802 & _GEN_101135 : ~(_GEN_101233 & _GEN_1802) & _GEN_101135) : _GEN_101135;
  wire        _GEN_101370 = _GEN_1012 ? (_GEN_101302 ? ~(&lcam_ldq_idx_1) & _GEN_101136 : _GEN_1014 ? ~(&lcam_ldq_idx_1) & _GEN_101136 : ~(_GEN_101233 & (&lcam_ldq_idx_1)) & _GEN_101136) : _GEN_101136;
  wire        _GEN_101573 = _GEN_1015 ? (_GEN_101536 ? (|lcam_ldq_idx_0) & _GEN_101339 : _GEN_1017 ? (|lcam_ldq_idx_0) & _GEN_101339 : ~(_GEN_101701 & ~(|lcam_ldq_idx_0)) & _GEN_101339) : _GEN_101339;
  wire        _GEN_101574 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1743 & _GEN_101340 : _GEN_1017 ? ~_GEN_1743 & _GEN_101340 : ~(_GEN_101701 & _GEN_1743) & _GEN_101340) : _GEN_101340;
  wire        _GEN_101575 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1744 & _GEN_101341 : _GEN_1017 ? ~_GEN_1744 & _GEN_101341 : ~(_GEN_101701 & _GEN_1744) & _GEN_101341) : _GEN_101341;
  wire        _GEN_101576 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1745 & _GEN_101342 : _GEN_1017 ? ~_GEN_1745 & _GEN_101342 : ~(_GEN_101701 & _GEN_1745) & _GEN_101342) : _GEN_101342;
  wire        _GEN_101577 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1746 & _GEN_101343 : _GEN_1017 ? ~_GEN_1746 & _GEN_101343 : ~(_GEN_101701 & _GEN_1746) & _GEN_101343) : _GEN_101343;
  wire        _GEN_101578 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1747 & _GEN_101344 : _GEN_1017 ? ~_GEN_1747 & _GEN_101344 : ~(_GEN_101701 & _GEN_1747) & _GEN_101344) : _GEN_101344;
  wire        _GEN_101579 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1748 & _GEN_101345 : _GEN_1017 ? ~_GEN_1748 & _GEN_101345 : ~(_GEN_101701 & _GEN_1748) & _GEN_101345) : _GEN_101345;
  wire        _GEN_101580 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1749 & _GEN_101346 : _GEN_1017 ? ~_GEN_1749 & _GEN_101346 : ~(_GEN_101701 & _GEN_1749) & _GEN_101346) : _GEN_101346;
  wire        _GEN_101581 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1750 & _GEN_101347 : _GEN_1017 ? ~_GEN_1750 & _GEN_101347 : ~(_GEN_101701 & _GEN_1750) & _GEN_101347) : _GEN_101347;
  wire        _GEN_101582 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1751 & _GEN_101348 : _GEN_1017 ? ~_GEN_1751 & _GEN_101348 : ~(_GEN_101701 & _GEN_1751) & _GEN_101348) : _GEN_101348;
  wire        _GEN_101583 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1752 & _GEN_101349 : _GEN_1017 ? ~_GEN_1752 & _GEN_101349 : ~(_GEN_101701 & _GEN_1752) & _GEN_101349) : _GEN_101349;
  wire        _GEN_101584 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1753 & _GEN_101350 : _GEN_1017 ? ~_GEN_1753 & _GEN_101350 : ~(_GEN_101701 & _GEN_1753) & _GEN_101350) : _GEN_101350;
  wire        _GEN_101585 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1754 & _GEN_101351 : _GEN_1017 ? ~_GEN_1754 & _GEN_101351 : ~(_GEN_101701 & _GEN_1754) & _GEN_101351) : _GEN_101351;
  wire        _GEN_101586 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1755 & _GEN_101352 : _GEN_1017 ? ~_GEN_1755 & _GEN_101352 : ~(_GEN_101701 & _GEN_1755) & _GEN_101352) : _GEN_101352;
  wire        _GEN_101587 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1756 & _GEN_101353 : _GEN_1017 ? ~_GEN_1756 & _GEN_101353 : ~(_GEN_101701 & _GEN_1756) & _GEN_101353) : _GEN_101353;
  wire        _GEN_101588 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1757 & _GEN_101354 : _GEN_1017 ? ~_GEN_1757 & _GEN_101354 : ~(_GEN_101701 & _GEN_1757) & _GEN_101354) : _GEN_101354;
  wire        _GEN_101589 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1758 & _GEN_101355 : _GEN_1017 ? ~_GEN_1758 & _GEN_101355 : ~(_GEN_101701 & _GEN_1758) & _GEN_101355) : _GEN_101355;
  wire        _GEN_101590 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1759 & _GEN_101356 : _GEN_1017 ? ~_GEN_1759 & _GEN_101356 : ~(_GEN_101701 & _GEN_1759) & _GEN_101356) : _GEN_101356;
  wire        _GEN_101591 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1760 & _GEN_101357 : _GEN_1017 ? ~_GEN_1760 & _GEN_101357 : ~(_GEN_101701 & _GEN_1760) & _GEN_101357) : _GEN_101357;
  wire        _GEN_101592 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1761 & _GEN_101358 : _GEN_1017 ? ~_GEN_1761 & _GEN_101358 : ~(_GEN_101701 & _GEN_1761) & _GEN_101358) : _GEN_101358;
  wire        _GEN_101593 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1762 & _GEN_101359 : _GEN_1017 ? ~_GEN_1762 & _GEN_101359 : ~(_GEN_101701 & _GEN_1762) & _GEN_101359) : _GEN_101359;
  wire        _GEN_101594 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1763 & _GEN_101360 : _GEN_1017 ? ~_GEN_1763 & _GEN_101360 : ~(_GEN_101701 & _GEN_1763) & _GEN_101360) : _GEN_101360;
  wire        _GEN_101595 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1764 & _GEN_101361 : _GEN_1017 ? ~_GEN_1764 & _GEN_101361 : ~(_GEN_101701 & _GEN_1764) & _GEN_101361) : _GEN_101361;
  wire        _GEN_101596 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1765 & _GEN_101362 : _GEN_1017 ? ~_GEN_1765 & _GEN_101362 : ~(_GEN_101701 & _GEN_1765) & _GEN_101362) : _GEN_101362;
  wire        _GEN_101597 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1766 & _GEN_101363 : _GEN_1017 ? ~_GEN_1766 & _GEN_101363 : ~(_GEN_101701 & _GEN_1766) & _GEN_101363) : _GEN_101363;
  wire        _GEN_101598 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1767 & _GEN_101364 : _GEN_1017 ? ~_GEN_1767 & _GEN_101364 : ~(_GEN_101701 & _GEN_1767) & _GEN_101364) : _GEN_101364;
  wire        _GEN_101599 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1768 & _GEN_101365 : _GEN_1017 ? ~_GEN_1768 & _GEN_101365 : ~(_GEN_101701 & _GEN_1768) & _GEN_101365) : _GEN_101365;
  wire        _GEN_101600 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1769 & _GEN_101366 : _GEN_1017 ? ~_GEN_1769 & _GEN_101366 : ~(_GEN_101701 & _GEN_1769) & _GEN_101366) : _GEN_101366;
  wire        _GEN_101601 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1770 & _GEN_101367 : _GEN_1017 ? ~_GEN_1770 & _GEN_101367 : ~(_GEN_101701 & _GEN_1770) & _GEN_101367) : _GEN_101367;
  wire        _GEN_101602 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1771 & _GEN_101368 : _GEN_1017 ? ~_GEN_1771 & _GEN_101368 : ~(_GEN_101701 & _GEN_1771) & _GEN_101368) : _GEN_101368;
  wire        _GEN_101603 = _GEN_1015 ? (_GEN_101536 ? ~_GEN_1772 & _GEN_101369 : _GEN_1017 ? ~_GEN_1772 & _GEN_101369 : ~(_GEN_101701 & _GEN_1772) & _GEN_101369) : _GEN_101369;
  wire        _GEN_101604 = _GEN_1015 ? (_GEN_101536 ? ~(&lcam_ldq_idx_0) & _GEN_101370 : _GEN_1017 ? ~(&lcam_ldq_idx_0) & _GEN_101370 : ~(_GEN_101701 & (&lcam_ldq_idx_0)) & _GEN_101370) : _GEN_101370;
  wire        _GEN_101807 = _GEN_1018 ? (_GEN_101770 ? (|lcam_ldq_idx_1) & _GEN_101573 : _GEN_1020 ? (|lcam_ldq_idx_1) & _GEN_101573 : ~(_GEN_101701 & ~(|lcam_ldq_idx_1)) & _GEN_101573) : _GEN_101573;
  wire        _GEN_101808 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1773 & _GEN_101574 : _GEN_1020 ? ~_GEN_1773 & _GEN_101574 : ~(_GEN_101701 & _GEN_1773) & _GEN_101574) : _GEN_101574;
  wire        _GEN_101809 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1774 & _GEN_101575 : _GEN_1020 ? ~_GEN_1774 & _GEN_101575 : ~(_GEN_101701 & _GEN_1774) & _GEN_101575) : _GEN_101575;
  wire        _GEN_101810 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1775 & _GEN_101576 : _GEN_1020 ? ~_GEN_1775 & _GEN_101576 : ~(_GEN_101701 & _GEN_1775) & _GEN_101576) : _GEN_101576;
  wire        _GEN_101811 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1776 & _GEN_101577 : _GEN_1020 ? ~_GEN_1776 & _GEN_101577 : ~(_GEN_101701 & _GEN_1776) & _GEN_101577) : _GEN_101577;
  wire        _GEN_101812 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1777 & _GEN_101578 : _GEN_1020 ? ~_GEN_1777 & _GEN_101578 : ~(_GEN_101701 & _GEN_1777) & _GEN_101578) : _GEN_101578;
  wire        _GEN_101813 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1778 & _GEN_101579 : _GEN_1020 ? ~_GEN_1778 & _GEN_101579 : ~(_GEN_101701 & _GEN_1778) & _GEN_101579) : _GEN_101579;
  wire        _GEN_101814 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1779 & _GEN_101580 : _GEN_1020 ? ~_GEN_1779 & _GEN_101580 : ~(_GEN_101701 & _GEN_1779) & _GEN_101580) : _GEN_101580;
  wire        _GEN_101815 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1780 & _GEN_101581 : _GEN_1020 ? ~_GEN_1780 & _GEN_101581 : ~(_GEN_101701 & _GEN_1780) & _GEN_101581) : _GEN_101581;
  wire        _GEN_101816 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1781 & _GEN_101582 : _GEN_1020 ? ~_GEN_1781 & _GEN_101582 : ~(_GEN_101701 & _GEN_1781) & _GEN_101582) : _GEN_101582;
  wire        _GEN_101817 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1782 & _GEN_101583 : _GEN_1020 ? ~_GEN_1782 & _GEN_101583 : ~(_GEN_101701 & _GEN_1782) & _GEN_101583) : _GEN_101583;
  wire        _GEN_101818 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1783 & _GEN_101584 : _GEN_1020 ? ~_GEN_1783 & _GEN_101584 : ~(_GEN_101701 & _GEN_1783) & _GEN_101584) : _GEN_101584;
  wire        _GEN_101819 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1784 & _GEN_101585 : _GEN_1020 ? ~_GEN_1784 & _GEN_101585 : ~(_GEN_101701 & _GEN_1784) & _GEN_101585) : _GEN_101585;
  wire        _GEN_101820 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1785 & _GEN_101586 : _GEN_1020 ? ~_GEN_1785 & _GEN_101586 : ~(_GEN_101701 & _GEN_1785) & _GEN_101586) : _GEN_101586;
  wire        _GEN_101821 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1786 & _GEN_101587 : _GEN_1020 ? ~_GEN_1786 & _GEN_101587 : ~(_GEN_101701 & _GEN_1786) & _GEN_101587) : _GEN_101587;
  wire        _GEN_101822 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1787 & _GEN_101588 : _GEN_1020 ? ~_GEN_1787 & _GEN_101588 : ~(_GEN_101701 & _GEN_1787) & _GEN_101588) : _GEN_101588;
  wire        _GEN_101823 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1788 & _GEN_101589 : _GEN_1020 ? ~_GEN_1788 & _GEN_101589 : ~(_GEN_101701 & _GEN_1788) & _GEN_101589) : _GEN_101589;
  wire        _GEN_101824 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1789 & _GEN_101590 : _GEN_1020 ? ~_GEN_1789 & _GEN_101590 : ~(_GEN_101701 & _GEN_1789) & _GEN_101590) : _GEN_101590;
  wire        _GEN_101825 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1790 & _GEN_101591 : _GEN_1020 ? ~_GEN_1790 & _GEN_101591 : ~(_GEN_101701 & _GEN_1790) & _GEN_101591) : _GEN_101591;
  wire        _GEN_101826 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1791 & _GEN_101592 : _GEN_1020 ? ~_GEN_1791 & _GEN_101592 : ~(_GEN_101701 & _GEN_1791) & _GEN_101592) : _GEN_101592;
  wire        _GEN_101827 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1792 & _GEN_101593 : _GEN_1020 ? ~_GEN_1792 & _GEN_101593 : ~(_GEN_101701 & _GEN_1792) & _GEN_101593) : _GEN_101593;
  wire        _GEN_101828 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1793 & _GEN_101594 : _GEN_1020 ? ~_GEN_1793 & _GEN_101594 : ~(_GEN_101701 & _GEN_1793) & _GEN_101594) : _GEN_101594;
  wire        _GEN_101829 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1794 & _GEN_101595 : _GEN_1020 ? ~_GEN_1794 & _GEN_101595 : ~(_GEN_101701 & _GEN_1794) & _GEN_101595) : _GEN_101595;
  wire        _GEN_101830 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1795 & _GEN_101596 : _GEN_1020 ? ~_GEN_1795 & _GEN_101596 : ~(_GEN_101701 & _GEN_1795) & _GEN_101596) : _GEN_101596;
  wire        _GEN_101831 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1796 & _GEN_101597 : _GEN_1020 ? ~_GEN_1796 & _GEN_101597 : ~(_GEN_101701 & _GEN_1796) & _GEN_101597) : _GEN_101597;
  wire        _GEN_101832 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1797 & _GEN_101598 : _GEN_1020 ? ~_GEN_1797 & _GEN_101598 : ~(_GEN_101701 & _GEN_1797) & _GEN_101598) : _GEN_101598;
  wire        _GEN_101833 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1798 & _GEN_101599 : _GEN_1020 ? ~_GEN_1798 & _GEN_101599 : ~(_GEN_101701 & _GEN_1798) & _GEN_101599) : _GEN_101599;
  wire        _GEN_101834 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1799 & _GEN_101600 : _GEN_1020 ? ~_GEN_1799 & _GEN_101600 : ~(_GEN_101701 & _GEN_1799) & _GEN_101600) : _GEN_101600;
  wire        _GEN_101835 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1800 & _GEN_101601 : _GEN_1020 ? ~_GEN_1800 & _GEN_101601 : ~(_GEN_101701 & _GEN_1800) & _GEN_101601) : _GEN_101601;
  wire        _GEN_101836 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1801 & _GEN_101602 : _GEN_1020 ? ~_GEN_1801 & _GEN_101602 : ~(_GEN_101701 & _GEN_1801) & _GEN_101602) : _GEN_101602;
  wire        _GEN_101837 = _GEN_1018 ? (_GEN_101770 ? ~_GEN_1802 & _GEN_101603 : _GEN_1020 ? ~_GEN_1802 & _GEN_101603 : ~(_GEN_101701 & _GEN_1802) & _GEN_101603) : _GEN_101603;
  wire        _GEN_101838 = _GEN_1018 ? (_GEN_101770 ? ~(&lcam_ldq_idx_1) & _GEN_101604 : _GEN_1020 ? ~(&lcam_ldq_idx_1) & _GEN_101604 : ~(_GEN_101701 & (&lcam_ldq_idx_1)) & _GEN_101604) : _GEN_101604;
  wire        _GEN_102041 = _GEN_1021 ? (_GEN_102004 ? (|lcam_ldq_idx_0) & _GEN_101807 : _GEN_1023 ? (|lcam_ldq_idx_0) & _GEN_101807 : ~(_GEN_102169 & ~(|lcam_ldq_idx_0)) & _GEN_101807) : _GEN_101807;
  wire        _GEN_102042 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1743 & _GEN_101808 : _GEN_1023 ? ~_GEN_1743 & _GEN_101808 : ~(_GEN_102169 & _GEN_1743) & _GEN_101808) : _GEN_101808;
  wire        _GEN_102043 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1744 & _GEN_101809 : _GEN_1023 ? ~_GEN_1744 & _GEN_101809 : ~(_GEN_102169 & _GEN_1744) & _GEN_101809) : _GEN_101809;
  wire        _GEN_102044 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1745 & _GEN_101810 : _GEN_1023 ? ~_GEN_1745 & _GEN_101810 : ~(_GEN_102169 & _GEN_1745) & _GEN_101810) : _GEN_101810;
  wire        _GEN_102045 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1746 & _GEN_101811 : _GEN_1023 ? ~_GEN_1746 & _GEN_101811 : ~(_GEN_102169 & _GEN_1746) & _GEN_101811) : _GEN_101811;
  wire        _GEN_102046 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1747 & _GEN_101812 : _GEN_1023 ? ~_GEN_1747 & _GEN_101812 : ~(_GEN_102169 & _GEN_1747) & _GEN_101812) : _GEN_101812;
  wire        _GEN_102047 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1748 & _GEN_101813 : _GEN_1023 ? ~_GEN_1748 & _GEN_101813 : ~(_GEN_102169 & _GEN_1748) & _GEN_101813) : _GEN_101813;
  wire        _GEN_102048 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1749 & _GEN_101814 : _GEN_1023 ? ~_GEN_1749 & _GEN_101814 : ~(_GEN_102169 & _GEN_1749) & _GEN_101814) : _GEN_101814;
  wire        _GEN_102049 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1750 & _GEN_101815 : _GEN_1023 ? ~_GEN_1750 & _GEN_101815 : ~(_GEN_102169 & _GEN_1750) & _GEN_101815) : _GEN_101815;
  wire        _GEN_102050 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1751 & _GEN_101816 : _GEN_1023 ? ~_GEN_1751 & _GEN_101816 : ~(_GEN_102169 & _GEN_1751) & _GEN_101816) : _GEN_101816;
  wire        _GEN_102051 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1752 & _GEN_101817 : _GEN_1023 ? ~_GEN_1752 & _GEN_101817 : ~(_GEN_102169 & _GEN_1752) & _GEN_101817) : _GEN_101817;
  wire        _GEN_102052 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1753 & _GEN_101818 : _GEN_1023 ? ~_GEN_1753 & _GEN_101818 : ~(_GEN_102169 & _GEN_1753) & _GEN_101818) : _GEN_101818;
  wire        _GEN_102053 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1754 & _GEN_101819 : _GEN_1023 ? ~_GEN_1754 & _GEN_101819 : ~(_GEN_102169 & _GEN_1754) & _GEN_101819) : _GEN_101819;
  wire        _GEN_102054 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1755 & _GEN_101820 : _GEN_1023 ? ~_GEN_1755 & _GEN_101820 : ~(_GEN_102169 & _GEN_1755) & _GEN_101820) : _GEN_101820;
  wire        _GEN_102055 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1756 & _GEN_101821 : _GEN_1023 ? ~_GEN_1756 & _GEN_101821 : ~(_GEN_102169 & _GEN_1756) & _GEN_101821) : _GEN_101821;
  wire        _GEN_102056 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1757 & _GEN_101822 : _GEN_1023 ? ~_GEN_1757 & _GEN_101822 : ~(_GEN_102169 & _GEN_1757) & _GEN_101822) : _GEN_101822;
  wire        _GEN_102057 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1758 & _GEN_101823 : _GEN_1023 ? ~_GEN_1758 & _GEN_101823 : ~(_GEN_102169 & _GEN_1758) & _GEN_101823) : _GEN_101823;
  wire        _GEN_102058 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1759 & _GEN_101824 : _GEN_1023 ? ~_GEN_1759 & _GEN_101824 : ~(_GEN_102169 & _GEN_1759) & _GEN_101824) : _GEN_101824;
  wire        _GEN_102059 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1760 & _GEN_101825 : _GEN_1023 ? ~_GEN_1760 & _GEN_101825 : ~(_GEN_102169 & _GEN_1760) & _GEN_101825) : _GEN_101825;
  wire        _GEN_102060 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1761 & _GEN_101826 : _GEN_1023 ? ~_GEN_1761 & _GEN_101826 : ~(_GEN_102169 & _GEN_1761) & _GEN_101826) : _GEN_101826;
  wire        _GEN_102061 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1762 & _GEN_101827 : _GEN_1023 ? ~_GEN_1762 & _GEN_101827 : ~(_GEN_102169 & _GEN_1762) & _GEN_101827) : _GEN_101827;
  wire        _GEN_102062 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1763 & _GEN_101828 : _GEN_1023 ? ~_GEN_1763 & _GEN_101828 : ~(_GEN_102169 & _GEN_1763) & _GEN_101828) : _GEN_101828;
  wire        _GEN_102063 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1764 & _GEN_101829 : _GEN_1023 ? ~_GEN_1764 & _GEN_101829 : ~(_GEN_102169 & _GEN_1764) & _GEN_101829) : _GEN_101829;
  wire        _GEN_102064 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1765 & _GEN_101830 : _GEN_1023 ? ~_GEN_1765 & _GEN_101830 : ~(_GEN_102169 & _GEN_1765) & _GEN_101830) : _GEN_101830;
  wire        _GEN_102065 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1766 & _GEN_101831 : _GEN_1023 ? ~_GEN_1766 & _GEN_101831 : ~(_GEN_102169 & _GEN_1766) & _GEN_101831) : _GEN_101831;
  wire        _GEN_102066 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1767 & _GEN_101832 : _GEN_1023 ? ~_GEN_1767 & _GEN_101832 : ~(_GEN_102169 & _GEN_1767) & _GEN_101832) : _GEN_101832;
  wire        _GEN_102067 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1768 & _GEN_101833 : _GEN_1023 ? ~_GEN_1768 & _GEN_101833 : ~(_GEN_102169 & _GEN_1768) & _GEN_101833) : _GEN_101833;
  wire        _GEN_102068 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1769 & _GEN_101834 : _GEN_1023 ? ~_GEN_1769 & _GEN_101834 : ~(_GEN_102169 & _GEN_1769) & _GEN_101834) : _GEN_101834;
  wire        _GEN_102069 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1770 & _GEN_101835 : _GEN_1023 ? ~_GEN_1770 & _GEN_101835 : ~(_GEN_102169 & _GEN_1770) & _GEN_101835) : _GEN_101835;
  wire        _GEN_102070 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1771 & _GEN_101836 : _GEN_1023 ? ~_GEN_1771 & _GEN_101836 : ~(_GEN_102169 & _GEN_1771) & _GEN_101836) : _GEN_101836;
  wire        _GEN_102071 = _GEN_1021 ? (_GEN_102004 ? ~_GEN_1772 & _GEN_101837 : _GEN_1023 ? ~_GEN_1772 & _GEN_101837 : ~(_GEN_102169 & _GEN_1772) & _GEN_101837) : _GEN_101837;
  wire        _GEN_102072 = _GEN_1021 ? (_GEN_102004 ? ~(&lcam_ldq_idx_0) & _GEN_101838 : _GEN_1023 ? ~(&lcam_ldq_idx_0) & _GEN_101838 : ~(_GEN_102169 & (&lcam_ldq_idx_0)) & _GEN_101838) : _GEN_101838;
  wire        _GEN_102275 = _GEN_1024 ? (_GEN_102238 ? (|lcam_ldq_idx_1) & _GEN_102041 : _GEN_1026 ? (|lcam_ldq_idx_1) & _GEN_102041 : ~(_GEN_102169 & ~(|lcam_ldq_idx_1)) & _GEN_102041) : _GEN_102041;
  wire        _GEN_102276 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1773 & _GEN_102042 : _GEN_1026 ? ~_GEN_1773 & _GEN_102042 : ~(_GEN_102169 & _GEN_1773) & _GEN_102042) : _GEN_102042;
  wire        _GEN_102277 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1774 & _GEN_102043 : _GEN_1026 ? ~_GEN_1774 & _GEN_102043 : ~(_GEN_102169 & _GEN_1774) & _GEN_102043) : _GEN_102043;
  wire        _GEN_102278 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1775 & _GEN_102044 : _GEN_1026 ? ~_GEN_1775 & _GEN_102044 : ~(_GEN_102169 & _GEN_1775) & _GEN_102044) : _GEN_102044;
  wire        _GEN_102279 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1776 & _GEN_102045 : _GEN_1026 ? ~_GEN_1776 & _GEN_102045 : ~(_GEN_102169 & _GEN_1776) & _GEN_102045) : _GEN_102045;
  wire        _GEN_102280 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1777 & _GEN_102046 : _GEN_1026 ? ~_GEN_1777 & _GEN_102046 : ~(_GEN_102169 & _GEN_1777) & _GEN_102046) : _GEN_102046;
  wire        _GEN_102281 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1778 & _GEN_102047 : _GEN_1026 ? ~_GEN_1778 & _GEN_102047 : ~(_GEN_102169 & _GEN_1778) & _GEN_102047) : _GEN_102047;
  wire        _GEN_102282 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1779 & _GEN_102048 : _GEN_1026 ? ~_GEN_1779 & _GEN_102048 : ~(_GEN_102169 & _GEN_1779) & _GEN_102048) : _GEN_102048;
  wire        _GEN_102283 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1780 & _GEN_102049 : _GEN_1026 ? ~_GEN_1780 & _GEN_102049 : ~(_GEN_102169 & _GEN_1780) & _GEN_102049) : _GEN_102049;
  wire        _GEN_102284 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1781 & _GEN_102050 : _GEN_1026 ? ~_GEN_1781 & _GEN_102050 : ~(_GEN_102169 & _GEN_1781) & _GEN_102050) : _GEN_102050;
  wire        _GEN_102285 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1782 & _GEN_102051 : _GEN_1026 ? ~_GEN_1782 & _GEN_102051 : ~(_GEN_102169 & _GEN_1782) & _GEN_102051) : _GEN_102051;
  wire        _GEN_102286 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1783 & _GEN_102052 : _GEN_1026 ? ~_GEN_1783 & _GEN_102052 : ~(_GEN_102169 & _GEN_1783) & _GEN_102052) : _GEN_102052;
  wire        _GEN_102287 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1784 & _GEN_102053 : _GEN_1026 ? ~_GEN_1784 & _GEN_102053 : ~(_GEN_102169 & _GEN_1784) & _GEN_102053) : _GEN_102053;
  wire        _GEN_102288 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1785 & _GEN_102054 : _GEN_1026 ? ~_GEN_1785 & _GEN_102054 : ~(_GEN_102169 & _GEN_1785) & _GEN_102054) : _GEN_102054;
  wire        _GEN_102289 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1786 & _GEN_102055 : _GEN_1026 ? ~_GEN_1786 & _GEN_102055 : ~(_GEN_102169 & _GEN_1786) & _GEN_102055) : _GEN_102055;
  wire        _GEN_102290 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1787 & _GEN_102056 : _GEN_1026 ? ~_GEN_1787 & _GEN_102056 : ~(_GEN_102169 & _GEN_1787) & _GEN_102056) : _GEN_102056;
  wire        _GEN_102291 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1788 & _GEN_102057 : _GEN_1026 ? ~_GEN_1788 & _GEN_102057 : ~(_GEN_102169 & _GEN_1788) & _GEN_102057) : _GEN_102057;
  wire        _GEN_102292 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1789 & _GEN_102058 : _GEN_1026 ? ~_GEN_1789 & _GEN_102058 : ~(_GEN_102169 & _GEN_1789) & _GEN_102058) : _GEN_102058;
  wire        _GEN_102293 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1790 & _GEN_102059 : _GEN_1026 ? ~_GEN_1790 & _GEN_102059 : ~(_GEN_102169 & _GEN_1790) & _GEN_102059) : _GEN_102059;
  wire        _GEN_102294 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1791 & _GEN_102060 : _GEN_1026 ? ~_GEN_1791 & _GEN_102060 : ~(_GEN_102169 & _GEN_1791) & _GEN_102060) : _GEN_102060;
  wire        _GEN_102295 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1792 & _GEN_102061 : _GEN_1026 ? ~_GEN_1792 & _GEN_102061 : ~(_GEN_102169 & _GEN_1792) & _GEN_102061) : _GEN_102061;
  wire        _GEN_102296 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1793 & _GEN_102062 : _GEN_1026 ? ~_GEN_1793 & _GEN_102062 : ~(_GEN_102169 & _GEN_1793) & _GEN_102062) : _GEN_102062;
  wire        _GEN_102297 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1794 & _GEN_102063 : _GEN_1026 ? ~_GEN_1794 & _GEN_102063 : ~(_GEN_102169 & _GEN_1794) & _GEN_102063) : _GEN_102063;
  wire        _GEN_102298 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1795 & _GEN_102064 : _GEN_1026 ? ~_GEN_1795 & _GEN_102064 : ~(_GEN_102169 & _GEN_1795) & _GEN_102064) : _GEN_102064;
  wire        _GEN_102299 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1796 & _GEN_102065 : _GEN_1026 ? ~_GEN_1796 & _GEN_102065 : ~(_GEN_102169 & _GEN_1796) & _GEN_102065) : _GEN_102065;
  wire        _GEN_102300 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1797 & _GEN_102066 : _GEN_1026 ? ~_GEN_1797 & _GEN_102066 : ~(_GEN_102169 & _GEN_1797) & _GEN_102066) : _GEN_102066;
  wire        _GEN_102301 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1798 & _GEN_102067 : _GEN_1026 ? ~_GEN_1798 & _GEN_102067 : ~(_GEN_102169 & _GEN_1798) & _GEN_102067) : _GEN_102067;
  wire        _GEN_102302 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1799 & _GEN_102068 : _GEN_1026 ? ~_GEN_1799 & _GEN_102068 : ~(_GEN_102169 & _GEN_1799) & _GEN_102068) : _GEN_102068;
  wire        _GEN_102303 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1800 & _GEN_102069 : _GEN_1026 ? ~_GEN_1800 & _GEN_102069 : ~(_GEN_102169 & _GEN_1800) & _GEN_102069) : _GEN_102069;
  wire        _GEN_102304 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1801 & _GEN_102070 : _GEN_1026 ? ~_GEN_1801 & _GEN_102070 : ~(_GEN_102169 & _GEN_1801) & _GEN_102070) : _GEN_102070;
  wire        _GEN_102305 = _GEN_1024 ? (_GEN_102238 ? ~_GEN_1802 & _GEN_102071 : _GEN_1026 ? ~_GEN_1802 & _GEN_102071 : ~(_GEN_102169 & _GEN_1802) & _GEN_102071) : _GEN_102071;
  wire        _GEN_102306 = _GEN_1024 ? (_GEN_102238 ? ~(&lcam_ldq_idx_1) & _GEN_102072 : _GEN_1026 ? ~(&lcam_ldq_idx_1) & _GEN_102072 : ~(_GEN_102169 & (&lcam_ldq_idx_1)) & _GEN_102072) : _GEN_102072;
  wire        _GEN_102509 = _GEN_1027 ? (_GEN_102472 ? (|lcam_ldq_idx_0) & _GEN_102275 : _GEN_1029 ? (|lcam_ldq_idx_0) & _GEN_102275 : ~(_GEN_102637 & ~(|lcam_ldq_idx_0)) & _GEN_102275) : _GEN_102275;
  wire        _GEN_102510 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1743 & _GEN_102276 : _GEN_1029 ? ~_GEN_1743 & _GEN_102276 : ~(_GEN_102637 & _GEN_1743) & _GEN_102276) : _GEN_102276;
  wire        _GEN_102511 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1744 & _GEN_102277 : _GEN_1029 ? ~_GEN_1744 & _GEN_102277 : ~(_GEN_102637 & _GEN_1744) & _GEN_102277) : _GEN_102277;
  wire        _GEN_102512 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1745 & _GEN_102278 : _GEN_1029 ? ~_GEN_1745 & _GEN_102278 : ~(_GEN_102637 & _GEN_1745) & _GEN_102278) : _GEN_102278;
  wire        _GEN_102513 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1746 & _GEN_102279 : _GEN_1029 ? ~_GEN_1746 & _GEN_102279 : ~(_GEN_102637 & _GEN_1746) & _GEN_102279) : _GEN_102279;
  wire        _GEN_102514 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1747 & _GEN_102280 : _GEN_1029 ? ~_GEN_1747 & _GEN_102280 : ~(_GEN_102637 & _GEN_1747) & _GEN_102280) : _GEN_102280;
  wire        _GEN_102515 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1748 & _GEN_102281 : _GEN_1029 ? ~_GEN_1748 & _GEN_102281 : ~(_GEN_102637 & _GEN_1748) & _GEN_102281) : _GEN_102281;
  wire        _GEN_102516 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1749 & _GEN_102282 : _GEN_1029 ? ~_GEN_1749 & _GEN_102282 : ~(_GEN_102637 & _GEN_1749) & _GEN_102282) : _GEN_102282;
  wire        _GEN_102517 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1750 & _GEN_102283 : _GEN_1029 ? ~_GEN_1750 & _GEN_102283 : ~(_GEN_102637 & _GEN_1750) & _GEN_102283) : _GEN_102283;
  wire        _GEN_102518 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1751 & _GEN_102284 : _GEN_1029 ? ~_GEN_1751 & _GEN_102284 : ~(_GEN_102637 & _GEN_1751) & _GEN_102284) : _GEN_102284;
  wire        _GEN_102519 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1752 & _GEN_102285 : _GEN_1029 ? ~_GEN_1752 & _GEN_102285 : ~(_GEN_102637 & _GEN_1752) & _GEN_102285) : _GEN_102285;
  wire        _GEN_102520 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1753 & _GEN_102286 : _GEN_1029 ? ~_GEN_1753 & _GEN_102286 : ~(_GEN_102637 & _GEN_1753) & _GEN_102286) : _GEN_102286;
  wire        _GEN_102521 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1754 & _GEN_102287 : _GEN_1029 ? ~_GEN_1754 & _GEN_102287 : ~(_GEN_102637 & _GEN_1754) & _GEN_102287) : _GEN_102287;
  wire        _GEN_102522 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1755 & _GEN_102288 : _GEN_1029 ? ~_GEN_1755 & _GEN_102288 : ~(_GEN_102637 & _GEN_1755) & _GEN_102288) : _GEN_102288;
  wire        _GEN_102523 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1756 & _GEN_102289 : _GEN_1029 ? ~_GEN_1756 & _GEN_102289 : ~(_GEN_102637 & _GEN_1756) & _GEN_102289) : _GEN_102289;
  wire        _GEN_102524 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1757 & _GEN_102290 : _GEN_1029 ? ~_GEN_1757 & _GEN_102290 : ~(_GEN_102637 & _GEN_1757) & _GEN_102290) : _GEN_102290;
  wire        _GEN_102525 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1758 & _GEN_102291 : _GEN_1029 ? ~_GEN_1758 & _GEN_102291 : ~(_GEN_102637 & _GEN_1758) & _GEN_102291) : _GEN_102291;
  wire        _GEN_102526 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1759 & _GEN_102292 : _GEN_1029 ? ~_GEN_1759 & _GEN_102292 : ~(_GEN_102637 & _GEN_1759) & _GEN_102292) : _GEN_102292;
  wire        _GEN_102527 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1760 & _GEN_102293 : _GEN_1029 ? ~_GEN_1760 & _GEN_102293 : ~(_GEN_102637 & _GEN_1760) & _GEN_102293) : _GEN_102293;
  wire        _GEN_102528 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1761 & _GEN_102294 : _GEN_1029 ? ~_GEN_1761 & _GEN_102294 : ~(_GEN_102637 & _GEN_1761) & _GEN_102294) : _GEN_102294;
  wire        _GEN_102529 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1762 & _GEN_102295 : _GEN_1029 ? ~_GEN_1762 & _GEN_102295 : ~(_GEN_102637 & _GEN_1762) & _GEN_102295) : _GEN_102295;
  wire        _GEN_102530 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1763 & _GEN_102296 : _GEN_1029 ? ~_GEN_1763 & _GEN_102296 : ~(_GEN_102637 & _GEN_1763) & _GEN_102296) : _GEN_102296;
  wire        _GEN_102531 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1764 & _GEN_102297 : _GEN_1029 ? ~_GEN_1764 & _GEN_102297 : ~(_GEN_102637 & _GEN_1764) & _GEN_102297) : _GEN_102297;
  wire        _GEN_102532 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1765 & _GEN_102298 : _GEN_1029 ? ~_GEN_1765 & _GEN_102298 : ~(_GEN_102637 & _GEN_1765) & _GEN_102298) : _GEN_102298;
  wire        _GEN_102533 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1766 & _GEN_102299 : _GEN_1029 ? ~_GEN_1766 & _GEN_102299 : ~(_GEN_102637 & _GEN_1766) & _GEN_102299) : _GEN_102299;
  wire        _GEN_102534 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1767 & _GEN_102300 : _GEN_1029 ? ~_GEN_1767 & _GEN_102300 : ~(_GEN_102637 & _GEN_1767) & _GEN_102300) : _GEN_102300;
  wire        _GEN_102535 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1768 & _GEN_102301 : _GEN_1029 ? ~_GEN_1768 & _GEN_102301 : ~(_GEN_102637 & _GEN_1768) & _GEN_102301) : _GEN_102301;
  wire        _GEN_102536 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1769 & _GEN_102302 : _GEN_1029 ? ~_GEN_1769 & _GEN_102302 : ~(_GEN_102637 & _GEN_1769) & _GEN_102302) : _GEN_102302;
  wire        _GEN_102537 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1770 & _GEN_102303 : _GEN_1029 ? ~_GEN_1770 & _GEN_102303 : ~(_GEN_102637 & _GEN_1770) & _GEN_102303) : _GEN_102303;
  wire        _GEN_102538 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1771 & _GEN_102304 : _GEN_1029 ? ~_GEN_1771 & _GEN_102304 : ~(_GEN_102637 & _GEN_1771) & _GEN_102304) : _GEN_102304;
  wire        _GEN_102539 = _GEN_1027 ? (_GEN_102472 ? ~_GEN_1772 & _GEN_102305 : _GEN_1029 ? ~_GEN_1772 & _GEN_102305 : ~(_GEN_102637 & _GEN_1772) & _GEN_102305) : _GEN_102305;
  wire        _GEN_102540 = _GEN_1027 ? (_GEN_102472 ? ~(&lcam_ldq_idx_0) & _GEN_102306 : _GEN_1029 ? ~(&lcam_ldq_idx_0) & _GEN_102306 : ~(_GEN_102637 & (&lcam_ldq_idx_0)) & _GEN_102306) : _GEN_102306;
  wire        _GEN_102743 = _GEN_1030 ? (_GEN_102706 ? (|lcam_ldq_idx_1) & _GEN_102509 : _GEN_1032 ? (|lcam_ldq_idx_1) & _GEN_102509 : ~(_GEN_102637 & ~(|lcam_ldq_idx_1)) & _GEN_102509) : _GEN_102509;
  wire        _GEN_102744 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1773 & _GEN_102510 : _GEN_1032 ? ~_GEN_1773 & _GEN_102510 : ~(_GEN_102637 & _GEN_1773) & _GEN_102510) : _GEN_102510;
  wire        _GEN_102745 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1774 & _GEN_102511 : _GEN_1032 ? ~_GEN_1774 & _GEN_102511 : ~(_GEN_102637 & _GEN_1774) & _GEN_102511) : _GEN_102511;
  wire        _GEN_102746 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1775 & _GEN_102512 : _GEN_1032 ? ~_GEN_1775 & _GEN_102512 : ~(_GEN_102637 & _GEN_1775) & _GEN_102512) : _GEN_102512;
  wire        _GEN_102747 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1776 & _GEN_102513 : _GEN_1032 ? ~_GEN_1776 & _GEN_102513 : ~(_GEN_102637 & _GEN_1776) & _GEN_102513) : _GEN_102513;
  wire        _GEN_102748 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1777 & _GEN_102514 : _GEN_1032 ? ~_GEN_1777 & _GEN_102514 : ~(_GEN_102637 & _GEN_1777) & _GEN_102514) : _GEN_102514;
  wire        _GEN_102749 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1778 & _GEN_102515 : _GEN_1032 ? ~_GEN_1778 & _GEN_102515 : ~(_GEN_102637 & _GEN_1778) & _GEN_102515) : _GEN_102515;
  wire        _GEN_102750 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1779 & _GEN_102516 : _GEN_1032 ? ~_GEN_1779 & _GEN_102516 : ~(_GEN_102637 & _GEN_1779) & _GEN_102516) : _GEN_102516;
  wire        _GEN_102751 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1780 & _GEN_102517 : _GEN_1032 ? ~_GEN_1780 & _GEN_102517 : ~(_GEN_102637 & _GEN_1780) & _GEN_102517) : _GEN_102517;
  wire        _GEN_102752 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1781 & _GEN_102518 : _GEN_1032 ? ~_GEN_1781 & _GEN_102518 : ~(_GEN_102637 & _GEN_1781) & _GEN_102518) : _GEN_102518;
  wire        _GEN_102753 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1782 & _GEN_102519 : _GEN_1032 ? ~_GEN_1782 & _GEN_102519 : ~(_GEN_102637 & _GEN_1782) & _GEN_102519) : _GEN_102519;
  wire        _GEN_102754 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1783 & _GEN_102520 : _GEN_1032 ? ~_GEN_1783 & _GEN_102520 : ~(_GEN_102637 & _GEN_1783) & _GEN_102520) : _GEN_102520;
  wire        _GEN_102755 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1784 & _GEN_102521 : _GEN_1032 ? ~_GEN_1784 & _GEN_102521 : ~(_GEN_102637 & _GEN_1784) & _GEN_102521) : _GEN_102521;
  wire        _GEN_102756 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1785 & _GEN_102522 : _GEN_1032 ? ~_GEN_1785 & _GEN_102522 : ~(_GEN_102637 & _GEN_1785) & _GEN_102522) : _GEN_102522;
  wire        _GEN_102757 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1786 & _GEN_102523 : _GEN_1032 ? ~_GEN_1786 & _GEN_102523 : ~(_GEN_102637 & _GEN_1786) & _GEN_102523) : _GEN_102523;
  wire        _GEN_102758 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1787 & _GEN_102524 : _GEN_1032 ? ~_GEN_1787 & _GEN_102524 : ~(_GEN_102637 & _GEN_1787) & _GEN_102524) : _GEN_102524;
  wire        _GEN_102759 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1788 & _GEN_102525 : _GEN_1032 ? ~_GEN_1788 & _GEN_102525 : ~(_GEN_102637 & _GEN_1788) & _GEN_102525) : _GEN_102525;
  wire        _GEN_102760 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1789 & _GEN_102526 : _GEN_1032 ? ~_GEN_1789 & _GEN_102526 : ~(_GEN_102637 & _GEN_1789) & _GEN_102526) : _GEN_102526;
  wire        _GEN_102761 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1790 & _GEN_102527 : _GEN_1032 ? ~_GEN_1790 & _GEN_102527 : ~(_GEN_102637 & _GEN_1790) & _GEN_102527) : _GEN_102527;
  wire        _GEN_102762 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1791 & _GEN_102528 : _GEN_1032 ? ~_GEN_1791 & _GEN_102528 : ~(_GEN_102637 & _GEN_1791) & _GEN_102528) : _GEN_102528;
  wire        _GEN_102763 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1792 & _GEN_102529 : _GEN_1032 ? ~_GEN_1792 & _GEN_102529 : ~(_GEN_102637 & _GEN_1792) & _GEN_102529) : _GEN_102529;
  wire        _GEN_102764 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1793 & _GEN_102530 : _GEN_1032 ? ~_GEN_1793 & _GEN_102530 : ~(_GEN_102637 & _GEN_1793) & _GEN_102530) : _GEN_102530;
  wire        _GEN_102765 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1794 & _GEN_102531 : _GEN_1032 ? ~_GEN_1794 & _GEN_102531 : ~(_GEN_102637 & _GEN_1794) & _GEN_102531) : _GEN_102531;
  wire        _GEN_102766 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1795 & _GEN_102532 : _GEN_1032 ? ~_GEN_1795 & _GEN_102532 : ~(_GEN_102637 & _GEN_1795) & _GEN_102532) : _GEN_102532;
  wire        _GEN_102767 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1796 & _GEN_102533 : _GEN_1032 ? ~_GEN_1796 & _GEN_102533 : ~(_GEN_102637 & _GEN_1796) & _GEN_102533) : _GEN_102533;
  wire        _GEN_102768 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1797 & _GEN_102534 : _GEN_1032 ? ~_GEN_1797 & _GEN_102534 : ~(_GEN_102637 & _GEN_1797) & _GEN_102534) : _GEN_102534;
  wire        _GEN_102769 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1798 & _GEN_102535 : _GEN_1032 ? ~_GEN_1798 & _GEN_102535 : ~(_GEN_102637 & _GEN_1798) & _GEN_102535) : _GEN_102535;
  wire        _GEN_102770 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1799 & _GEN_102536 : _GEN_1032 ? ~_GEN_1799 & _GEN_102536 : ~(_GEN_102637 & _GEN_1799) & _GEN_102536) : _GEN_102536;
  wire        _GEN_102771 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1800 & _GEN_102537 : _GEN_1032 ? ~_GEN_1800 & _GEN_102537 : ~(_GEN_102637 & _GEN_1800) & _GEN_102537) : _GEN_102537;
  wire        _GEN_102772 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1801 & _GEN_102538 : _GEN_1032 ? ~_GEN_1801 & _GEN_102538 : ~(_GEN_102637 & _GEN_1801) & _GEN_102538) : _GEN_102538;
  wire        _GEN_102773 = _GEN_1030 ? (_GEN_102706 ? ~_GEN_1802 & _GEN_102539 : _GEN_1032 ? ~_GEN_1802 & _GEN_102539 : ~(_GEN_102637 & _GEN_1802) & _GEN_102539) : _GEN_102539;
  wire        _GEN_102774 = _GEN_1030 ? (_GEN_102706 ? ~(&lcam_ldq_idx_1) & _GEN_102540 : _GEN_1032 ? ~(&lcam_ldq_idx_1) & _GEN_102540 : ~(_GEN_102637 & (&lcam_ldq_idx_1)) & _GEN_102540) : _GEN_102540;
  wire        _GEN_102977 = _GEN_1033 ? (_GEN_102940 ? (|lcam_ldq_idx_0) & _GEN_102743 : _GEN_1035 ? (|lcam_ldq_idx_0) & _GEN_102743 : ~(_GEN_103105 & ~(|lcam_ldq_idx_0)) & _GEN_102743) : _GEN_102743;
  wire        _GEN_102978 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1743 & _GEN_102744 : _GEN_1035 ? ~_GEN_1743 & _GEN_102744 : ~(_GEN_103105 & _GEN_1743) & _GEN_102744) : _GEN_102744;
  wire        _GEN_102979 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1744 & _GEN_102745 : _GEN_1035 ? ~_GEN_1744 & _GEN_102745 : ~(_GEN_103105 & _GEN_1744) & _GEN_102745) : _GEN_102745;
  wire        _GEN_102980 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1745 & _GEN_102746 : _GEN_1035 ? ~_GEN_1745 & _GEN_102746 : ~(_GEN_103105 & _GEN_1745) & _GEN_102746) : _GEN_102746;
  wire        _GEN_102981 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1746 & _GEN_102747 : _GEN_1035 ? ~_GEN_1746 & _GEN_102747 : ~(_GEN_103105 & _GEN_1746) & _GEN_102747) : _GEN_102747;
  wire        _GEN_102982 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1747 & _GEN_102748 : _GEN_1035 ? ~_GEN_1747 & _GEN_102748 : ~(_GEN_103105 & _GEN_1747) & _GEN_102748) : _GEN_102748;
  wire        _GEN_102983 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1748 & _GEN_102749 : _GEN_1035 ? ~_GEN_1748 & _GEN_102749 : ~(_GEN_103105 & _GEN_1748) & _GEN_102749) : _GEN_102749;
  wire        _GEN_102984 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1749 & _GEN_102750 : _GEN_1035 ? ~_GEN_1749 & _GEN_102750 : ~(_GEN_103105 & _GEN_1749) & _GEN_102750) : _GEN_102750;
  wire        _GEN_102985 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1750 & _GEN_102751 : _GEN_1035 ? ~_GEN_1750 & _GEN_102751 : ~(_GEN_103105 & _GEN_1750) & _GEN_102751) : _GEN_102751;
  wire        _GEN_102986 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1751 & _GEN_102752 : _GEN_1035 ? ~_GEN_1751 & _GEN_102752 : ~(_GEN_103105 & _GEN_1751) & _GEN_102752) : _GEN_102752;
  wire        _GEN_102987 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1752 & _GEN_102753 : _GEN_1035 ? ~_GEN_1752 & _GEN_102753 : ~(_GEN_103105 & _GEN_1752) & _GEN_102753) : _GEN_102753;
  wire        _GEN_102988 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1753 & _GEN_102754 : _GEN_1035 ? ~_GEN_1753 & _GEN_102754 : ~(_GEN_103105 & _GEN_1753) & _GEN_102754) : _GEN_102754;
  wire        _GEN_102989 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1754 & _GEN_102755 : _GEN_1035 ? ~_GEN_1754 & _GEN_102755 : ~(_GEN_103105 & _GEN_1754) & _GEN_102755) : _GEN_102755;
  wire        _GEN_102990 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1755 & _GEN_102756 : _GEN_1035 ? ~_GEN_1755 & _GEN_102756 : ~(_GEN_103105 & _GEN_1755) & _GEN_102756) : _GEN_102756;
  wire        _GEN_102991 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1756 & _GEN_102757 : _GEN_1035 ? ~_GEN_1756 & _GEN_102757 : ~(_GEN_103105 & _GEN_1756) & _GEN_102757) : _GEN_102757;
  wire        _GEN_102992 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1757 & _GEN_102758 : _GEN_1035 ? ~_GEN_1757 & _GEN_102758 : ~(_GEN_103105 & _GEN_1757) & _GEN_102758) : _GEN_102758;
  wire        _GEN_102993 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1758 & _GEN_102759 : _GEN_1035 ? ~_GEN_1758 & _GEN_102759 : ~(_GEN_103105 & _GEN_1758) & _GEN_102759) : _GEN_102759;
  wire        _GEN_102994 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1759 & _GEN_102760 : _GEN_1035 ? ~_GEN_1759 & _GEN_102760 : ~(_GEN_103105 & _GEN_1759) & _GEN_102760) : _GEN_102760;
  wire        _GEN_102995 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1760 & _GEN_102761 : _GEN_1035 ? ~_GEN_1760 & _GEN_102761 : ~(_GEN_103105 & _GEN_1760) & _GEN_102761) : _GEN_102761;
  wire        _GEN_102996 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1761 & _GEN_102762 : _GEN_1035 ? ~_GEN_1761 & _GEN_102762 : ~(_GEN_103105 & _GEN_1761) & _GEN_102762) : _GEN_102762;
  wire        _GEN_102997 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1762 & _GEN_102763 : _GEN_1035 ? ~_GEN_1762 & _GEN_102763 : ~(_GEN_103105 & _GEN_1762) & _GEN_102763) : _GEN_102763;
  wire        _GEN_102998 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1763 & _GEN_102764 : _GEN_1035 ? ~_GEN_1763 & _GEN_102764 : ~(_GEN_103105 & _GEN_1763) & _GEN_102764) : _GEN_102764;
  wire        _GEN_102999 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1764 & _GEN_102765 : _GEN_1035 ? ~_GEN_1764 & _GEN_102765 : ~(_GEN_103105 & _GEN_1764) & _GEN_102765) : _GEN_102765;
  wire        _GEN_103000 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1765 & _GEN_102766 : _GEN_1035 ? ~_GEN_1765 & _GEN_102766 : ~(_GEN_103105 & _GEN_1765) & _GEN_102766) : _GEN_102766;
  wire        _GEN_103001 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1766 & _GEN_102767 : _GEN_1035 ? ~_GEN_1766 & _GEN_102767 : ~(_GEN_103105 & _GEN_1766) & _GEN_102767) : _GEN_102767;
  wire        _GEN_103002 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1767 & _GEN_102768 : _GEN_1035 ? ~_GEN_1767 & _GEN_102768 : ~(_GEN_103105 & _GEN_1767) & _GEN_102768) : _GEN_102768;
  wire        _GEN_103003 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1768 & _GEN_102769 : _GEN_1035 ? ~_GEN_1768 & _GEN_102769 : ~(_GEN_103105 & _GEN_1768) & _GEN_102769) : _GEN_102769;
  wire        _GEN_103004 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1769 & _GEN_102770 : _GEN_1035 ? ~_GEN_1769 & _GEN_102770 : ~(_GEN_103105 & _GEN_1769) & _GEN_102770) : _GEN_102770;
  wire        _GEN_103005 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1770 & _GEN_102771 : _GEN_1035 ? ~_GEN_1770 & _GEN_102771 : ~(_GEN_103105 & _GEN_1770) & _GEN_102771) : _GEN_102771;
  wire        _GEN_103006 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1771 & _GEN_102772 : _GEN_1035 ? ~_GEN_1771 & _GEN_102772 : ~(_GEN_103105 & _GEN_1771) & _GEN_102772) : _GEN_102772;
  wire        _GEN_103007 = _GEN_1033 ? (_GEN_102940 ? ~_GEN_1772 & _GEN_102773 : _GEN_1035 ? ~_GEN_1772 & _GEN_102773 : ~(_GEN_103105 & _GEN_1772) & _GEN_102773) : _GEN_102773;
  wire        _GEN_103008 = _GEN_1033 ? (_GEN_102940 ? ~(&lcam_ldq_idx_0) & _GEN_102774 : _GEN_1035 ? ~(&lcam_ldq_idx_0) & _GEN_102774 : ~(_GEN_103105 & (&lcam_ldq_idx_0)) & _GEN_102774) : _GEN_102774;
  wire        _GEN_103211 = _GEN_1036 ? (_GEN_103174 ? (|lcam_ldq_idx_1) & _GEN_102977 : _GEN_1038 ? (|lcam_ldq_idx_1) & _GEN_102977 : ~(_GEN_103105 & ~(|lcam_ldq_idx_1)) & _GEN_102977) : _GEN_102977;
  wire        _GEN_103212 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1773 & _GEN_102978 : _GEN_1038 ? ~_GEN_1773 & _GEN_102978 : ~(_GEN_103105 & _GEN_1773) & _GEN_102978) : _GEN_102978;
  wire        _GEN_103213 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1774 & _GEN_102979 : _GEN_1038 ? ~_GEN_1774 & _GEN_102979 : ~(_GEN_103105 & _GEN_1774) & _GEN_102979) : _GEN_102979;
  wire        _GEN_103214 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1775 & _GEN_102980 : _GEN_1038 ? ~_GEN_1775 & _GEN_102980 : ~(_GEN_103105 & _GEN_1775) & _GEN_102980) : _GEN_102980;
  wire        _GEN_103215 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1776 & _GEN_102981 : _GEN_1038 ? ~_GEN_1776 & _GEN_102981 : ~(_GEN_103105 & _GEN_1776) & _GEN_102981) : _GEN_102981;
  wire        _GEN_103216 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1777 & _GEN_102982 : _GEN_1038 ? ~_GEN_1777 & _GEN_102982 : ~(_GEN_103105 & _GEN_1777) & _GEN_102982) : _GEN_102982;
  wire        _GEN_103217 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1778 & _GEN_102983 : _GEN_1038 ? ~_GEN_1778 & _GEN_102983 : ~(_GEN_103105 & _GEN_1778) & _GEN_102983) : _GEN_102983;
  wire        _GEN_103218 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1779 & _GEN_102984 : _GEN_1038 ? ~_GEN_1779 & _GEN_102984 : ~(_GEN_103105 & _GEN_1779) & _GEN_102984) : _GEN_102984;
  wire        _GEN_103219 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1780 & _GEN_102985 : _GEN_1038 ? ~_GEN_1780 & _GEN_102985 : ~(_GEN_103105 & _GEN_1780) & _GEN_102985) : _GEN_102985;
  wire        _GEN_103220 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1781 & _GEN_102986 : _GEN_1038 ? ~_GEN_1781 & _GEN_102986 : ~(_GEN_103105 & _GEN_1781) & _GEN_102986) : _GEN_102986;
  wire        _GEN_103221 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1782 & _GEN_102987 : _GEN_1038 ? ~_GEN_1782 & _GEN_102987 : ~(_GEN_103105 & _GEN_1782) & _GEN_102987) : _GEN_102987;
  wire        _GEN_103222 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1783 & _GEN_102988 : _GEN_1038 ? ~_GEN_1783 & _GEN_102988 : ~(_GEN_103105 & _GEN_1783) & _GEN_102988) : _GEN_102988;
  wire        _GEN_103223 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1784 & _GEN_102989 : _GEN_1038 ? ~_GEN_1784 & _GEN_102989 : ~(_GEN_103105 & _GEN_1784) & _GEN_102989) : _GEN_102989;
  wire        _GEN_103224 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1785 & _GEN_102990 : _GEN_1038 ? ~_GEN_1785 & _GEN_102990 : ~(_GEN_103105 & _GEN_1785) & _GEN_102990) : _GEN_102990;
  wire        _GEN_103225 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1786 & _GEN_102991 : _GEN_1038 ? ~_GEN_1786 & _GEN_102991 : ~(_GEN_103105 & _GEN_1786) & _GEN_102991) : _GEN_102991;
  wire        _GEN_103226 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1787 & _GEN_102992 : _GEN_1038 ? ~_GEN_1787 & _GEN_102992 : ~(_GEN_103105 & _GEN_1787) & _GEN_102992) : _GEN_102992;
  wire        _GEN_103227 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1788 & _GEN_102993 : _GEN_1038 ? ~_GEN_1788 & _GEN_102993 : ~(_GEN_103105 & _GEN_1788) & _GEN_102993) : _GEN_102993;
  wire        _GEN_103228 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1789 & _GEN_102994 : _GEN_1038 ? ~_GEN_1789 & _GEN_102994 : ~(_GEN_103105 & _GEN_1789) & _GEN_102994) : _GEN_102994;
  wire        _GEN_103229 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1790 & _GEN_102995 : _GEN_1038 ? ~_GEN_1790 & _GEN_102995 : ~(_GEN_103105 & _GEN_1790) & _GEN_102995) : _GEN_102995;
  wire        _GEN_103230 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1791 & _GEN_102996 : _GEN_1038 ? ~_GEN_1791 & _GEN_102996 : ~(_GEN_103105 & _GEN_1791) & _GEN_102996) : _GEN_102996;
  wire        _GEN_103231 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1792 & _GEN_102997 : _GEN_1038 ? ~_GEN_1792 & _GEN_102997 : ~(_GEN_103105 & _GEN_1792) & _GEN_102997) : _GEN_102997;
  wire        _GEN_103232 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1793 & _GEN_102998 : _GEN_1038 ? ~_GEN_1793 & _GEN_102998 : ~(_GEN_103105 & _GEN_1793) & _GEN_102998) : _GEN_102998;
  wire        _GEN_103233 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1794 & _GEN_102999 : _GEN_1038 ? ~_GEN_1794 & _GEN_102999 : ~(_GEN_103105 & _GEN_1794) & _GEN_102999) : _GEN_102999;
  wire        _GEN_103234 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1795 & _GEN_103000 : _GEN_1038 ? ~_GEN_1795 & _GEN_103000 : ~(_GEN_103105 & _GEN_1795) & _GEN_103000) : _GEN_103000;
  wire        _GEN_103235 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1796 & _GEN_103001 : _GEN_1038 ? ~_GEN_1796 & _GEN_103001 : ~(_GEN_103105 & _GEN_1796) & _GEN_103001) : _GEN_103001;
  wire        _GEN_103236 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1797 & _GEN_103002 : _GEN_1038 ? ~_GEN_1797 & _GEN_103002 : ~(_GEN_103105 & _GEN_1797) & _GEN_103002) : _GEN_103002;
  wire        _GEN_103237 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1798 & _GEN_103003 : _GEN_1038 ? ~_GEN_1798 & _GEN_103003 : ~(_GEN_103105 & _GEN_1798) & _GEN_103003) : _GEN_103003;
  wire        _GEN_103238 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1799 & _GEN_103004 : _GEN_1038 ? ~_GEN_1799 & _GEN_103004 : ~(_GEN_103105 & _GEN_1799) & _GEN_103004) : _GEN_103004;
  wire        _GEN_103239 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1800 & _GEN_103005 : _GEN_1038 ? ~_GEN_1800 & _GEN_103005 : ~(_GEN_103105 & _GEN_1800) & _GEN_103005) : _GEN_103005;
  wire        _GEN_103240 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1801 & _GEN_103006 : _GEN_1038 ? ~_GEN_1801 & _GEN_103006 : ~(_GEN_103105 & _GEN_1801) & _GEN_103006) : _GEN_103006;
  wire        _GEN_103241 = _GEN_1036 ? (_GEN_103174 ? ~_GEN_1802 & _GEN_103007 : _GEN_1038 ? ~_GEN_1802 & _GEN_103007 : ~(_GEN_103105 & _GEN_1802) & _GEN_103007) : _GEN_103007;
  wire        _GEN_103242 = _GEN_1036 ? (_GEN_103174 ? ~(&lcam_ldq_idx_1) & _GEN_103008 : _GEN_1038 ? ~(&lcam_ldq_idx_1) & _GEN_103008 : ~(_GEN_103105 & (&lcam_ldq_idx_1)) & _GEN_103008) : _GEN_103008;
  wire        _GEN_103445 = _GEN_1039 ? (_GEN_103408 ? (|lcam_ldq_idx_0) & _GEN_103211 : _GEN_1041 ? (|lcam_ldq_idx_0) & _GEN_103211 : ~(_GEN_103573 & ~(|lcam_ldq_idx_0)) & _GEN_103211) : _GEN_103211;
  wire        _GEN_103446 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1743 & _GEN_103212 : _GEN_1041 ? ~_GEN_1743 & _GEN_103212 : ~(_GEN_103573 & _GEN_1743) & _GEN_103212) : _GEN_103212;
  wire        _GEN_103447 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1744 & _GEN_103213 : _GEN_1041 ? ~_GEN_1744 & _GEN_103213 : ~(_GEN_103573 & _GEN_1744) & _GEN_103213) : _GEN_103213;
  wire        _GEN_103448 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1745 & _GEN_103214 : _GEN_1041 ? ~_GEN_1745 & _GEN_103214 : ~(_GEN_103573 & _GEN_1745) & _GEN_103214) : _GEN_103214;
  wire        _GEN_103449 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1746 & _GEN_103215 : _GEN_1041 ? ~_GEN_1746 & _GEN_103215 : ~(_GEN_103573 & _GEN_1746) & _GEN_103215) : _GEN_103215;
  wire        _GEN_103450 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1747 & _GEN_103216 : _GEN_1041 ? ~_GEN_1747 & _GEN_103216 : ~(_GEN_103573 & _GEN_1747) & _GEN_103216) : _GEN_103216;
  wire        _GEN_103451 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1748 & _GEN_103217 : _GEN_1041 ? ~_GEN_1748 & _GEN_103217 : ~(_GEN_103573 & _GEN_1748) & _GEN_103217) : _GEN_103217;
  wire        _GEN_103452 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1749 & _GEN_103218 : _GEN_1041 ? ~_GEN_1749 & _GEN_103218 : ~(_GEN_103573 & _GEN_1749) & _GEN_103218) : _GEN_103218;
  wire        _GEN_103453 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1750 & _GEN_103219 : _GEN_1041 ? ~_GEN_1750 & _GEN_103219 : ~(_GEN_103573 & _GEN_1750) & _GEN_103219) : _GEN_103219;
  wire        _GEN_103454 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1751 & _GEN_103220 : _GEN_1041 ? ~_GEN_1751 & _GEN_103220 : ~(_GEN_103573 & _GEN_1751) & _GEN_103220) : _GEN_103220;
  wire        _GEN_103455 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1752 & _GEN_103221 : _GEN_1041 ? ~_GEN_1752 & _GEN_103221 : ~(_GEN_103573 & _GEN_1752) & _GEN_103221) : _GEN_103221;
  wire        _GEN_103456 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1753 & _GEN_103222 : _GEN_1041 ? ~_GEN_1753 & _GEN_103222 : ~(_GEN_103573 & _GEN_1753) & _GEN_103222) : _GEN_103222;
  wire        _GEN_103457 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1754 & _GEN_103223 : _GEN_1041 ? ~_GEN_1754 & _GEN_103223 : ~(_GEN_103573 & _GEN_1754) & _GEN_103223) : _GEN_103223;
  wire        _GEN_103458 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1755 & _GEN_103224 : _GEN_1041 ? ~_GEN_1755 & _GEN_103224 : ~(_GEN_103573 & _GEN_1755) & _GEN_103224) : _GEN_103224;
  wire        _GEN_103459 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1756 & _GEN_103225 : _GEN_1041 ? ~_GEN_1756 & _GEN_103225 : ~(_GEN_103573 & _GEN_1756) & _GEN_103225) : _GEN_103225;
  wire        _GEN_103460 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1757 & _GEN_103226 : _GEN_1041 ? ~_GEN_1757 & _GEN_103226 : ~(_GEN_103573 & _GEN_1757) & _GEN_103226) : _GEN_103226;
  wire        _GEN_103461 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1758 & _GEN_103227 : _GEN_1041 ? ~_GEN_1758 & _GEN_103227 : ~(_GEN_103573 & _GEN_1758) & _GEN_103227) : _GEN_103227;
  wire        _GEN_103462 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1759 & _GEN_103228 : _GEN_1041 ? ~_GEN_1759 & _GEN_103228 : ~(_GEN_103573 & _GEN_1759) & _GEN_103228) : _GEN_103228;
  wire        _GEN_103463 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1760 & _GEN_103229 : _GEN_1041 ? ~_GEN_1760 & _GEN_103229 : ~(_GEN_103573 & _GEN_1760) & _GEN_103229) : _GEN_103229;
  wire        _GEN_103464 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1761 & _GEN_103230 : _GEN_1041 ? ~_GEN_1761 & _GEN_103230 : ~(_GEN_103573 & _GEN_1761) & _GEN_103230) : _GEN_103230;
  wire        _GEN_103465 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1762 & _GEN_103231 : _GEN_1041 ? ~_GEN_1762 & _GEN_103231 : ~(_GEN_103573 & _GEN_1762) & _GEN_103231) : _GEN_103231;
  wire        _GEN_103466 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1763 & _GEN_103232 : _GEN_1041 ? ~_GEN_1763 & _GEN_103232 : ~(_GEN_103573 & _GEN_1763) & _GEN_103232) : _GEN_103232;
  wire        _GEN_103467 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1764 & _GEN_103233 : _GEN_1041 ? ~_GEN_1764 & _GEN_103233 : ~(_GEN_103573 & _GEN_1764) & _GEN_103233) : _GEN_103233;
  wire        _GEN_103468 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1765 & _GEN_103234 : _GEN_1041 ? ~_GEN_1765 & _GEN_103234 : ~(_GEN_103573 & _GEN_1765) & _GEN_103234) : _GEN_103234;
  wire        _GEN_103469 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1766 & _GEN_103235 : _GEN_1041 ? ~_GEN_1766 & _GEN_103235 : ~(_GEN_103573 & _GEN_1766) & _GEN_103235) : _GEN_103235;
  wire        _GEN_103470 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1767 & _GEN_103236 : _GEN_1041 ? ~_GEN_1767 & _GEN_103236 : ~(_GEN_103573 & _GEN_1767) & _GEN_103236) : _GEN_103236;
  wire        _GEN_103471 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1768 & _GEN_103237 : _GEN_1041 ? ~_GEN_1768 & _GEN_103237 : ~(_GEN_103573 & _GEN_1768) & _GEN_103237) : _GEN_103237;
  wire        _GEN_103472 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1769 & _GEN_103238 : _GEN_1041 ? ~_GEN_1769 & _GEN_103238 : ~(_GEN_103573 & _GEN_1769) & _GEN_103238) : _GEN_103238;
  wire        _GEN_103473 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1770 & _GEN_103239 : _GEN_1041 ? ~_GEN_1770 & _GEN_103239 : ~(_GEN_103573 & _GEN_1770) & _GEN_103239) : _GEN_103239;
  wire        _GEN_103474 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1771 & _GEN_103240 : _GEN_1041 ? ~_GEN_1771 & _GEN_103240 : ~(_GEN_103573 & _GEN_1771) & _GEN_103240) : _GEN_103240;
  wire        _GEN_103475 = _GEN_1039 ? (_GEN_103408 ? ~_GEN_1772 & _GEN_103241 : _GEN_1041 ? ~_GEN_1772 & _GEN_103241 : ~(_GEN_103573 & _GEN_1772) & _GEN_103241) : _GEN_103241;
  wire        _GEN_103476 = _GEN_1039 ? (_GEN_103408 ? ~(&lcam_ldq_idx_0) & _GEN_103242 : _GEN_1041 ? ~(&lcam_ldq_idx_0) & _GEN_103242 : ~(_GEN_103573 & (&lcam_ldq_idx_0)) & _GEN_103242) : _GEN_103242;
  wire        _GEN_103679 = _GEN_1042 ? (_GEN_103642 ? (|lcam_ldq_idx_1) & _GEN_103445 : _GEN_1044 ? (|lcam_ldq_idx_1) & _GEN_103445 : ~(_GEN_103573 & ~(|lcam_ldq_idx_1)) & _GEN_103445) : _GEN_103445;
  wire        _GEN_103680 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1773 & _GEN_103446 : _GEN_1044 ? ~_GEN_1773 & _GEN_103446 : ~(_GEN_103573 & _GEN_1773) & _GEN_103446) : _GEN_103446;
  wire        _GEN_103681 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1774 & _GEN_103447 : _GEN_1044 ? ~_GEN_1774 & _GEN_103447 : ~(_GEN_103573 & _GEN_1774) & _GEN_103447) : _GEN_103447;
  wire        _GEN_103682 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1775 & _GEN_103448 : _GEN_1044 ? ~_GEN_1775 & _GEN_103448 : ~(_GEN_103573 & _GEN_1775) & _GEN_103448) : _GEN_103448;
  wire        _GEN_103683 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1776 & _GEN_103449 : _GEN_1044 ? ~_GEN_1776 & _GEN_103449 : ~(_GEN_103573 & _GEN_1776) & _GEN_103449) : _GEN_103449;
  wire        _GEN_103684 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1777 & _GEN_103450 : _GEN_1044 ? ~_GEN_1777 & _GEN_103450 : ~(_GEN_103573 & _GEN_1777) & _GEN_103450) : _GEN_103450;
  wire        _GEN_103685 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1778 & _GEN_103451 : _GEN_1044 ? ~_GEN_1778 & _GEN_103451 : ~(_GEN_103573 & _GEN_1778) & _GEN_103451) : _GEN_103451;
  wire        _GEN_103686 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1779 & _GEN_103452 : _GEN_1044 ? ~_GEN_1779 & _GEN_103452 : ~(_GEN_103573 & _GEN_1779) & _GEN_103452) : _GEN_103452;
  wire        _GEN_103687 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1780 & _GEN_103453 : _GEN_1044 ? ~_GEN_1780 & _GEN_103453 : ~(_GEN_103573 & _GEN_1780) & _GEN_103453) : _GEN_103453;
  wire        _GEN_103688 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1781 & _GEN_103454 : _GEN_1044 ? ~_GEN_1781 & _GEN_103454 : ~(_GEN_103573 & _GEN_1781) & _GEN_103454) : _GEN_103454;
  wire        _GEN_103689 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1782 & _GEN_103455 : _GEN_1044 ? ~_GEN_1782 & _GEN_103455 : ~(_GEN_103573 & _GEN_1782) & _GEN_103455) : _GEN_103455;
  wire        _GEN_103690 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1783 & _GEN_103456 : _GEN_1044 ? ~_GEN_1783 & _GEN_103456 : ~(_GEN_103573 & _GEN_1783) & _GEN_103456) : _GEN_103456;
  wire        _GEN_103691 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1784 & _GEN_103457 : _GEN_1044 ? ~_GEN_1784 & _GEN_103457 : ~(_GEN_103573 & _GEN_1784) & _GEN_103457) : _GEN_103457;
  wire        _GEN_103692 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1785 & _GEN_103458 : _GEN_1044 ? ~_GEN_1785 & _GEN_103458 : ~(_GEN_103573 & _GEN_1785) & _GEN_103458) : _GEN_103458;
  wire        _GEN_103693 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1786 & _GEN_103459 : _GEN_1044 ? ~_GEN_1786 & _GEN_103459 : ~(_GEN_103573 & _GEN_1786) & _GEN_103459) : _GEN_103459;
  wire        _GEN_103694 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1787 & _GEN_103460 : _GEN_1044 ? ~_GEN_1787 & _GEN_103460 : ~(_GEN_103573 & _GEN_1787) & _GEN_103460) : _GEN_103460;
  wire        _GEN_103695 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1788 & _GEN_103461 : _GEN_1044 ? ~_GEN_1788 & _GEN_103461 : ~(_GEN_103573 & _GEN_1788) & _GEN_103461) : _GEN_103461;
  wire        _GEN_103696 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1789 & _GEN_103462 : _GEN_1044 ? ~_GEN_1789 & _GEN_103462 : ~(_GEN_103573 & _GEN_1789) & _GEN_103462) : _GEN_103462;
  wire        _GEN_103697 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1790 & _GEN_103463 : _GEN_1044 ? ~_GEN_1790 & _GEN_103463 : ~(_GEN_103573 & _GEN_1790) & _GEN_103463) : _GEN_103463;
  wire        _GEN_103698 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1791 & _GEN_103464 : _GEN_1044 ? ~_GEN_1791 & _GEN_103464 : ~(_GEN_103573 & _GEN_1791) & _GEN_103464) : _GEN_103464;
  wire        _GEN_103699 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1792 & _GEN_103465 : _GEN_1044 ? ~_GEN_1792 & _GEN_103465 : ~(_GEN_103573 & _GEN_1792) & _GEN_103465) : _GEN_103465;
  wire        _GEN_103700 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1793 & _GEN_103466 : _GEN_1044 ? ~_GEN_1793 & _GEN_103466 : ~(_GEN_103573 & _GEN_1793) & _GEN_103466) : _GEN_103466;
  wire        _GEN_103701 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1794 & _GEN_103467 : _GEN_1044 ? ~_GEN_1794 & _GEN_103467 : ~(_GEN_103573 & _GEN_1794) & _GEN_103467) : _GEN_103467;
  wire        _GEN_103702 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1795 & _GEN_103468 : _GEN_1044 ? ~_GEN_1795 & _GEN_103468 : ~(_GEN_103573 & _GEN_1795) & _GEN_103468) : _GEN_103468;
  wire        _GEN_103703 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1796 & _GEN_103469 : _GEN_1044 ? ~_GEN_1796 & _GEN_103469 : ~(_GEN_103573 & _GEN_1796) & _GEN_103469) : _GEN_103469;
  wire        _GEN_103704 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1797 & _GEN_103470 : _GEN_1044 ? ~_GEN_1797 & _GEN_103470 : ~(_GEN_103573 & _GEN_1797) & _GEN_103470) : _GEN_103470;
  wire        _GEN_103705 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1798 & _GEN_103471 : _GEN_1044 ? ~_GEN_1798 & _GEN_103471 : ~(_GEN_103573 & _GEN_1798) & _GEN_103471) : _GEN_103471;
  wire        _GEN_103706 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1799 & _GEN_103472 : _GEN_1044 ? ~_GEN_1799 & _GEN_103472 : ~(_GEN_103573 & _GEN_1799) & _GEN_103472) : _GEN_103472;
  wire        _GEN_103707 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1800 & _GEN_103473 : _GEN_1044 ? ~_GEN_1800 & _GEN_103473 : ~(_GEN_103573 & _GEN_1800) & _GEN_103473) : _GEN_103473;
  wire        _GEN_103708 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1801 & _GEN_103474 : _GEN_1044 ? ~_GEN_1801 & _GEN_103474 : ~(_GEN_103573 & _GEN_1801) & _GEN_103474) : _GEN_103474;
  wire        _GEN_103709 = _GEN_1042 ? (_GEN_103642 ? ~_GEN_1802 & _GEN_103475 : _GEN_1044 ? ~_GEN_1802 & _GEN_103475 : ~(_GEN_103573 & _GEN_1802) & _GEN_103475) : _GEN_103475;
  wire        _GEN_103710 = _GEN_1042 ? (_GEN_103642 ? ~(&lcam_ldq_idx_1) & _GEN_103476 : _GEN_1044 ? ~(&lcam_ldq_idx_1) & _GEN_103476 : ~(_GEN_103573 & (&lcam_ldq_idx_1)) & _GEN_103476) : _GEN_103476;
  wire        _GEN_103913 = _GEN_1045 ? (_GEN_103876 ? (|lcam_ldq_idx_0) & _GEN_103679 : _GEN_1047 ? (|lcam_ldq_idx_0) & _GEN_103679 : ~(_GEN_104041 & ~(|lcam_ldq_idx_0)) & _GEN_103679) : _GEN_103679;
  wire        _GEN_103914 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1743 & _GEN_103680 : _GEN_1047 ? ~_GEN_1743 & _GEN_103680 : ~(_GEN_104041 & _GEN_1743) & _GEN_103680) : _GEN_103680;
  wire        _GEN_103915 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1744 & _GEN_103681 : _GEN_1047 ? ~_GEN_1744 & _GEN_103681 : ~(_GEN_104041 & _GEN_1744) & _GEN_103681) : _GEN_103681;
  wire        _GEN_103916 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1745 & _GEN_103682 : _GEN_1047 ? ~_GEN_1745 & _GEN_103682 : ~(_GEN_104041 & _GEN_1745) & _GEN_103682) : _GEN_103682;
  wire        _GEN_103917 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1746 & _GEN_103683 : _GEN_1047 ? ~_GEN_1746 & _GEN_103683 : ~(_GEN_104041 & _GEN_1746) & _GEN_103683) : _GEN_103683;
  wire        _GEN_103918 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1747 & _GEN_103684 : _GEN_1047 ? ~_GEN_1747 & _GEN_103684 : ~(_GEN_104041 & _GEN_1747) & _GEN_103684) : _GEN_103684;
  wire        _GEN_103919 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1748 & _GEN_103685 : _GEN_1047 ? ~_GEN_1748 & _GEN_103685 : ~(_GEN_104041 & _GEN_1748) & _GEN_103685) : _GEN_103685;
  wire        _GEN_103920 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1749 & _GEN_103686 : _GEN_1047 ? ~_GEN_1749 & _GEN_103686 : ~(_GEN_104041 & _GEN_1749) & _GEN_103686) : _GEN_103686;
  wire        _GEN_103921 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1750 & _GEN_103687 : _GEN_1047 ? ~_GEN_1750 & _GEN_103687 : ~(_GEN_104041 & _GEN_1750) & _GEN_103687) : _GEN_103687;
  wire        _GEN_103922 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1751 & _GEN_103688 : _GEN_1047 ? ~_GEN_1751 & _GEN_103688 : ~(_GEN_104041 & _GEN_1751) & _GEN_103688) : _GEN_103688;
  wire        _GEN_103923 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1752 & _GEN_103689 : _GEN_1047 ? ~_GEN_1752 & _GEN_103689 : ~(_GEN_104041 & _GEN_1752) & _GEN_103689) : _GEN_103689;
  wire        _GEN_103924 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1753 & _GEN_103690 : _GEN_1047 ? ~_GEN_1753 & _GEN_103690 : ~(_GEN_104041 & _GEN_1753) & _GEN_103690) : _GEN_103690;
  wire        _GEN_103925 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1754 & _GEN_103691 : _GEN_1047 ? ~_GEN_1754 & _GEN_103691 : ~(_GEN_104041 & _GEN_1754) & _GEN_103691) : _GEN_103691;
  wire        _GEN_103926 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1755 & _GEN_103692 : _GEN_1047 ? ~_GEN_1755 & _GEN_103692 : ~(_GEN_104041 & _GEN_1755) & _GEN_103692) : _GEN_103692;
  wire        _GEN_103927 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1756 & _GEN_103693 : _GEN_1047 ? ~_GEN_1756 & _GEN_103693 : ~(_GEN_104041 & _GEN_1756) & _GEN_103693) : _GEN_103693;
  wire        _GEN_103928 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1757 & _GEN_103694 : _GEN_1047 ? ~_GEN_1757 & _GEN_103694 : ~(_GEN_104041 & _GEN_1757) & _GEN_103694) : _GEN_103694;
  wire        _GEN_103929 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1758 & _GEN_103695 : _GEN_1047 ? ~_GEN_1758 & _GEN_103695 : ~(_GEN_104041 & _GEN_1758) & _GEN_103695) : _GEN_103695;
  wire        _GEN_103930 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1759 & _GEN_103696 : _GEN_1047 ? ~_GEN_1759 & _GEN_103696 : ~(_GEN_104041 & _GEN_1759) & _GEN_103696) : _GEN_103696;
  wire        _GEN_103931 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1760 & _GEN_103697 : _GEN_1047 ? ~_GEN_1760 & _GEN_103697 : ~(_GEN_104041 & _GEN_1760) & _GEN_103697) : _GEN_103697;
  wire        _GEN_103932 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1761 & _GEN_103698 : _GEN_1047 ? ~_GEN_1761 & _GEN_103698 : ~(_GEN_104041 & _GEN_1761) & _GEN_103698) : _GEN_103698;
  wire        _GEN_103933 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1762 & _GEN_103699 : _GEN_1047 ? ~_GEN_1762 & _GEN_103699 : ~(_GEN_104041 & _GEN_1762) & _GEN_103699) : _GEN_103699;
  wire        _GEN_103934 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1763 & _GEN_103700 : _GEN_1047 ? ~_GEN_1763 & _GEN_103700 : ~(_GEN_104041 & _GEN_1763) & _GEN_103700) : _GEN_103700;
  wire        _GEN_103935 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1764 & _GEN_103701 : _GEN_1047 ? ~_GEN_1764 & _GEN_103701 : ~(_GEN_104041 & _GEN_1764) & _GEN_103701) : _GEN_103701;
  wire        _GEN_103936 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1765 & _GEN_103702 : _GEN_1047 ? ~_GEN_1765 & _GEN_103702 : ~(_GEN_104041 & _GEN_1765) & _GEN_103702) : _GEN_103702;
  wire        _GEN_103937 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1766 & _GEN_103703 : _GEN_1047 ? ~_GEN_1766 & _GEN_103703 : ~(_GEN_104041 & _GEN_1766) & _GEN_103703) : _GEN_103703;
  wire        _GEN_103938 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1767 & _GEN_103704 : _GEN_1047 ? ~_GEN_1767 & _GEN_103704 : ~(_GEN_104041 & _GEN_1767) & _GEN_103704) : _GEN_103704;
  wire        _GEN_103939 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1768 & _GEN_103705 : _GEN_1047 ? ~_GEN_1768 & _GEN_103705 : ~(_GEN_104041 & _GEN_1768) & _GEN_103705) : _GEN_103705;
  wire        _GEN_103940 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1769 & _GEN_103706 : _GEN_1047 ? ~_GEN_1769 & _GEN_103706 : ~(_GEN_104041 & _GEN_1769) & _GEN_103706) : _GEN_103706;
  wire        _GEN_103941 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1770 & _GEN_103707 : _GEN_1047 ? ~_GEN_1770 & _GEN_103707 : ~(_GEN_104041 & _GEN_1770) & _GEN_103707) : _GEN_103707;
  wire        _GEN_103942 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1771 & _GEN_103708 : _GEN_1047 ? ~_GEN_1771 & _GEN_103708 : ~(_GEN_104041 & _GEN_1771) & _GEN_103708) : _GEN_103708;
  wire        _GEN_103943 = _GEN_1045 ? (_GEN_103876 ? ~_GEN_1772 & _GEN_103709 : _GEN_1047 ? ~_GEN_1772 & _GEN_103709 : ~(_GEN_104041 & _GEN_1772) & _GEN_103709) : _GEN_103709;
  wire        _GEN_103944 = _GEN_1045 ? (_GEN_103876 ? ~(&lcam_ldq_idx_0) & _GEN_103710 : _GEN_1047 ? ~(&lcam_ldq_idx_0) & _GEN_103710 : ~(_GEN_104041 & (&lcam_ldq_idx_0)) & _GEN_103710) : _GEN_103710;
  wire        _GEN_104147 = _GEN_1048 ? (_GEN_104110 ? (|lcam_ldq_idx_1) & _GEN_103913 : _GEN_1050 ? (|lcam_ldq_idx_1) & _GEN_103913 : ~(_GEN_104041 & ~(|lcam_ldq_idx_1)) & _GEN_103913) : _GEN_103913;
  wire        _GEN_104148 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1773 & _GEN_103914 : _GEN_1050 ? ~_GEN_1773 & _GEN_103914 : ~(_GEN_104041 & _GEN_1773) & _GEN_103914) : _GEN_103914;
  wire        _GEN_104149 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1774 & _GEN_103915 : _GEN_1050 ? ~_GEN_1774 & _GEN_103915 : ~(_GEN_104041 & _GEN_1774) & _GEN_103915) : _GEN_103915;
  wire        _GEN_104150 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1775 & _GEN_103916 : _GEN_1050 ? ~_GEN_1775 & _GEN_103916 : ~(_GEN_104041 & _GEN_1775) & _GEN_103916) : _GEN_103916;
  wire        _GEN_104151 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1776 & _GEN_103917 : _GEN_1050 ? ~_GEN_1776 & _GEN_103917 : ~(_GEN_104041 & _GEN_1776) & _GEN_103917) : _GEN_103917;
  wire        _GEN_104152 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1777 & _GEN_103918 : _GEN_1050 ? ~_GEN_1777 & _GEN_103918 : ~(_GEN_104041 & _GEN_1777) & _GEN_103918) : _GEN_103918;
  wire        _GEN_104153 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1778 & _GEN_103919 : _GEN_1050 ? ~_GEN_1778 & _GEN_103919 : ~(_GEN_104041 & _GEN_1778) & _GEN_103919) : _GEN_103919;
  wire        _GEN_104154 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1779 & _GEN_103920 : _GEN_1050 ? ~_GEN_1779 & _GEN_103920 : ~(_GEN_104041 & _GEN_1779) & _GEN_103920) : _GEN_103920;
  wire        _GEN_104155 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1780 & _GEN_103921 : _GEN_1050 ? ~_GEN_1780 & _GEN_103921 : ~(_GEN_104041 & _GEN_1780) & _GEN_103921) : _GEN_103921;
  wire        _GEN_104156 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1781 & _GEN_103922 : _GEN_1050 ? ~_GEN_1781 & _GEN_103922 : ~(_GEN_104041 & _GEN_1781) & _GEN_103922) : _GEN_103922;
  wire        _GEN_104157 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1782 & _GEN_103923 : _GEN_1050 ? ~_GEN_1782 & _GEN_103923 : ~(_GEN_104041 & _GEN_1782) & _GEN_103923) : _GEN_103923;
  wire        _GEN_104158 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1783 & _GEN_103924 : _GEN_1050 ? ~_GEN_1783 & _GEN_103924 : ~(_GEN_104041 & _GEN_1783) & _GEN_103924) : _GEN_103924;
  wire        _GEN_104159 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1784 & _GEN_103925 : _GEN_1050 ? ~_GEN_1784 & _GEN_103925 : ~(_GEN_104041 & _GEN_1784) & _GEN_103925) : _GEN_103925;
  wire        _GEN_104160 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1785 & _GEN_103926 : _GEN_1050 ? ~_GEN_1785 & _GEN_103926 : ~(_GEN_104041 & _GEN_1785) & _GEN_103926) : _GEN_103926;
  wire        _GEN_104161 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1786 & _GEN_103927 : _GEN_1050 ? ~_GEN_1786 & _GEN_103927 : ~(_GEN_104041 & _GEN_1786) & _GEN_103927) : _GEN_103927;
  wire        _GEN_104162 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1787 & _GEN_103928 : _GEN_1050 ? ~_GEN_1787 & _GEN_103928 : ~(_GEN_104041 & _GEN_1787) & _GEN_103928) : _GEN_103928;
  wire        _GEN_104163 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1788 & _GEN_103929 : _GEN_1050 ? ~_GEN_1788 & _GEN_103929 : ~(_GEN_104041 & _GEN_1788) & _GEN_103929) : _GEN_103929;
  wire        _GEN_104164 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1789 & _GEN_103930 : _GEN_1050 ? ~_GEN_1789 & _GEN_103930 : ~(_GEN_104041 & _GEN_1789) & _GEN_103930) : _GEN_103930;
  wire        _GEN_104165 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1790 & _GEN_103931 : _GEN_1050 ? ~_GEN_1790 & _GEN_103931 : ~(_GEN_104041 & _GEN_1790) & _GEN_103931) : _GEN_103931;
  wire        _GEN_104166 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1791 & _GEN_103932 : _GEN_1050 ? ~_GEN_1791 & _GEN_103932 : ~(_GEN_104041 & _GEN_1791) & _GEN_103932) : _GEN_103932;
  wire        _GEN_104167 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1792 & _GEN_103933 : _GEN_1050 ? ~_GEN_1792 & _GEN_103933 : ~(_GEN_104041 & _GEN_1792) & _GEN_103933) : _GEN_103933;
  wire        _GEN_104168 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1793 & _GEN_103934 : _GEN_1050 ? ~_GEN_1793 & _GEN_103934 : ~(_GEN_104041 & _GEN_1793) & _GEN_103934) : _GEN_103934;
  wire        _GEN_104169 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1794 & _GEN_103935 : _GEN_1050 ? ~_GEN_1794 & _GEN_103935 : ~(_GEN_104041 & _GEN_1794) & _GEN_103935) : _GEN_103935;
  wire        _GEN_104170 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1795 & _GEN_103936 : _GEN_1050 ? ~_GEN_1795 & _GEN_103936 : ~(_GEN_104041 & _GEN_1795) & _GEN_103936) : _GEN_103936;
  wire        _GEN_104171 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1796 & _GEN_103937 : _GEN_1050 ? ~_GEN_1796 & _GEN_103937 : ~(_GEN_104041 & _GEN_1796) & _GEN_103937) : _GEN_103937;
  wire        _GEN_104172 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1797 & _GEN_103938 : _GEN_1050 ? ~_GEN_1797 & _GEN_103938 : ~(_GEN_104041 & _GEN_1797) & _GEN_103938) : _GEN_103938;
  wire        _GEN_104173 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1798 & _GEN_103939 : _GEN_1050 ? ~_GEN_1798 & _GEN_103939 : ~(_GEN_104041 & _GEN_1798) & _GEN_103939) : _GEN_103939;
  wire        _GEN_104174 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1799 & _GEN_103940 : _GEN_1050 ? ~_GEN_1799 & _GEN_103940 : ~(_GEN_104041 & _GEN_1799) & _GEN_103940) : _GEN_103940;
  wire        _GEN_104175 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1800 & _GEN_103941 : _GEN_1050 ? ~_GEN_1800 & _GEN_103941 : ~(_GEN_104041 & _GEN_1800) & _GEN_103941) : _GEN_103941;
  wire        _GEN_104176 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1801 & _GEN_103942 : _GEN_1050 ? ~_GEN_1801 & _GEN_103942 : ~(_GEN_104041 & _GEN_1801) & _GEN_103942) : _GEN_103942;
  wire        _GEN_104177 = _GEN_1048 ? (_GEN_104110 ? ~_GEN_1802 & _GEN_103943 : _GEN_1050 ? ~_GEN_1802 & _GEN_103943 : ~(_GEN_104041 & _GEN_1802) & _GEN_103943) : _GEN_103943;
  wire        _GEN_104178 = _GEN_1048 ? (_GEN_104110 ? ~(&lcam_ldq_idx_1) & _GEN_103944 : _GEN_1050 ? ~(&lcam_ldq_idx_1) & _GEN_103944 : ~(_GEN_104041 & (&lcam_ldq_idx_1)) & _GEN_103944) : _GEN_103944;
  wire        _GEN_104381 = _GEN_1051 ? (_GEN_104344 ? (|lcam_ldq_idx_0) & _GEN_104147 : _GEN_1053 ? (|lcam_ldq_idx_0) & _GEN_104147 : ~(_GEN_104509 & ~(|lcam_ldq_idx_0)) & _GEN_104147) : _GEN_104147;
  wire        _GEN_104382 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1743 & _GEN_104148 : _GEN_1053 ? ~_GEN_1743 & _GEN_104148 : ~(_GEN_104509 & _GEN_1743) & _GEN_104148) : _GEN_104148;
  wire        _GEN_104383 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1744 & _GEN_104149 : _GEN_1053 ? ~_GEN_1744 & _GEN_104149 : ~(_GEN_104509 & _GEN_1744) & _GEN_104149) : _GEN_104149;
  wire        _GEN_104384 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1745 & _GEN_104150 : _GEN_1053 ? ~_GEN_1745 & _GEN_104150 : ~(_GEN_104509 & _GEN_1745) & _GEN_104150) : _GEN_104150;
  wire        _GEN_104385 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1746 & _GEN_104151 : _GEN_1053 ? ~_GEN_1746 & _GEN_104151 : ~(_GEN_104509 & _GEN_1746) & _GEN_104151) : _GEN_104151;
  wire        _GEN_104386 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1747 & _GEN_104152 : _GEN_1053 ? ~_GEN_1747 & _GEN_104152 : ~(_GEN_104509 & _GEN_1747) & _GEN_104152) : _GEN_104152;
  wire        _GEN_104387 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1748 & _GEN_104153 : _GEN_1053 ? ~_GEN_1748 & _GEN_104153 : ~(_GEN_104509 & _GEN_1748) & _GEN_104153) : _GEN_104153;
  wire        _GEN_104388 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1749 & _GEN_104154 : _GEN_1053 ? ~_GEN_1749 & _GEN_104154 : ~(_GEN_104509 & _GEN_1749) & _GEN_104154) : _GEN_104154;
  wire        _GEN_104389 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1750 & _GEN_104155 : _GEN_1053 ? ~_GEN_1750 & _GEN_104155 : ~(_GEN_104509 & _GEN_1750) & _GEN_104155) : _GEN_104155;
  wire        _GEN_104390 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1751 & _GEN_104156 : _GEN_1053 ? ~_GEN_1751 & _GEN_104156 : ~(_GEN_104509 & _GEN_1751) & _GEN_104156) : _GEN_104156;
  wire        _GEN_104391 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1752 & _GEN_104157 : _GEN_1053 ? ~_GEN_1752 & _GEN_104157 : ~(_GEN_104509 & _GEN_1752) & _GEN_104157) : _GEN_104157;
  wire        _GEN_104392 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1753 & _GEN_104158 : _GEN_1053 ? ~_GEN_1753 & _GEN_104158 : ~(_GEN_104509 & _GEN_1753) & _GEN_104158) : _GEN_104158;
  wire        _GEN_104393 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1754 & _GEN_104159 : _GEN_1053 ? ~_GEN_1754 & _GEN_104159 : ~(_GEN_104509 & _GEN_1754) & _GEN_104159) : _GEN_104159;
  wire        _GEN_104394 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1755 & _GEN_104160 : _GEN_1053 ? ~_GEN_1755 & _GEN_104160 : ~(_GEN_104509 & _GEN_1755) & _GEN_104160) : _GEN_104160;
  wire        _GEN_104395 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1756 & _GEN_104161 : _GEN_1053 ? ~_GEN_1756 & _GEN_104161 : ~(_GEN_104509 & _GEN_1756) & _GEN_104161) : _GEN_104161;
  wire        _GEN_104396 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1757 & _GEN_104162 : _GEN_1053 ? ~_GEN_1757 & _GEN_104162 : ~(_GEN_104509 & _GEN_1757) & _GEN_104162) : _GEN_104162;
  wire        _GEN_104397 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1758 & _GEN_104163 : _GEN_1053 ? ~_GEN_1758 & _GEN_104163 : ~(_GEN_104509 & _GEN_1758) & _GEN_104163) : _GEN_104163;
  wire        _GEN_104398 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1759 & _GEN_104164 : _GEN_1053 ? ~_GEN_1759 & _GEN_104164 : ~(_GEN_104509 & _GEN_1759) & _GEN_104164) : _GEN_104164;
  wire        _GEN_104399 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1760 & _GEN_104165 : _GEN_1053 ? ~_GEN_1760 & _GEN_104165 : ~(_GEN_104509 & _GEN_1760) & _GEN_104165) : _GEN_104165;
  wire        _GEN_104400 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1761 & _GEN_104166 : _GEN_1053 ? ~_GEN_1761 & _GEN_104166 : ~(_GEN_104509 & _GEN_1761) & _GEN_104166) : _GEN_104166;
  wire        _GEN_104401 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1762 & _GEN_104167 : _GEN_1053 ? ~_GEN_1762 & _GEN_104167 : ~(_GEN_104509 & _GEN_1762) & _GEN_104167) : _GEN_104167;
  wire        _GEN_104402 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1763 & _GEN_104168 : _GEN_1053 ? ~_GEN_1763 & _GEN_104168 : ~(_GEN_104509 & _GEN_1763) & _GEN_104168) : _GEN_104168;
  wire        _GEN_104403 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1764 & _GEN_104169 : _GEN_1053 ? ~_GEN_1764 & _GEN_104169 : ~(_GEN_104509 & _GEN_1764) & _GEN_104169) : _GEN_104169;
  wire        _GEN_104404 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1765 & _GEN_104170 : _GEN_1053 ? ~_GEN_1765 & _GEN_104170 : ~(_GEN_104509 & _GEN_1765) & _GEN_104170) : _GEN_104170;
  wire        _GEN_104405 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1766 & _GEN_104171 : _GEN_1053 ? ~_GEN_1766 & _GEN_104171 : ~(_GEN_104509 & _GEN_1766) & _GEN_104171) : _GEN_104171;
  wire        _GEN_104406 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1767 & _GEN_104172 : _GEN_1053 ? ~_GEN_1767 & _GEN_104172 : ~(_GEN_104509 & _GEN_1767) & _GEN_104172) : _GEN_104172;
  wire        _GEN_104407 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1768 & _GEN_104173 : _GEN_1053 ? ~_GEN_1768 & _GEN_104173 : ~(_GEN_104509 & _GEN_1768) & _GEN_104173) : _GEN_104173;
  wire        _GEN_104408 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1769 & _GEN_104174 : _GEN_1053 ? ~_GEN_1769 & _GEN_104174 : ~(_GEN_104509 & _GEN_1769) & _GEN_104174) : _GEN_104174;
  wire        _GEN_104409 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1770 & _GEN_104175 : _GEN_1053 ? ~_GEN_1770 & _GEN_104175 : ~(_GEN_104509 & _GEN_1770) & _GEN_104175) : _GEN_104175;
  wire        _GEN_104410 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1771 & _GEN_104176 : _GEN_1053 ? ~_GEN_1771 & _GEN_104176 : ~(_GEN_104509 & _GEN_1771) & _GEN_104176) : _GEN_104176;
  wire        _GEN_104411 = _GEN_1051 ? (_GEN_104344 ? ~_GEN_1772 & _GEN_104177 : _GEN_1053 ? ~_GEN_1772 & _GEN_104177 : ~(_GEN_104509 & _GEN_1772) & _GEN_104177) : _GEN_104177;
  wire        _GEN_104412 = _GEN_1051 ? (_GEN_104344 ? ~(&lcam_ldq_idx_0) & _GEN_104178 : _GEN_1053 ? ~(&lcam_ldq_idx_0) & _GEN_104178 : ~(_GEN_104509 & (&lcam_ldq_idx_0)) & _GEN_104178) : _GEN_104178;
  wire        _GEN_104615 = _GEN_1054 ? (_GEN_104578 ? (|lcam_ldq_idx_1) & _GEN_104381 : _GEN_1056 ? (|lcam_ldq_idx_1) & _GEN_104381 : ~(_GEN_104509 & ~(|lcam_ldq_idx_1)) & _GEN_104381) : _GEN_104381;
  wire        _GEN_104616 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1773 & _GEN_104382 : _GEN_1056 ? ~_GEN_1773 & _GEN_104382 : ~(_GEN_104509 & _GEN_1773) & _GEN_104382) : _GEN_104382;
  wire        _GEN_104617 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1774 & _GEN_104383 : _GEN_1056 ? ~_GEN_1774 & _GEN_104383 : ~(_GEN_104509 & _GEN_1774) & _GEN_104383) : _GEN_104383;
  wire        _GEN_104618 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1775 & _GEN_104384 : _GEN_1056 ? ~_GEN_1775 & _GEN_104384 : ~(_GEN_104509 & _GEN_1775) & _GEN_104384) : _GEN_104384;
  wire        _GEN_104619 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1776 & _GEN_104385 : _GEN_1056 ? ~_GEN_1776 & _GEN_104385 : ~(_GEN_104509 & _GEN_1776) & _GEN_104385) : _GEN_104385;
  wire        _GEN_104620 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1777 & _GEN_104386 : _GEN_1056 ? ~_GEN_1777 & _GEN_104386 : ~(_GEN_104509 & _GEN_1777) & _GEN_104386) : _GEN_104386;
  wire        _GEN_104621 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1778 & _GEN_104387 : _GEN_1056 ? ~_GEN_1778 & _GEN_104387 : ~(_GEN_104509 & _GEN_1778) & _GEN_104387) : _GEN_104387;
  wire        _GEN_104622 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1779 & _GEN_104388 : _GEN_1056 ? ~_GEN_1779 & _GEN_104388 : ~(_GEN_104509 & _GEN_1779) & _GEN_104388) : _GEN_104388;
  wire        _GEN_104623 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1780 & _GEN_104389 : _GEN_1056 ? ~_GEN_1780 & _GEN_104389 : ~(_GEN_104509 & _GEN_1780) & _GEN_104389) : _GEN_104389;
  wire        _GEN_104624 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1781 & _GEN_104390 : _GEN_1056 ? ~_GEN_1781 & _GEN_104390 : ~(_GEN_104509 & _GEN_1781) & _GEN_104390) : _GEN_104390;
  wire        _GEN_104625 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1782 & _GEN_104391 : _GEN_1056 ? ~_GEN_1782 & _GEN_104391 : ~(_GEN_104509 & _GEN_1782) & _GEN_104391) : _GEN_104391;
  wire        _GEN_104626 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1783 & _GEN_104392 : _GEN_1056 ? ~_GEN_1783 & _GEN_104392 : ~(_GEN_104509 & _GEN_1783) & _GEN_104392) : _GEN_104392;
  wire        _GEN_104627 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1784 & _GEN_104393 : _GEN_1056 ? ~_GEN_1784 & _GEN_104393 : ~(_GEN_104509 & _GEN_1784) & _GEN_104393) : _GEN_104393;
  wire        _GEN_104628 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1785 & _GEN_104394 : _GEN_1056 ? ~_GEN_1785 & _GEN_104394 : ~(_GEN_104509 & _GEN_1785) & _GEN_104394) : _GEN_104394;
  wire        _GEN_104629 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1786 & _GEN_104395 : _GEN_1056 ? ~_GEN_1786 & _GEN_104395 : ~(_GEN_104509 & _GEN_1786) & _GEN_104395) : _GEN_104395;
  wire        _GEN_104630 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1787 & _GEN_104396 : _GEN_1056 ? ~_GEN_1787 & _GEN_104396 : ~(_GEN_104509 & _GEN_1787) & _GEN_104396) : _GEN_104396;
  wire        _GEN_104631 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1788 & _GEN_104397 : _GEN_1056 ? ~_GEN_1788 & _GEN_104397 : ~(_GEN_104509 & _GEN_1788) & _GEN_104397) : _GEN_104397;
  wire        _GEN_104632 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1789 & _GEN_104398 : _GEN_1056 ? ~_GEN_1789 & _GEN_104398 : ~(_GEN_104509 & _GEN_1789) & _GEN_104398) : _GEN_104398;
  wire        _GEN_104633 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1790 & _GEN_104399 : _GEN_1056 ? ~_GEN_1790 & _GEN_104399 : ~(_GEN_104509 & _GEN_1790) & _GEN_104399) : _GEN_104399;
  wire        _GEN_104634 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1791 & _GEN_104400 : _GEN_1056 ? ~_GEN_1791 & _GEN_104400 : ~(_GEN_104509 & _GEN_1791) & _GEN_104400) : _GEN_104400;
  wire        _GEN_104635 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1792 & _GEN_104401 : _GEN_1056 ? ~_GEN_1792 & _GEN_104401 : ~(_GEN_104509 & _GEN_1792) & _GEN_104401) : _GEN_104401;
  wire        _GEN_104636 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1793 & _GEN_104402 : _GEN_1056 ? ~_GEN_1793 & _GEN_104402 : ~(_GEN_104509 & _GEN_1793) & _GEN_104402) : _GEN_104402;
  wire        _GEN_104637 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1794 & _GEN_104403 : _GEN_1056 ? ~_GEN_1794 & _GEN_104403 : ~(_GEN_104509 & _GEN_1794) & _GEN_104403) : _GEN_104403;
  wire        _GEN_104638 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1795 & _GEN_104404 : _GEN_1056 ? ~_GEN_1795 & _GEN_104404 : ~(_GEN_104509 & _GEN_1795) & _GEN_104404) : _GEN_104404;
  wire        _GEN_104639 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1796 & _GEN_104405 : _GEN_1056 ? ~_GEN_1796 & _GEN_104405 : ~(_GEN_104509 & _GEN_1796) & _GEN_104405) : _GEN_104405;
  wire        _GEN_104640 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1797 & _GEN_104406 : _GEN_1056 ? ~_GEN_1797 & _GEN_104406 : ~(_GEN_104509 & _GEN_1797) & _GEN_104406) : _GEN_104406;
  wire        _GEN_104641 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1798 & _GEN_104407 : _GEN_1056 ? ~_GEN_1798 & _GEN_104407 : ~(_GEN_104509 & _GEN_1798) & _GEN_104407) : _GEN_104407;
  wire        _GEN_104642 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1799 & _GEN_104408 : _GEN_1056 ? ~_GEN_1799 & _GEN_104408 : ~(_GEN_104509 & _GEN_1799) & _GEN_104408) : _GEN_104408;
  wire        _GEN_104643 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1800 & _GEN_104409 : _GEN_1056 ? ~_GEN_1800 & _GEN_104409 : ~(_GEN_104509 & _GEN_1800) & _GEN_104409) : _GEN_104409;
  wire        _GEN_104644 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1801 & _GEN_104410 : _GEN_1056 ? ~_GEN_1801 & _GEN_104410 : ~(_GEN_104509 & _GEN_1801) & _GEN_104410) : _GEN_104410;
  wire        _GEN_104645 = _GEN_1054 ? (_GEN_104578 ? ~_GEN_1802 & _GEN_104411 : _GEN_1056 ? ~_GEN_1802 & _GEN_104411 : ~(_GEN_104509 & _GEN_1802) & _GEN_104411) : _GEN_104411;
  wire        _GEN_104646 = _GEN_1054 ? (_GEN_104578 ? ~(&lcam_ldq_idx_1) & _GEN_104412 : _GEN_1056 ? ~(&lcam_ldq_idx_1) & _GEN_104412 : ~(_GEN_104509 & (&lcam_ldq_idx_1)) & _GEN_104412) : _GEN_104412;
  wire        _GEN_104849 = _GEN_1057 ? (_GEN_104812 ? (|lcam_ldq_idx_0) & _GEN_104615 : _GEN_1059 ? (|lcam_ldq_idx_0) & _GEN_104615 : ~(_GEN_104977 & ~(|lcam_ldq_idx_0)) & _GEN_104615) : _GEN_104615;
  wire        _GEN_104850 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1743 & _GEN_104616 : _GEN_1059 ? ~_GEN_1743 & _GEN_104616 : ~(_GEN_104977 & _GEN_1743) & _GEN_104616) : _GEN_104616;
  wire        _GEN_104851 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1744 & _GEN_104617 : _GEN_1059 ? ~_GEN_1744 & _GEN_104617 : ~(_GEN_104977 & _GEN_1744) & _GEN_104617) : _GEN_104617;
  wire        _GEN_104852 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1745 & _GEN_104618 : _GEN_1059 ? ~_GEN_1745 & _GEN_104618 : ~(_GEN_104977 & _GEN_1745) & _GEN_104618) : _GEN_104618;
  wire        _GEN_104853 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1746 & _GEN_104619 : _GEN_1059 ? ~_GEN_1746 & _GEN_104619 : ~(_GEN_104977 & _GEN_1746) & _GEN_104619) : _GEN_104619;
  wire        _GEN_104854 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1747 & _GEN_104620 : _GEN_1059 ? ~_GEN_1747 & _GEN_104620 : ~(_GEN_104977 & _GEN_1747) & _GEN_104620) : _GEN_104620;
  wire        _GEN_104855 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1748 & _GEN_104621 : _GEN_1059 ? ~_GEN_1748 & _GEN_104621 : ~(_GEN_104977 & _GEN_1748) & _GEN_104621) : _GEN_104621;
  wire        _GEN_104856 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1749 & _GEN_104622 : _GEN_1059 ? ~_GEN_1749 & _GEN_104622 : ~(_GEN_104977 & _GEN_1749) & _GEN_104622) : _GEN_104622;
  wire        _GEN_104857 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1750 & _GEN_104623 : _GEN_1059 ? ~_GEN_1750 & _GEN_104623 : ~(_GEN_104977 & _GEN_1750) & _GEN_104623) : _GEN_104623;
  wire        _GEN_104858 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1751 & _GEN_104624 : _GEN_1059 ? ~_GEN_1751 & _GEN_104624 : ~(_GEN_104977 & _GEN_1751) & _GEN_104624) : _GEN_104624;
  wire        _GEN_104859 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1752 & _GEN_104625 : _GEN_1059 ? ~_GEN_1752 & _GEN_104625 : ~(_GEN_104977 & _GEN_1752) & _GEN_104625) : _GEN_104625;
  wire        _GEN_104860 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1753 & _GEN_104626 : _GEN_1059 ? ~_GEN_1753 & _GEN_104626 : ~(_GEN_104977 & _GEN_1753) & _GEN_104626) : _GEN_104626;
  wire        _GEN_104861 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1754 & _GEN_104627 : _GEN_1059 ? ~_GEN_1754 & _GEN_104627 : ~(_GEN_104977 & _GEN_1754) & _GEN_104627) : _GEN_104627;
  wire        _GEN_104862 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1755 & _GEN_104628 : _GEN_1059 ? ~_GEN_1755 & _GEN_104628 : ~(_GEN_104977 & _GEN_1755) & _GEN_104628) : _GEN_104628;
  wire        _GEN_104863 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1756 & _GEN_104629 : _GEN_1059 ? ~_GEN_1756 & _GEN_104629 : ~(_GEN_104977 & _GEN_1756) & _GEN_104629) : _GEN_104629;
  wire        _GEN_104864 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1757 & _GEN_104630 : _GEN_1059 ? ~_GEN_1757 & _GEN_104630 : ~(_GEN_104977 & _GEN_1757) & _GEN_104630) : _GEN_104630;
  wire        _GEN_104865 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1758 & _GEN_104631 : _GEN_1059 ? ~_GEN_1758 & _GEN_104631 : ~(_GEN_104977 & _GEN_1758) & _GEN_104631) : _GEN_104631;
  wire        _GEN_104866 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1759 & _GEN_104632 : _GEN_1059 ? ~_GEN_1759 & _GEN_104632 : ~(_GEN_104977 & _GEN_1759) & _GEN_104632) : _GEN_104632;
  wire        _GEN_104867 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1760 & _GEN_104633 : _GEN_1059 ? ~_GEN_1760 & _GEN_104633 : ~(_GEN_104977 & _GEN_1760) & _GEN_104633) : _GEN_104633;
  wire        _GEN_104868 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1761 & _GEN_104634 : _GEN_1059 ? ~_GEN_1761 & _GEN_104634 : ~(_GEN_104977 & _GEN_1761) & _GEN_104634) : _GEN_104634;
  wire        _GEN_104869 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1762 & _GEN_104635 : _GEN_1059 ? ~_GEN_1762 & _GEN_104635 : ~(_GEN_104977 & _GEN_1762) & _GEN_104635) : _GEN_104635;
  wire        _GEN_104870 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1763 & _GEN_104636 : _GEN_1059 ? ~_GEN_1763 & _GEN_104636 : ~(_GEN_104977 & _GEN_1763) & _GEN_104636) : _GEN_104636;
  wire        _GEN_104871 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1764 & _GEN_104637 : _GEN_1059 ? ~_GEN_1764 & _GEN_104637 : ~(_GEN_104977 & _GEN_1764) & _GEN_104637) : _GEN_104637;
  wire        _GEN_104872 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1765 & _GEN_104638 : _GEN_1059 ? ~_GEN_1765 & _GEN_104638 : ~(_GEN_104977 & _GEN_1765) & _GEN_104638) : _GEN_104638;
  wire        _GEN_104873 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1766 & _GEN_104639 : _GEN_1059 ? ~_GEN_1766 & _GEN_104639 : ~(_GEN_104977 & _GEN_1766) & _GEN_104639) : _GEN_104639;
  wire        _GEN_104874 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1767 & _GEN_104640 : _GEN_1059 ? ~_GEN_1767 & _GEN_104640 : ~(_GEN_104977 & _GEN_1767) & _GEN_104640) : _GEN_104640;
  wire        _GEN_104875 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1768 & _GEN_104641 : _GEN_1059 ? ~_GEN_1768 & _GEN_104641 : ~(_GEN_104977 & _GEN_1768) & _GEN_104641) : _GEN_104641;
  wire        _GEN_104876 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1769 & _GEN_104642 : _GEN_1059 ? ~_GEN_1769 & _GEN_104642 : ~(_GEN_104977 & _GEN_1769) & _GEN_104642) : _GEN_104642;
  wire        _GEN_104877 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1770 & _GEN_104643 : _GEN_1059 ? ~_GEN_1770 & _GEN_104643 : ~(_GEN_104977 & _GEN_1770) & _GEN_104643) : _GEN_104643;
  wire        _GEN_104878 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1771 & _GEN_104644 : _GEN_1059 ? ~_GEN_1771 & _GEN_104644 : ~(_GEN_104977 & _GEN_1771) & _GEN_104644) : _GEN_104644;
  wire        _GEN_104879 = _GEN_1057 ? (_GEN_104812 ? ~_GEN_1772 & _GEN_104645 : _GEN_1059 ? ~_GEN_1772 & _GEN_104645 : ~(_GEN_104977 & _GEN_1772) & _GEN_104645) : _GEN_104645;
  wire        _GEN_104880 = _GEN_1057 ? (_GEN_104812 ? ~(&lcam_ldq_idx_0) & _GEN_104646 : _GEN_1059 ? ~(&lcam_ldq_idx_0) & _GEN_104646 : ~(_GEN_104977 & (&lcam_ldq_idx_0)) & _GEN_104646) : _GEN_104646;
  wire        _GEN_105083 = _GEN_1060 ? (_GEN_105046 ? (|lcam_ldq_idx_1) & _GEN_104849 : _GEN_1062 ? (|lcam_ldq_idx_1) & _GEN_104849 : ~(_GEN_104977 & ~(|lcam_ldq_idx_1)) & _GEN_104849) : _GEN_104849;
  wire        _GEN_105084 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1773 & _GEN_104850 : _GEN_1062 ? ~_GEN_1773 & _GEN_104850 : ~(_GEN_104977 & _GEN_1773) & _GEN_104850) : _GEN_104850;
  wire        _GEN_105085 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1774 & _GEN_104851 : _GEN_1062 ? ~_GEN_1774 & _GEN_104851 : ~(_GEN_104977 & _GEN_1774) & _GEN_104851) : _GEN_104851;
  wire        _GEN_105086 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1775 & _GEN_104852 : _GEN_1062 ? ~_GEN_1775 & _GEN_104852 : ~(_GEN_104977 & _GEN_1775) & _GEN_104852) : _GEN_104852;
  wire        _GEN_105087 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1776 & _GEN_104853 : _GEN_1062 ? ~_GEN_1776 & _GEN_104853 : ~(_GEN_104977 & _GEN_1776) & _GEN_104853) : _GEN_104853;
  wire        _GEN_105088 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1777 & _GEN_104854 : _GEN_1062 ? ~_GEN_1777 & _GEN_104854 : ~(_GEN_104977 & _GEN_1777) & _GEN_104854) : _GEN_104854;
  wire        _GEN_105089 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1778 & _GEN_104855 : _GEN_1062 ? ~_GEN_1778 & _GEN_104855 : ~(_GEN_104977 & _GEN_1778) & _GEN_104855) : _GEN_104855;
  wire        _GEN_105090 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1779 & _GEN_104856 : _GEN_1062 ? ~_GEN_1779 & _GEN_104856 : ~(_GEN_104977 & _GEN_1779) & _GEN_104856) : _GEN_104856;
  wire        _GEN_105091 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1780 & _GEN_104857 : _GEN_1062 ? ~_GEN_1780 & _GEN_104857 : ~(_GEN_104977 & _GEN_1780) & _GEN_104857) : _GEN_104857;
  wire        _GEN_105092 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1781 & _GEN_104858 : _GEN_1062 ? ~_GEN_1781 & _GEN_104858 : ~(_GEN_104977 & _GEN_1781) & _GEN_104858) : _GEN_104858;
  wire        _GEN_105093 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1782 & _GEN_104859 : _GEN_1062 ? ~_GEN_1782 & _GEN_104859 : ~(_GEN_104977 & _GEN_1782) & _GEN_104859) : _GEN_104859;
  wire        _GEN_105094 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1783 & _GEN_104860 : _GEN_1062 ? ~_GEN_1783 & _GEN_104860 : ~(_GEN_104977 & _GEN_1783) & _GEN_104860) : _GEN_104860;
  wire        _GEN_105095 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1784 & _GEN_104861 : _GEN_1062 ? ~_GEN_1784 & _GEN_104861 : ~(_GEN_104977 & _GEN_1784) & _GEN_104861) : _GEN_104861;
  wire        _GEN_105096 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1785 & _GEN_104862 : _GEN_1062 ? ~_GEN_1785 & _GEN_104862 : ~(_GEN_104977 & _GEN_1785) & _GEN_104862) : _GEN_104862;
  wire        _GEN_105097 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1786 & _GEN_104863 : _GEN_1062 ? ~_GEN_1786 & _GEN_104863 : ~(_GEN_104977 & _GEN_1786) & _GEN_104863) : _GEN_104863;
  wire        _GEN_105098 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1787 & _GEN_104864 : _GEN_1062 ? ~_GEN_1787 & _GEN_104864 : ~(_GEN_104977 & _GEN_1787) & _GEN_104864) : _GEN_104864;
  wire        _GEN_105099 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1788 & _GEN_104865 : _GEN_1062 ? ~_GEN_1788 & _GEN_104865 : ~(_GEN_104977 & _GEN_1788) & _GEN_104865) : _GEN_104865;
  wire        _GEN_105100 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1789 & _GEN_104866 : _GEN_1062 ? ~_GEN_1789 & _GEN_104866 : ~(_GEN_104977 & _GEN_1789) & _GEN_104866) : _GEN_104866;
  wire        _GEN_105101 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1790 & _GEN_104867 : _GEN_1062 ? ~_GEN_1790 & _GEN_104867 : ~(_GEN_104977 & _GEN_1790) & _GEN_104867) : _GEN_104867;
  wire        _GEN_105102 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1791 & _GEN_104868 : _GEN_1062 ? ~_GEN_1791 & _GEN_104868 : ~(_GEN_104977 & _GEN_1791) & _GEN_104868) : _GEN_104868;
  wire        _GEN_105103 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1792 & _GEN_104869 : _GEN_1062 ? ~_GEN_1792 & _GEN_104869 : ~(_GEN_104977 & _GEN_1792) & _GEN_104869) : _GEN_104869;
  wire        _GEN_105104 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1793 & _GEN_104870 : _GEN_1062 ? ~_GEN_1793 & _GEN_104870 : ~(_GEN_104977 & _GEN_1793) & _GEN_104870) : _GEN_104870;
  wire        _GEN_105105 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1794 & _GEN_104871 : _GEN_1062 ? ~_GEN_1794 & _GEN_104871 : ~(_GEN_104977 & _GEN_1794) & _GEN_104871) : _GEN_104871;
  wire        _GEN_105106 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1795 & _GEN_104872 : _GEN_1062 ? ~_GEN_1795 & _GEN_104872 : ~(_GEN_104977 & _GEN_1795) & _GEN_104872) : _GEN_104872;
  wire        _GEN_105107 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1796 & _GEN_104873 : _GEN_1062 ? ~_GEN_1796 & _GEN_104873 : ~(_GEN_104977 & _GEN_1796) & _GEN_104873) : _GEN_104873;
  wire        _GEN_105108 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1797 & _GEN_104874 : _GEN_1062 ? ~_GEN_1797 & _GEN_104874 : ~(_GEN_104977 & _GEN_1797) & _GEN_104874) : _GEN_104874;
  wire        _GEN_105109 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1798 & _GEN_104875 : _GEN_1062 ? ~_GEN_1798 & _GEN_104875 : ~(_GEN_104977 & _GEN_1798) & _GEN_104875) : _GEN_104875;
  wire        _GEN_105110 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1799 & _GEN_104876 : _GEN_1062 ? ~_GEN_1799 & _GEN_104876 : ~(_GEN_104977 & _GEN_1799) & _GEN_104876) : _GEN_104876;
  wire        _GEN_105111 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1800 & _GEN_104877 : _GEN_1062 ? ~_GEN_1800 & _GEN_104877 : ~(_GEN_104977 & _GEN_1800) & _GEN_104877) : _GEN_104877;
  wire        _GEN_105112 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1801 & _GEN_104878 : _GEN_1062 ? ~_GEN_1801 & _GEN_104878 : ~(_GEN_104977 & _GEN_1801) & _GEN_104878) : _GEN_104878;
  wire        _GEN_105113 = _GEN_1060 ? (_GEN_105046 ? ~_GEN_1802 & _GEN_104879 : _GEN_1062 ? ~_GEN_1802 & _GEN_104879 : ~(_GEN_104977 & _GEN_1802) & _GEN_104879) : _GEN_104879;
  wire        _GEN_105114 = _GEN_1060 ? (_GEN_105046 ? ~(&lcam_ldq_idx_1) & _GEN_104880 : _GEN_1062 ? ~(&lcam_ldq_idx_1) & _GEN_104880 : ~(_GEN_104977 & (&lcam_ldq_idx_1)) & _GEN_104880) : _GEN_104880;
  wire        _GEN_105317 = _GEN_1063 ? (_GEN_105280 ? (|lcam_ldq_idx_0) & _GEN_105083 : _GEN_1065 ? (|lcam_ldq_idx_0) & _GEN_105083 : ~(_GEN_105445 & ~(|lcam_ldq_idx_0)) & _GEN_105083) : _GEN_105083;
  wire        _GEN_105318 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1743 & _GEN_105084 : _GEN_1065 ? ~_GEN_1743 & _GEN_105084 : ~(_GEN_105445 & _GEN_1743) & _GEN_105084) : _GEN_105084;
  wire        _GEN_105319 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1744 & _GEN_105085 : _GEN_1065 ? ~_GEN_1744 & _GEN_105085 : ~(_GEN_105445 & _GEN_1744) & _GEN_105085) : _GEN_105085;
  wire        _GEN_105320 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1745 & _GEN_105086 : _GEN_1065 ? ~_GEN_1745 & _GEN_105086 : ~(_GEN_105445 & _GEN_1745) & _GEN_105086) : _GEN_105086;
  wire        _GEN_105321 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1746 & _GEN_105087 : _GEN_1065 ? ~_GEN_1746 & _GEN_105087 : ~(_GEN_105445 & _GEN_1746) & _GEN_105087) : _GEN_105087;
  wire        _GEN_105322 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1747 & _GEN_105088 : _GEN_1065 ? ~_GEN_1747 & _GEN_105088 : ~(_GEN_105445 & _GEN_1747) & _GEN_105088) : _GEN_105088;
  wire        _GEN_105323 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1748 & _GEN_105089 : _GEN_1065 ? ~_GEN_1748 & _GEN_105089 : ~(_GEN_105445 & _GEN_1748) & _GEN_105089) : _GEN_105089;
  wire        _GEN_105324 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1749 & _GEN_105090 : _GEN_1065 ? ~_GEN_1749 & _GEN_105090 : ~(_GEN_105445 & _GEN_1749) & _GEN_105090) : _GEN_105090;
  wire        _GEN_105325 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1750 & _GEN_105091 : _GEN_1065 ? ~_GEN_1750 & _GEN_105091 : ~(_GEN_105445 & _GEN_1750) & _GEN_105091) : _GEN_105091;
  wire        _GEN_105326 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1751 & _GEN_105092 : _GEN_1065 ? ~_GEN_1751 & _GEN_105092 : ~(_GEN_105445 & _GEN_1751) & _GEN_105092) : _GEN_105092;
  wire        _GEN_105327 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1752 & _GEN_105093 : _GEN_1065 ? ~_GEN_1752 & _GEN_105093 : ~(_GEN_105445 & _GEN_1752) & _GEN_105093) : _GEN_105093;
  wire        _GEN_105328 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1753 & _GEN_105094 : _GEN_1065 ? ~_GEN_1753 & _GEN_105094 : ~(_GEN_105445 & _GEN_1753) & _GEN_105094) : _GEN_105094;
  wire        _GEN_105329 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1754 & _GEN_105095 : _GEN_1065 ? ~_GEN_1754 & _GEN_105095 : ~(_GEN_105445 & _GEN_1754) & _GEN_105095) : _GEN_105095;
  wire        _GEN_105330 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1755 & _GEN_105096 : _GEN_1065 ? ~_GEN_1755 & _GEN_105096 : ~(_GEN_105445 & _GEN_1755) & _GEN_105096) : _GEN_105096;
  wire        _GEN_105331 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1756 & _GEN_105097 : _GEN_1065 ? ~_GEN_1756 & _GEN_105097 : ~(_GEN_105445 & _GEN_1756) & _GEN_105097) : _GEN_105097;
  wire        _GEN_105332 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1757 & _GEN_105098 : _GEN_1065 ? ~_GEN_1757 & _GEN_105098 : ~(_GEN_105445 & _GEN_1757) & _GEN_105098) : _GEN_105098;
  wire        _GEN_105333 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1758 & _GEN_105099 : _GEN_1065 ? ~_GEN_1758 & _GEN_105099 : ~(_GEN_105445 & _GEN_1758) & _GEN_105099) : _GEN_105099;
  wire        _GEN_105334 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1759 & _GEN_105100 : _GEN_1065 ? ~_GEN_1759 & _GEN_105100 : ~(_GEN_105445 & _GEN_1759) & _GEN_105100) : _GEN_105100;
  wire        _GEN_105335 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1760 & _GEN_105101 : _GEN_1065 ? ~_GEN_1760 & _GEN_105101 : ~(_GEN_105445 & _GEN_1760) & _GEN_105101) : _GEN_105101;
  wire        _GEN_105336 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1761 & _GEN_105102 : _GEN_1065 ? ~_GEN_1761 & _GEN_105102 : ~(_GEN_105445 & _GEN_1761) & _GEN_105102) : _GEN_105102;
  wire        _GEN_105337 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1762 & _GEN_105103 : _GEN_1065 ? ~_GEN_1762 & _GEN_105103 : ~(_GEN_105445 & _GEN_1762) & _GEN_105103) : _GEN_105103;
  wire        _GEN_105338 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1763 & _GEN_105104 : _GEN_1065 ? ~_GEN_1763 & _GEN_105104 : ~(_GEN_105445 & _GEN_1763) & _GEN_105104) : _GEN_105104;
  wire        _GEN_105339 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1764 & _GEN_105105 : _GEN_1065 ? ~_GEN_1764 & _GEN_105105 : ~(_GEN_105445 & _GEN_1764) & _GEN_105105) : _GEN_105105;
  wire        _GEN_105340 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1765 & _GEN_105106 : _GEN_1065 ? ~_GEN_1765 & _GEN_105106 : ~(_GEN_105445 & _GEN_1765) & _GEN_105106) : _GEN_105106;
  wire        _GEN_105341 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1766 & _GEN_105107 : _GEN_1065 ? ~_GEN_1766 & _GEN_105107 : ~(_GEN_105445 & _GEN_1766) & _GEN_105107) : _GEN_105107;
  wire        _GEN_105342 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1767 & _GEN_105108 : _GEN_1065 ? ~_GEN_1767 & _GEN_105108 : ~(_GEN_105445 & _GEN_1767) & _GEN_105108) : _GEN_105108;
  wire        _GEN_105343 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1768 & _GEN_105109 : _GEN_1065 ? ~_GEN_1768 & _GEN_105109 : ~(_GEN_105445 & _GEN_1768) & _GEN_105109) : _GEN_105109;
  wire        _GEN_105344 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1769 & _GEN_105110 : _GEN_1065 ? ~_GEN_1769 & _GEN_105110 : ~(_GEN_105445 & _GEN_1769) & _GEN_105110) : _GEN_105110;
  wire        _GEN_105345 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1770 & _GEN_105111 : _GEN_1065 ? ~_GEN_1770 & _GEN_105111 : ~(_GEN_105445 & _GEN_1770) & _GEN_105111) : _GEN_105111;
  wire        _GEN_105346 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1771 & _GEN_105112 : _GEN_1065 ? ~_GEN_1771 & _GEN_105112 : ~(_GEN_105445 & _GEN_1771) & _GEN_105112) : _GEN_105112;
  wire        _GEN_105347 = _GEN_1063 ? (_GEN_105280 ? ~_GEN_1772 & _GEN_105113 : _GEN_1065 ? ~_GEN_1772 & _GEN_105113 : ~(_GEN_105445 & _GEN_1772) & _GEN_105113) : _GEN_105113;
  wire        _GEN_105348 = _GEN_1063 ? (_GEN_105280 ? ~(&lcam_ldq_idx_0) & _GEN_105114 : _GEN_1065 ? ~(&lcam_ldq_idx_0) & _GEN_105114 : ~(_GEN_105445 & (&lcam_ldq_idx_0)) & _GEN_105114) : _GEN_105114;
  wire        _GEN_105551 = _GEN_1066 ? (_GEN_105514 ? (|lcam_ldq_idx_1) & _GEN_105317 : _GEN_1068 ? (|lcam_ldq_idx_1) & _GEN_105317 : ~(_GEN_105445 & ~(|lcam_ldq_idx_1)) & _GEN_105317) : _GEN_105317;
  wire        _GEN_105552 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1773 & _GEN_105318 : _GEN_1068 ? ~_GEN_1773 & _GEN_105318 : ~(_GEN_105445 & _GEN_1773) & _GEN_105318) : _GEN_105318;
  wire        _GEN_105553 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1774 & _GEN_105319 : _GEN_1068 ? ~_GEN_1774 & _GEN_105319 : ~(_GEN_105445 & _GEN_1774) & _GEN_105319) : _GEN_105319;
  wire        _GEN_105554 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1775 & _GEN_105320 : _GEN_1068 ? ~_GEN_1775 & _GEN_105320 : ~(_GEN_105445 & _GEN_1775) & _GEN_105320) : _GEN_105320;
  wire        _GEN_105555 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1776 & _GEN_105321 : _GEN_1068 ? ~_GEN_1776 & _GEN_105321 : ~(_GEN_105445 & _GEN_1776) & _GEN_105321) : _GEN_105321;
  wire        _GEN_105556 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1777 & _GEN_105322 : _GEN_1068 ? ~_GEN_1777 & _GEN_105322 : ~(_GEN_105445 & _GEN_1777) & _GEN_105322) : _GEN_105322;
  wire        _GEN_105557 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1778 & _GEN_105323 : _GEN_1068 ? ~_GEN_1778 & _GEN_105323 : ~(_GEN_105445 & _GEN_1778) & _GEN_105323) : _GEN_105323;
  wire        _GEN_105558 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1779 & _GEN_105324 : _GEN_1068 ? ~_GEN_1779 & _GEN_105324 : ~(_GEN_105445 & _GEN_1779) & _GEN_105324) : _GEN_105324;
  wire        _GEN_105559 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1780 & _GEN_105325 : _GEN_1068 ? ~_GEN_1780 & _GEN_105325 : ~(_GEN_105445 & _GEN_1780) & _GEN_105325) : _GEN_105325;
  wire        _GEN_105560 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1781 & _GEN_105326 : _GEN_1068 ? ~_GEN_1781 & _GEN_105326 : ~(_GEN_105445 & _GEN_1781) & _GEN_105326) : _GEN_105326;
  wire        _GEN_105561 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1782 & _GEN_105327 : _GEN_1068 ? ~_GEN_1782 & _GEN_105327 : ~(_GEN_105445 & _GEN_1782) & _GEN_105327) : _GEN_105327;
  wire        _GEN_105562 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1783 & _GEN_105328 : _GEN_1068 ? ~_GEN_1783 & _GEN_105328 : ~(_GEN_105445 & _GEN_1783) & _GEN_105328) : _GEN_105328;
  wire        _GEN_105563 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1784 & _GEN_105329 : _GEN_1068 ? ~_GEN_1784 & _GEN_105329 : ~(_GEN_105445 & _GEN_1784) & _GEN_105329) : _GEN_105329;
  wire        _GEN_105564 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1785 & _GEN_105330 : _GEN_1068 ? ~_GEN_1785 & _GEN_105330 : ~(_GEN_105445 & _GEN_1785) & _GEN_105330) : _GEN_105330;
  wire        _GEN_105565 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1786 & _GEN_105331 : _GEN_1068 ? ~_GEN_1786 & _GEN_105331 : ~(_GEN_105445 & _GEN_1786) & _GEN_105331) : _GEN_105331;
  wire        _GEN_105566 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1787 & _GEN_105332 : _GEN_1068 ? ~_GEN_1787 & _GEN_105332 : ~(_GEN_105445 & _GEN_1787) & _GEN_105332) : _GEN_105332;
  wire        _GEN_105567 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1788 & _GEN_105333 : _GEN_1068 ? ~_GEN_1788 & _GEN_105333 : ~(_GEN_105445 & _GEN_1788) & _GEN_105333) : _GEN_105333;
  wire        _GEN_105568 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1789 & _GEN_105334 : _GEN_1068 ? ~_GEN_1789 & _GEN_105334 : ~(_GEN_105445 & _GEN_1789) & _GEN_105334) : _GEN_105334;
  wire        _GEN_105569 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1790 & _GEN_105335 : _GEN_1068 ? ~_GEN_1790 & _GEN_105335 : ~(_GEN_105445 & _GEN_1790) & _GEN_105335) : _GEN_105335;
  wire        _GEN_105570 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1791 & _GEN_105336 : _GEN_1068 ? ~_GEN_1791 & _GEN_105336 : ~(_GEN_105445 & _GEN_1791) & _GEN_105336) : _GEN_105336;
  wire        _GEN_105571 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1792 & _GEN_105337 : _GEN_1068 ? ~_GEN_1792 & _GEN_105337 : ~(_GEN_105445 & _GEN_1792) & _GEN_105337) : _GEN_105337;
  wire        _GEN_105572 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1793 & _GEN_105338 : _GEN_1068 ? ~_GEN_1793 & _GEN_105338 : ~(_GEN_105445 & _GEN_1793) & _GEN_105338) : _GEN_105338;
  wire        _GEN_105573 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1794 & _GEN_105339 : _GEN_1068 ? ~_GEN_1794 & _GEN_105339 : ~(_GEN_105445 & _GEN_1794) & _GEN_105339) : _GEN_105339;
  wire        _GEN_105574 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1795 & _GEN_105340 : _GEN_1068 ? ~_GEN_1795 & _GEN_105340 : ~(_GEN_105445 & _GEN_1795) & _GEN_105340) : _GEN_105340;
  wire        _GEN_105575 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1796 & _GEN_105341 : _GEN_1068 ? ~_GEN_1796 & _GEN_105341 : ~(_GEN_105445 & _GEN_1796) & _GEN_105341) : _GEN_105341;
  wire        _GEN_105576 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1797 & _GEN_105342 : _GEN_1068 ? ~_GEN_1797 & _GEN_105342 : ~(_GEN_105445 & _GEN_1797) & _GEN_105342) : _GEN_105342;
  wire        _GEN_105577 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1798 & _GEN_105343 : _GEN_1068 ? ~_GEN_1798 & _GEN_105343 : ~(_GEN_105445 & _GEN_1798) & _GEN_105343) : _GEN_105343;
  wire        _GEN_105578 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1799 & _GEN_105344 : _GEN_1068 ? ~_GEN_1799 & _GEN_105344 : ~(_GEN_105445 & _GEN_1799) & _GEN_105344) : _GEN_105344;
  wire        _GEN_105579 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1800 & _GEN_105345 : _GEN_1068 ? ~_GEN_1800 & _GEN_105345 : ~(_GEN_105445 & _GEN_1800) & _GEN_105345) : _GEN_105345;
  wire        _GEN_105580 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1801 & _GEN_105346 : _GEN_1068 ? ~_GEN_1801 & _GEN_105346 : ~(_GEN_105445 & _GEN_1801) & _GEN_105346) : _GEN_105346;
  wire        _GEN_105581 = _GEN_1066 ? (_GEN_105514 ? ~_GEN_1802 & _GEN_105347 : _GEN_1068 ? ~_GEN_1802 & _GEN_105347 : ~(_GEN_105445 & _GEN_1802) & _GEN_105347) : _GEN_105347;
  wire        _GEN_105582 = _GEN_1066 ? (_GEN_105514 ? ~(&lcam_ldq_idx_1) & _GEN_105348 : _GEN_1068 ? ~(&lcam_ldq_idx_1) & _GEN_105348 : ~(_GEN_105445 & (&lcam_ldq_idx_1)) & _GEN_105348) : _GEN_105348;
  wire        _GEN_105785 = _GEN_1069 ? (_GEN_105748 ? (|lcam_ldq_idx_0) & _GEN_105551 : _GEN_1071 ? (|lcam_ldq_idx_0) & _GEN_105551 : ~(_GEN_105913 & ~(|lcam_ldq_idx_0)) & _GEN_105551) : _GEN_105551;
  wire        _GEN_105786 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1743 & _GEN_105552 : _GEN_1071 ? ~_GEN_1743 & _GEN_105552 : ~(_GEN_105913 & _GEN_1743) & _GEN_105552) : _GEN_105552;
  wire        _GEN_105787 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1744 & _GEN_105553 : _GEN_1071 ? ~_GEN_1744 & _GEN_105553 : ~(_GEN_105913 & _GEN_1744) & _GEN_105553) : _GEN_105553;
  wire        _GEN_105788 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1745 & _GEN_105554 : _GEN_1071 ? ~_GEN_1745 & _GEN_105554 : ~(_GEN_105913 & _GEN_1745) & _GEN_105554) : _GEN_105554;
  wire        _GEN_105789 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1746 & _GEN_105555 : _GEN_1071 ? ~_GEN_1746 & _GEN_105555 : ~(_GEN_105913 & _GEN_1746) & _GEN_105555) : _GEN_105555;
  wire        _GEN_105790 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1747 & _GEN_105556 : _GEN_1071 ? ~_GEN_1747 & _GEN_105556 : ~(_GEN_105913 & _GEN_1747) & _GEN_105556) : _GEN_105556;
  wire        _GEN_105791 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1748 & _GEN_105557 : _GEN_1071 ? ~_GEN_1748 & _GEN_105557 : ~(_GEN_105913 & _GEN_1748) & _GEN_105557) : _GEN_105557;
  wire        _GEN_105792 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1749 & _GEN_105558 : _GEN_1071 ? ~_GEN_1749 & _GEN_105558 : ~(_GEN_105913 & _GEN_1749) & _GEN_105558) : _GEN_105558;
  wire        _GEN_105793 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1750 & _GEN_105559 : _GEN_1071 ? ~_GEN_1750 & _GEN_105559 : ~(_GEN_105913 & _GEN_1750) & _GEN_105559) : _GEN_105559;
  wire        _GEN_105794 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1751 & _GEN_105560 : _GEN_1071 ? ~_GEN_1751 & _GEN_105560 : ~(_GEN_105913 & _GEN_1751) & _GEN_105560) : _GEN_105560;
  wire        _GEN_105795 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1752 & _GEN_105561 : _GEN_1071 ? ~_GEN_1752 & _GEN_105561 : ~(_GEN_105913 & _GEN_1752) & _GEN_105561) : _GEN_105561;
  wire        _GEN_105796 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1753 & _GEN_105562 : _GEN_1071 ? ~_GEN_1753 & _GEN_105562 : ~(_GEN_105913 & _GEN_1753) & _GEN_105562) : _GEN_105562;
  wire        _GEN_105797 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1754 & _GEN_105563 : _GEN_1071 ? ~_GEN_1754 & _GEN_105563 : ~(_GEN_105913 & _GEN_1754) & _GEN_105563) : _GEN_105563;
  wire        _GEN_105798 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1755 & _GEN_105564 : _GEN_1071 ? ~_GEN_1755 & _GEN_105564 : ~(_GEN_105913 & _GEN_1755) & _GEN_105564) : _GEN_105564;
  wire        _GEN_105799 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1756 & _GEN_105565 : _GEN_1071 ? ~_GEN_1756 & _GEN_105565 : ~(_GEN_105913 & _GEN_1756) & _GEN_105565) : _GEN_105565;
  wire        _GEN_105800 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1757 & _GEN_105566 : _GEN_1071 ? ~_GEN_1757 & _GEN_105566 : ~(_GEN_105913 & _GEN_1757) & _GEN_105566) : _GEN_105566;
  wire        _GEN_105801 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1758 & _GEN_105567 : _GEN_1071 ? ~_GEN_1758 & _GEN_105567 : ~(_GEN_105913 & _GEN_1758) & _GEN_105567) : _GEN_105567;
  wire        _GEN_105802 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1759 & _GEN_105568 : _GEN_1071 ? ~_GEN_1759 & _GEN_105568 : ~(_GEN_105913 & _GEN_1759) & _GEN_105568) : _GEN_105568;
  wire        _GEN_105803 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1760 & _GEN_105569 : _GEN_1071 ? ~_GEN_1760 & _GEN_105569 : ~(_GEN_105913 & _GEN_1760) & _GEN_105569) : _GEN_105569;
  wire        _GEN_105804 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1761 & _GEN_105570 : _GEN_1071 ? ~_GEN_1761 & _GEN_105570 : ~(_GEN_105913 & _GEN_1761) & _GEN_105570) : _GEN_105570;
  wire        _GEN_105805 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1762 & _GEN_105571 : _GEN_1071 ? ~_GEN_1762 & _GEN_105571 : ~(_GEN_105913 & _GEN_1762) & _GEN_105571) : _GEN_105571;
  wire        _GEN_105806 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1763 & _GEN_105572 : _GEN_1071 ? ~_GEN_1763 & _GEN_105572 : ~(_GEN_105913 & _GEN_1763) & _GEN_105572) : _GEN_105572;
  wire        _GEN_105807 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1764 & _GEN_105573 : _GEN_1071 ? ~_GEN_1764 & _GEN_105573 : ~(_GEN_105913 & _GEN_1764) & _GEN_105573) : _GEN_105573;
  wire        _GEN_105808 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1765 & _GEN_105574 : _GEN_1071 ? ~_GEN_1765 & _GEN_105574 : ~(_GEN_105913 & _GEN_1765) & _GEN_105574) : _GEN_105574;
  wire        _GEN_105809 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1766 & _GEN_105575 : _GEN_1071 ? ~_GEN_1766 & _GEN_105575 : ~(_GEN_105913 & _GEN_1766) & _GEN_105575) : _GEN_105575;
  wire        _GEN_105810 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1767 & _GEN_105576 : _GEN_1071 ? ~_GEN_1767 & _GEN_105576 : ~(_GEN_105913 & _GEN_1767) & _GEN_105576) : _GEN_105576;
  wire        _GEN_105811 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1768 & _GEN_105577 : _GEN_1071 ? ~_GEN_1768 & _GEN_105577 : ~(_GEN_105913 & _GEN_1768) & _GEN_105577) : _GEN_105577;
  wire        _GEN_105812 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1769 & _GEN_105578 : _GEN_1071 ? ~_GEN_1769 & _GEN_105578 : ~(_GEN_105913 & _GEN_1769) & _GEN_105578) : _GEN_105578;
  wire        _GEN_105813 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1770 & _GEN_105579 : _GEN_1071 ? ~_GEN_1770 & _GEN_105579 : ~(_GEN_105913 & _GEN_1770) & _GEN_105579) : _GEN_105579;
  wire        _GEN_105814 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1771 & _GEN_105580 : _GEN_1071 ? ~_GEN_1771 & _GEN_105580 : ~(_GEN_105913 & _GEN_1771) & _GEN_105580) : _GEN_105580;
  wire        _GEN_105815 = _GEN_1069 ? (_GEN_105748 ? ~_GEN_1772 & _GEN_105581 : _GEN_1071 ? ~_GEN_1772 & _GEN_105581 : ~(_GEN_105913 & _GEN_1772) & _GEN_105581) : _GEN_105581;
  wire        _GEN_105816 = _GEN_1069 ? (_GEN_105748 ? ~(&lcam_ldq_idx_0) & _GEN_105582 : _GEN_1071 ? ~(&lcam_ldq_idx_0) & _GEN_105582 : ~(_GEN_105913 & (&lcam_ldq_idx_0)) & _GEN_105582) : _GEN_105582;
  wire        _GEN_106019 = _GEN_1072 ? (_GEN_105982 ? (|lcam_ldq_idx_1) & _GEN_105785 : _GEN_1074 ? (|lcam_ldq_idx_1) & _GEN_105785 : ~(_GEN_105913 & ~(|lcam_ldq_idx_1)) & _GEN_105785) : _GEN_105785;
  wire        _GEN_106020 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1773 & _GEN_105786 : _GEN_1074 ? ~_GEN_1773 & _GEN_105786 : ~(_GEN_105913 & _GEN_1773) & _GEN_105786) : _GEN_105786;
  wire        _GEN_106021 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1774 & _GEN_105787 : _GEN_1074 ? ~_GEN_1774 & _GEN_105787 : ~(_GEN_105913 & _GEN_1774) & _GEN_105787) : _GEN_105787;
  wire        _GEN_106022 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1775 & _GEN_105788 : _GEN_1074 ? ~_GEN_1775 & _GEN_105788 : ~(_GEN_105913 & _GEN_1775) & _GEN_105788) : _GEN_105788;
  wire        _GEN_106023 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1776 & _GEN_105789 : _GEN_1074 ? ~_GEN_1776 & _GEN_105789 : ~(_GEN_105913 & _GEN_1776) & _GEN_105789) : _GEN_105789;
  wire        _GEN_106024 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1777 & _GEN_105790 : _GEN_1074 ? ~_GEN_1777 & _GEN_105790 : ~(_GEN_105913 & _GEN_1777) & _GEN_105790) : _GEN_105790;
  wire        _GEN_106025 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1778 & _GEN_105791 : _GEN_1074 ? ~_GEN_1778 & _GEN_105791 : ~(_GEN_105913 & _GEN_1778) & _GEN_105791) : _GEN_105791;
  wire        _GEN_106026 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1779 & _GEN_105792 : _GEN_1074 ? ~_GEN_1779 & _GEN_105792 : ~(_GEN_105913 & _GEN_1779) & _GEN_105792) : _GEN_105792;
  wire        _GEN_106027 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1780 & _GEN_105793 : _GEN_1074 ? ~_GEN_1780 & _GEN_105793 : ~(_GEN_105913 & _GEN_1780) & _GEN_105793) : _GEN_105793;
  wire        _GEN_106028 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1781 & _GEN_105794 : _GEN_1074 ? ~_GEN_1781 & _GEN_105794 : ~(_GEN_105913 & _GEN_1781) & _GEN_105794) : _GEN_105794;
  wire        _GEN_106029 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1782 & _GEN_105795 : _GEN_1074 ? ~_GEN_1782 & _GEN_105795 : ~(_GEN_105913 & _GEN_1782) & _GEN_105795) : _GEN_105795;
  wire        _GEN_106030 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1783 & _GEN_105796 : _GEN_1074 ? ~_GEN_1783 & _GEN_105796 : ~(_GEN_105913 & _GEN_1783) & _GEN_105796) : _GEN_105796;
  wire        _GEN_106031 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1784 & _GEN_105797 : _GEN_1074 ? ~_GEN_1784 & _GEN_105797 : ~(_GEN_105913 & _GEN_1784) & _GEN_105797) : _GEN_105797;
  wire        _GEN_106032 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1785 & _GEN_105798 : _GEN_1074 ? ~_GEN_1785 & _GEN_105798 : ~(_GEN_105913 & _GEN_1785) & _GEN_105798) : _GEN_105798;
  wire        _GEN_106033 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1786 & _GEN_105799 : _GEN_1074 ? ~_GEN_1786 & _GEN_105799 : ~(_GEN_105913 & _GEN_1786) & _GEN_105799) : _GEN_105799;
  wire        _GEN_106034 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1787 & _GEN_105800 : _GEN_1074 ? ~_GEN_1787 & _GEN_105800 : ~(_GEN_105913 & _GEN_1787) & _GEN_105800) : _GEN_105800;
  wire        _GEN_106035 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1788 & _GEN_105801 : _GEN_1074 ? ~_GEN_1788 & _GEN_105801 : ~(_GEN_105913 & _GEN_1788) & _GEN_105801) : _GEN_105801;
  wire        _GEN_106036 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1789 & _GEN_105802 : _GEN_1074 ? ~_GEN_1789 & _GEN_105802 : ~(_GEN_105913 & _GEN_1789) & _GEN_105802) : _GEN_105802;
  wire        _GEN_106037 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1790 & _GEN_105803 : _GEN_1074 ? ~_GEN_1790 & _GEN_105803 : ~(_GEN_105913 & _GEN_1790) & _GEN_105803) : _GEN_105803;
  wire        _GEN_106038 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1791 & _GEN_105804 : _GEN_1074 ? ~_GEN_1791 & _GEN_105804 : ~(_GEN_105913 & _GEN_1791) & _GEN_105804) : _GEN_105804;
  wire        _GEN_106039 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1792 & _GEN_105805 : _GEN_1074 ? ~_GEN_1792 & _GEN_105805 : ~(_GEN_105913 & _GEN_1792) & _GEN_105805) : _GEN_105805;
  wire        _GEN_106040 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1793 & _GEN_105806 : _GEN_1074 ? ~_GEN_1793 & _GEN_105806 : ~(_GEN_105913 & _GEN_1793) & _GEN_105806) : _GEN_105806;
  wire        _GEN_106041 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1794 & _GEN_105807 : _GEN_1074 ? ~_GEN_1794 & _GEN_105807 : ~(_GEN_105913 & _GEN_1794) & _GEN_105807) : _GEN_105807;
  wire        _GEN_106042 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1795 & _GEN_105808 : _GEN_1074 ? ~_GEN_1795 & _GEN_105808 : ~(_GEN_105913 & _GEN_1795) & _GEN_105808) : _GEN_105808;
  wire        _GEN_106043 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1796 & _GEN_105809 : _GEN_1074 ? ~_GEN_1796 & _GEN_105809 : ~(_GEN_105913 & _GEN_1796) & _GEN_105809) : _GEN_105809;
  wire        _GEN_106044 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1797 & _GEN_105810 : _GEN_1074 ? ~_GEN_1797 & _GEN_105810 : ~(_GEN_105913 & _GEN_1797) & _GEN_105810) : _GEN_105810;
  wire        _GEN_106045 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1798 & _GEN_105811 : _GEN_1074 ? ~_GEN_1798 & _GEN_105811 : ~(_GEN_105913 & _GEN_1798) & _GEN_105811) : _GEN_105811;
  wire        _GEN_106046 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1799 & _GEN_105812 : _GEN_1074 ? ~_GEN_1799 & _GEN_105812 : ~(_GEN_105913 & _GEN_1799) & _GEN_105812) : _GEN_105812;
  wire        _GEN_106047 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1800 & _GEN_105813 : _GEN_1074 ? ~_GEN_1800 & _GEN_105813 : ~(_GEN_105913 & _GEN_1800) & _GEN_105813) : _GEN_105813;
  wire        _GEN_106048 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1801 & _GEN_105814 : _GEN_1074 ? ~_GEN_1801 & _GEN_105814 : ~(_GEN_105913 & _GEN_1801) & _GEN_105814) : _GEN_105814;
  wire        _GEN_106049 = _GEN_1072 ? (_GEN_105982 ? ~_GEN_1802 & _GEN_105815 : _GEN_1074 ? ~_GEN_1802 & _GEN_105815 : ~(_GEN_105913 & _GEN_1802) & _GEN_105815) : _GEN_105815;
  wire        _GEN_106050 = _GEN_1072 ? (_GEN_105982 ? ~(&lcam_ldq_idx_1) & _GEN_105816 : _GEN_1074 ? ~(&lcam_ldq_idx_1) & _GEN_105816 : ~(_GEN_105913 & (&lcam_ldq_idx_1)) & _GEN_105816) : _GEN_105816;
  wire        _GEN_106253 = _GEN_1075 ? (_GEN_106216 ? (|lcam_ldq_idx_0) & _GEN_106019 : _GEN_1077 ? (|lcam_ldq_idx_0) & _GEN_106019 : ~(_GEN_106381 & ~(|lcam_ldq_idx_0)) & _GEN_106019) : _GEN_106019;
  wire        _GEN_106254 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1743 & _GEN_106020 : _GEN_1077 ? ~_GEN_1743 & _GEN_106020 : ~(_GEN_106381 & _GEN_1743) & _GEN_106020) : _GEN_106020;
  wire        _GEN_106255 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1744 & _GEN_106021 : _GEN_1077 ? ~_GEN_1744 & _GEN_106021 : ~(_GEN_106381 & _GEN_1744) & _GEN_106021) : _GEN_106021;
  wire        _GEN_106256 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1745 & _GEN_106022 : _GEN_1077 ? ~_GEN_1745 & _GEN_106022 : ~(_GEN_106381 & _GEN_1745) & _GEN_106022) : _GEN_106022;
  wire        _GEN_106257 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1746 & _GEN_106023 : _GEN_1077 ? ~_GEN_1746 & _GEN_106023 : ~(_GEN_106381 & _GEN_1746) & _GEN_106023) : _GEN_106023;
  wire        _GEN_106258 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1747 & _GEN_106024 : _GEN_1077 ? ~_GEN_1747 & _GEN_106024 : ~(_GEN_106381 & _GEN_1747) & _GEN_106024) : _GEN_106024;
  wire        _GEN_106259 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1748 & _GEN_106025 : _GEN_1077 ? ~_GEN_1748 & _GEN_106025 : ~(_GEN_106381 & _GEN_1748) & _GEN_106025) : _GEN_106025;
  wire        _GEN_106260 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1749 & _GEN_106026 : _GEN_1077 ? ~_GEN_1749 & _GEN_106026 : ~(_GEN_106381 & _GEN_1749) & _GEN_106026) : _GEN_106026;
  wire        _GEN_106261 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1750 & _GEN_106027 : _GEN_1077 ? ~_GEN_1750 & _GEN_106027 : ~(_GEN_106381 & _GEN_1750) & _GEN_106027) : _GEN_106027;
  wire        _GEN_106262 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1751 & _GEN_106028 : _GEN_1077 ? ~_GEN_1751 & _GEN_106028 : ~(_GEN_106381 & _GEN_1751) & _GEN_106028) : _GEN_106028;
  wire        _GEN_106263 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1752 & _GEN_106029 : _GEN_1077 ? ~_GEN_1752 & _GEN_106029 : ~(_GEN_106381 & _GEN_1752) & _GEN_106029) : _GEN_106029;
  wire        _GEN_106264 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1753 & _GEN_106030 : _GEN_1077 ? ~_GEN_1753 & _GEN_106030 : ~(_GEN_106381 & _GEN_1753) & _GEN_106030) : _GEN_106030;
  wire        _GEN_106265 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1754 & _GEN_106031 : _GEN_1077 ? ~_GEN_1754 & _GEN_106031 : ~(_GEN_106381 & _GEN_1754) & _GEN_106031) : _GEN_106031;
  wire        _GEN_106266 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1755 & _GEN_106032 : _GEN_1077 ? ~_GEN_1755 & _GEN_106032 : ~(_GEN_106381 & _GEN_1755) & _GEN_106032) : _GEN_106032;
  wire        _GEN_106267 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1756 & _GEN_106033 : _GEN_1077 ? ~_GEN_1756 & _GEN_106033 : ~(_GEN_106381 & _GEN_1756) & _GEN_106033) : _GEN_106033;
  wire        _GEN_106268 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1757 & _GEN_106034 : _GEN_1077 ? ~_GEN_1757 & _GEN_106034 : ~(_GEN_106381 & _GEN_1757) & _GEN_106034) : _GEN_106034;
  wire        _GEN_106269 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1758 & _GEN_106035 : _GEN_1077 ? ~_GEN_1758 & _GEN_106035 : ~(_GEN_106381 & _GEN_1758) & _GEN_106035) : _GEN_106035;
  wire        _GEN_106270 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1759 & _GEN_106036 : _GEN_1077 ? ~_GEN_1759 & _GEN_106036 : ~(_GEN_106381 & _GEN_1759) & _GEN_106036) : _GEN_106036;
  wire        _GEN_106271 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1760 & _GEN_106037 : _GEN_1077 ? ~_GEN_1760 & _GEN_106037 : ~(_GEN_106381 & _GEN_1760) & _GEN_106037) : _GEN_106037;
  wire        _GEN_106272 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1761 & _GEN_106038 : _GEN_1077 ? ~_GEN_1761 & _GEN_106038 : ~(_GEN_106381 & _GEN_1761) & _GEN_106038) : _GEN_106038;
  wire        _GEN_106273 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1762 & _GEN_106039 : _GEN_1077 ? ~_GEN_1762 & _GEN_106039 : ~(_GEN_106381 & _GEN_1762) & _GEN_106039) : _GEN_106039;
  wire        _GEN_106274 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1763 & _GEN_106040 : _GEN_1077 ? ~_GEN_1763 & _GEN_106040 : ~(_GEN_106381 & _GEN_1763) & _GEN_106040) : _GEN_106040;
  wire        _GEN_106275 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1764 & _GEN_106041 : _GEN_1077 ? ~_GEN_1764 & _GEN_106041 : ~(_GEN_106381 & _GEN_1764) & _GEN_106041) : _GEN_106041;
  wire        _GEN_106276 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1765 & _GEN_106042 : _GEN_1077 ? ~_GEN_1765 & _GEN_106042 : ~(_GEN_106381 & _GEN_1765) & _GEN_106042) : _GEN_106042;
  wire        _GEN_106277 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1766 & _GEN_106043 : _GEN_1077 ? ~_GEN_1766 & _GEN_106043 : ~(_GEN_106381 & _GEN_1766) & _GEN_106043) : _GEN_106043;
  wire        _GEN_106278 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1767 & _GEN_106044 : _GEN_1077 ? ~_GEN_1767 & _GEN_106044 : ~(_GEN_106381 & _GEN_1767) & _GEN_106044) : _GEN_106044;
  wire        _GEN_106279 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1768 & _GEN_106045 : _GEN_1077 ? ~_GEN_1768 & _GEN_106045 : ~(_GEN_106381 & _GEN_1768) & _GEN_106045) : _GEN_106045;
  wire        _GEN_106280 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1769 & _GEN_106046 : _GEN_1077 ? ~_GEN_1769 & _GEN_106046 : ~(_GEN_106381 & _GEN_1769) & _GEN_106046) : _GEN_106046;
  wire        _GEN_106281 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1770 & _GEN_106047 : _GEN_1077 ? ~_GEN_1770 & _GEN_106047 : ~(_GEN_106381 & _GEN_1770) & _GEN_106047) : _GEN_106047;
  wire        _GEN_106282 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1771 & _GEN_106048 : _GEN_1077 ? ~_GEN_1771 & _GEN_106048 : ~(_GEN_106381 & _GEN_1771) & _GEN_106048) : _GEN_106048;
  wire        _GEN_106283 = _GEN_1075 ? (_GEN_106216 ? ~_GEN_1772 & _GEN_106049 : _GEN_1077 ? ~_GEN_1772 & _GEN_106049 : ~(_GEN_106381 & _GEN_1772) & _GEN_106049) : _GEN_106049;
  wire        _GEN_106284 = _GEN_1075 ? (_GEN_106216 ? ~(&lcam_ldq_idx_0) & _GEN_106050 : _GEN_1077 ? ~(&lcam_ldq_idx_0) & _GEN_106050 : ~(_GEN_106381 & (&lcam_ldq_idx_0)) & _GEN_106050) : _GEN_106050;
  wire        _GEN_106487 = _GEN_1078 ? (_GEN_106450 ? (|lcam_ldq_idx_1) & _GEN_106253 : _GEN_1080 ? (|lcam_ldq_idx_1) & _GEN_106253 : ~(_GEN_106381 & ~(|lcam_ldq_idx_1)) & _GEN_106253) : _GEN_106253;
  wire        _GEN_106488 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1773 & _GEN_106254 : _GEN_1080 ? ~_GEN_1773 & _GEN_106254 : ~(_GEN_106381 & _GEN_1773) & _GEN_106254) : _GEN_106254;
  wire        _GEN_106489 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1774 & _GEN_106255 : _GEN_1080 ? ~_GEN_1774 & _GEN_106255 : ~(_GEN_106381 & _GEN_1774) & _GEN_106255) : _GEN_106255;
  wire        _GEN_106490 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1775 & _GEN_106256 : _GEN_1080 ? ~_GEN_1775 & _GEN_106256 : ~(_GEN_106381 & _GEN_1775) & _GEN_106256) : _GEN_106256;
  wire        _GEN_106491 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1776 & _GEN_106257 : _GEN_1080 ? ~_GEN_1776 & _GEN_106257 : ~(_GEN_106381 & _GEN_1776) & _GEN_106257) : _GEN_106257;
  wire        _GEN_106492 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1777 & _GEN_106258 : _GEN_1080 ? ~_GEN_1777 & _GEN_106258 : ~(_GEN_106381 & _GEN_1777) & _GEN_106258) : _GEN_106258;
  wire        _GEN_106493 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1778 & _GEN_106259 : _GEN_1080 ? ~_GEN_1778 & _GEN_106259 : ~(_GEN_106381 & _GEN_1778) & _GEN_106259) : _GEN_106259;
  wire        _GEN_106494 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1779 & _GEN_106260 : _GEN_1080 ? ~_GEN_1779 & _GEN_106260 : ~(_GEN_106381 & _GEN_1779) & _GEN_106260) : _GEN_106260;
  wire        _GEN_106495 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1780 & _GEN_106261 : _GEN_1080 ? ~_GEN_1780 & _GEN_106261 : ~(_GEN_106381 & _GEN_1780) & _GEN_106261) : _GEN_106261;
  wire        _GEN_106496 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1781 & _GEN_106262 : _GEN_1080 ? ~_GEN_1781 & _GEN_106262 : ~(_GEN_106381 & _GEN_1781) & _GEN_106262) : _GEN_106262;
  wire        _GEN_106497 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1782 & _GEN_106263 : _GEN_1080 ? ~_GEN_1782 & _GEN_106263 : ~(_GEN_106381 & _GEN_1782) & _GEN_106263) : _GEN_106263;
  wire        _GEN_106498 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1783 & _GEN_106264 : _GEN_1080 ? ~_GEN_1783 & _GEN_106264 : ~(_GEN_106381 & _GEN_1783) & _GEN_106264) : _GEN_106264;
  wire        _GEN_106499 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1784 & _GEN_106265 : _GEN_1080 ? ~_GEN_1784 & _GEN_106265 : ~(_GEN_106381 & _GEN_1784) & _GEN_106265) : _GEN_106265;
  wire        _GEN_106500 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1785 & _GEN_106266 : _GEN_1080 ? ~_GEN_1785 & _GEN_106266 : ~(_GEN_106381 & _GEN_1785) & _GEN_106266) : _GEN_106266;
  wire        _GEN_106501 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1786 & _GEN_106267 : _GEN_1080 ? ~_GEN_1786 & _GEN_106267 : ~(_GEN_106381 & _GEN_1786) & _GEN_106267) : _GEN_106267;
  wire        _GEN_106502 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1787 & _GEN_106268 : _GEN_1080 ? ~_GEN_1787 & _GEN_106268 : ~(_GEN_106381 & _GEN_1787) & _GEN_106268) : _GEN_106268;
  wire        _GEN_106503 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1788 & _GEN_106269 : _GEN_1080 ? ~_GEN_1788 & _GEN_106269 : ~(_GEN_106381 & _GEN_1788) & _GEN_106269) : _GEN_106269;
  wire        _GEN_106504 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1789 & _GEN_106270 : _GEN_1080 ? ~_GEN_1789 & _GEN_106270 : ~(_GEN_106381 & _GEN_1789) & _GEN_106270) : _GEN_106270;
  wire        _GEN_106505 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1790 & _GEN_106271 : _GEN_1080 ? ~_GEN_1790 & _GEN_106271 : ~(_GEN_106381 & _GEN_1790) & _GEN_106271) : _GEN_106271;
  wire        _GEN_106506 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1791 & _GEN_106272 : _GEN_1080 ? ~_GEN_1791 & _GEN_106272 : ~(_GEN_106381 & _GEN_1791) & _GEN_106272) : _GEN_106272;
  wire        _GEN_106507 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1792 & _GEN_106273 : _GEN_1080 ? ~_GEN_1792 & _GEN_106273 : ~(_GEN_106381 & _GEN_1792) & _GEN_106273) : _GEN_106273;
  wire        _GEN_106508 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1793 & _GEN_106274 : _GEN_1080 ? ~_GEN_1793 & _GEN_106274 : ~(_GEN_106381 & _GEN_1793) & _GEN_106274) : _GEN_106274;
  wire        _GEN_106509 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1794 & _GEN_106275 : _GEN_1080 ? ~_GEN_1794 & _GEN_106275 : ~(_GEN_106381 & _GEN_1794) & _GEN_106275) : _GEN_106275;
  wire        _GEN_106510 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1795 & _GEN_106276 : _GEN_1080 ? ~_GEN_1795 & _GEN_106276 : ~(_GEN_106381 & _GEN_1795) & _GEN_106276) : _GEN_106276;
  wire        _GEN_106511 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1796 & _GEN_106277 : _GEN_1080 ? ~_GEN_1796 & _GEN_106277 : ~(_GEN_106381 & _GEN_1796) & _GEN_106277) : _GEN_106277;
  wire        _GEN_106512 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1797 & _GEN_106278 : _GEN_1080 ? ~_GEN_1797 & _GEN_106278 : ~(_GEN_106381 & _GEN_1797) & _GEN_106278) : _GEN_106278;
  wire        _GEN_106513 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1798 & _GEN_106279 : _GEN_1080 ? ~_GEN_1798 & _GEN_106279 : ~(_GEN_106381 & _GEN_1798) & _GEN_106279) : _GEN_106279;
  wire        _GEN_106514 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1799 & _GEN_106280 : _GEN_1080 ? ~_GEN_1799 & _GEN_106280 : ~(_GEN_106381 & _GEN_1799) & _GEN_106280) : _GEN_106280;
  wire        _GEN_106515 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1800 & _GEN_106281 : _GEN_1080 ? ~_GEN_1800 & _GEN_106281 : ~(_GEN_106381 & _GEN_1800) & _GEN_106281) : _GEN_106281;
  wire        _GEN_106516 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1801 & _GEN_106282 : _GEN_1080 ? ~_GEN_1801 & _GEN_106282 : ~(_GEN_106381 & _GEN_1801) & _GEN_106282) : _GEN_106282;
  wire        _GEN_106517 = _GEN_1078 ? (_GEN_106450 ? ~_GEN_1802 & _GEN_106283 : _GEN_1080 ? ~_GEN_1802 & _GEN_106283 : ~(_GEN_106381 & _GEN_1802) & _GEN_106283) : _GEN_106283;
  wire        _GEN_106518 = _GEN_1078 ? (_GEN_106450 ? ~(&lcam_ldq_idx_1) & _GEN_106284 : _GEN_1080 ? ~(&lcam_ldq_idx_1) & _GEN_106284 : ~(_GEN_106381 & (&lcam_ldq_idx_1)) & _GEN_106284) : _GEN_106284;
  wire        _GEN_106721 = _GEN_1081 ? (_GEN_106684 ? (|lcam_ldq_idx_0) & _GEN_106487 : _GEN_1083 ? (|lcam_ldq_idx_0) & _GEN_106487 : ~(_GEN_106849 & ~(|lcam_ldq_idx_0)) & _GEN_106487) : _GEN_106487;
  wire        _GEN_106722 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1743 & _GEN_106488 : _GEN_1083 ? ~_GEN_1743 & _GEN_106488 : ~(_GEN_106849 & _GEN_1743) & _GEN_106488) : _GEN_106488;
  wire        _GEN_106723 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1744 & _GEN_106489 : _GEN_1083 ? ~_GEN_1744 & _GEN_106489 : ~(_GEN_106849 & _GEN_1744) & _GEN_106489) : _GEN_106489;
  wire        _GEN_106724 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1745 & _GEN_106490 : _GEN_1083 ? ~_GEN_1745 & _GEN_106490 : ~(_GEN_106849 & _GEN_1745) & _GEN_106490) : _GEN_106490;
  wire        _GEN_106725 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1746 & _GEN_106491 : _GEN_1083 ? ~_GEN_1746 & _GEN_106491 : ~(_GEN_106849 & _GEN_1746) & _GEN_106491) : _GEN_106491;
  wire        _GEN_106726 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1747 & _GEN_106492 : _GEN_1083 ? ~_GEN_1747 & _GEN_106492 : ~(_GEN_106849 & _GEN_1747) & _GEN_106492) : _GEN_106492;
  wire        _GEN_106727 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1748 & _GEN_106493 : _GEN_1083 ? ~_GEN_1748 & _GEN_106493 : ~(_GEN_106849 & _GEN_1748) & _GEN_106493) : _GEN_106493;
  wire        _GEN_106728 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1749 & _GEN_106494 : _GEN_1083 ? ~_GEN_1749 & _GEN_106494 : ~(_GEN_106849 & _GEN_1749) & _GEN_106494) : _GEN_106494;
  wire        _GEN_106729 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1750 & _GEN_106495 : _GEN_1083 ? ~_GEN_1750 & _GEN_106495 : ~(_GEN_106849 & _GEN_1750) & _GEN_106495) : _GEN_106495;
  wire        _GEN_106730 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1751 & _GEN_106496 : _GEN_1083 ? ~_GEN_1751 & _GEN_106496 : ~(_GEN_106849 & _GEN_1751) & _GEN_106496) : _GEN_106496;
  wire        _GEN_106731 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1752 & _GEN_106497 : _GEN_1083 ? ~_GEN_1752 & _GEN_106497 : ~(_GEN_106849 & _GEN_1752) & _GEN_106497) : _GEN_106497;
  wire        _GEN_106732 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1753 & _GEN_106498 : _GEN_1083 ? ~_GEN_1753 & _GEN_106498 : ~(_GEN_106849 & _GEN_1753) & _GEN_106498) : _GEN_106498;
  wire        _GEN_106733 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1754 & _GEN_106499 : _GEN_1083 ? ~_GEN_1754 & _GEN_106499 : ~(_GEN_106849 & _GEN_1754) & _GEN_106499) : _GEN_106499;
  wire        _GEN_106734 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1755 & _GEN_106500 : _GEN_1083 ? ~_GEN_1755 & _GEN_106500 : ~(_GEN_106849 & _GEN_1755) & _GEN_106500) : _GEN_106500;
  wire        _GEN_106735 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1756 & _GEN_106501 : _GEN_1083 ? ~_GEN_1756 & _GEN_106501 : ~(_GEN_106849 & _GEN_1756) & _GEN_106501) : _GEN_106501;
  wire        _GEN_106736 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1757 & _GEN_106502 : _GEN_1083 ? ~_GEN_1757 & _GEN_106502 : ~(_GEN_106849 & _GEN_1757) & _GEN_106502) : _GEN_106502;
  wire        _GEN_106737 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1758 & _GEN_106503 : _GEN_1083 ? ~_GEN_1758 & _GEN_106503 : ~(_GEN_106849 & _GEN_1758) & _GEN_106503) : _GEN_106503;
  wire        _GEN_106738 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1759 & _GEN_106504 : _GEN_1083 ? ~_GEN_1759 & _GEN_106504 : ~(_GEN_106849 & _GEN_1759) & _GEN_106504) : _GEN_106504;
  wire        _GEN_106739 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1760 & _GEN_106505 : _GEN_1083 ? ~_GEN_1760 & _GEN_106505 : ~(_GEN_106849 & _GEN_1760) & _GEN_106505) : _GEN_106505;
  wire        _GEN_106740 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1761 & _GEN_106506 : _GEN_1083 ? ~_GEN_1761 & _GEN_106506 : ~(_GEN_106849 & _GEN_1761) & _GEN_106506) : _GEN_106506;
  wire        _GEN_106741 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1762 & _GEN_106507 : _GEN_1083 ? ~_GEN_1762 & _GEN_106507 : ~(_GEN_106849 & _GEN_1762) & _GEN_106507) : _GEN_106507;
  wire        _GEN_106742 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1763 & _GEN_106508 : _GEN_1083 ? ~_GEN_1763 & _GEN_106508 : ~(_GEN_106849 & _GEN_1763) & _GEN_106508) : _GEN_106508;
  wire        _GEN_106743 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1764 & _GEN_106509 : _GEN_1083 ? ~_GEN_1764 & _GEN_106509 : ~(_GEN_106849 & _GEN_1764) & _GEN_106509) : _GEN_106509;
  wire        _GEN_106744 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1765 & _GEN_106510 : _GEN_1083 ? ~_GEN_1765 & _GEN_106510 : ~(_GEN_106849 & _GEN_1765) & _GEN_106510) : _GEN_106510;
  wire        _GEN_106745 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1766 & _GEN_106511 : _GEN_1083 ? ~_GEN_1766 & _GEN_106511 : ~(_GEN_106849 & _GEN_1766) & _GEN_106511) : _GEN_106511;
  wire        _GEN_106746 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1767 & _GEN_106512 : _GEN_1083 ? ~_GEN_1767 & _GEN_106512 : ~(_GEN_106849 & _GEN_1767) & _GEN_106512) : _GEN_106512;
  wire        _GEN_106747 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1768 & _GEN_106513 : _GEN_1083 ? ~_GEN_1768 & _GEN_106513 : ~(_GEN_106849 & _GEN_1768) & _GEN_106513) : _GEN_106513;
  wire        _GEN_106748 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1769 & _GEN_106514 : _GEN_1083 ? ~_GEN_1769 & _GEN_106514 : ~(_GEN_106849 & _GEN_1769) & _GEN_106514) : _GEN_106514;
  wire        _GEN_106749 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1770 & _GEN_106515 : _GEN_1083 ? ~_GEN_1770 & _GEN_106515 : ~(_GEN_106849 & _GEN_1770) & _GEN_106515) : _GEN_106515;
  wire        _GEN_106750 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1771 & _GEN_106516 : _GEN_1083 ? ~_GEN_1771 & _GEN_106516 : ~(_GEN_106849 & _GEN_1771) & _GEN_106516) : _GEN_106516;
  wire        _GEN_106751 = _GEN_1081 ? (_GEN_106684 ? ~_GEN_1772 & _GEN_106517 : _GEN_1083 ? ~_GEN_1772 & _GEN_106517 : ~(_GEN_106849 & _GEN_1772) & _GEN_106517) : _GEN_106517;
  wire        _GEN_106752 = _GEN_1081 ? (_GEN_106684 ? ~(&lcam_ldq_idx_0) & _GEN_106518 : _GEN_1083 ? ~(&lcam_ldq_idx_0) & _GEN_106518 : ~(_GEN_106849 & (&lcam_ldq_idx_0)) & _GEN_106518) : _GEN_106518;
  wire        _GEN_106955 = _GEN_1084 ? (_GEN_106918 ? (|lcam_ldq_idx_1) & _GEN_106721 : _GEN_1086 ? (|lcam_ldq_idx_1) & _GEN_106721 : ~(_GEN_106849 & ~(|lcam_ldq_idx_1)) & _GEN_106721) : _GEN_106721;
  wire        _GEN_106956 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1773 & _GEN_106722 : _GEN_1086 ? ~_GEN_1773 & _GEN_106722 : ~(_GEN_106849 & _GEN_1773) & _GEN_106722) : _GEN_106722;
  wire        _GEN_106957 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1774 & _GEN_106723 : _GEN_1086 ? ~_GEN_1774 & _GEN_106723 : ~(_GEN_106849 & _GEN_1774) & _GEN_106723) : _GEN_106723;
  wire        _GEN_106958 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1775 & _GEN_106724 : _GEN_1086 ? ~_GEN_1775 & _GEN_106724 : ~(_GEN_106849 & _GEN_1775) & _GEN_106724) : _GEN_106724;
  wire        _GEN_106959 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1776 & _GEN_106725 : _GEN_1086 ? ~_GEN_1776 & _GEN_106725 : ~(_GEN_106849 & _GEN_1776) & _GEN_106725) : _GEN_106725;
  wire        _GEN_106960 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1777 & _GEN_106726 : _GEN_1086 ? ~_GEN_1777 & _GEN_106726 : ~(_GEN_106849 & _GEN_1777) & _GEN_106726) : _GEN_106726;
  wire        _GEN_106961 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1778 & _GEN_106727 : _GEN_1086 ? ~_GEN_1778 & _GEN_106727 : ~(_GEN_106849 & _GEN_1778) & _GEN_106727) : _GEN_106727;
  wire        _GEN_106962 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1779 & _GEN_106728 : _GEN_1086 ? ~_GEN_1779 & _GEN_106728 : ~(_GEN_106849 & _GEN_1779) & _GEN_106728) : _GEN_106728;
  wire        _GEN_106963 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1780 & _GEN_106729 : _GEN_1086 ? ~_GEN_1780 & _GEN_106729 : ~(_GEN_106849 & _GEN_1780) & _GEN_106729) : _GEN_106729;
  wire        _GEN_106964 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1781 & _GEN_106730 : _GEN_1086 ? ~_GEN_1781 & _GEN_106730 : ~(_GEN_106849 & _GEN_1781) & _GEN_106730) : _GEN_106730;
  wire        _GEN_106965 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1782 & _GEN_106731 : _GEN_1086 ? ~_GEN_1782 & _GEN_106731 : ~(_GEN_106849 & _GEN_1782) & _GEN_106731) : _GEN_106731;
  wire        _GEN_106966 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1783 & _GEN_106732 : _GEN_1086 ? ~_GEN_1783 & _GEN_106732 : ~(_GEN_106849 & _GEN_1783) & _GEN_106732) : _GEN_106732;
  wire        _GEN_106967 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1784 & _GEN_106733 : _GEN_1086 ? ~_GEN_1784 & _GEN_106733 : ~(_GEN_106849 & _GEN_1784) & _GEN_106733) : _GEN_106733;
  wire        _GEN_106968 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1785 & _GEN_106734 : _GEN_1086 ? ~_GEN_1785 & _GEN_106734 : ~(_GEN_106849 & _GEN_1785) & _GEN_106734) : _GEN_106734;
  wire        _GEN_106969 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1786 & _GEN_106735 : _GEN_1086 ? ~_GEN_1786 & _GEN_106735 : ~(_GEN_106849 & _GEN_1786) & _GEN_106735) : _GEN_106735;
  wire        _GEN_106970 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1787 & _GEN_106736 : _GEN_1086 ? ~_GEN_1787 & _GEN_106736 : ~(_GEN_106849 & _GEN_1787) & _GEN_106736) : _GEN_106736;
  wire        _GEN_106971 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1788 & _GEN_106737 : _GEN_1086 ? ~_GEN_1788 & _GEN_106737 : ~(_GEN_106849 & _GEN_1788) & _GEN_106737) : _GEN_106737;
  wire        _GEN_106972 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1789 & _GEN_106738 : _GEN_1086 ? ~_GEN_1789 & _GEN_106738 : ~(_GEN_106849 & _GEN_1789) & _GEN_106738) : _GEN_106738;
  wire        _GEN_106973 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1790 & _GEN_106739 : _GEN_1086 ? ~_GEN_1790 & _GEN_106739 : ~(_GEN_106849 & _GEN_1790) & _GEN_106739) : _GEN_106739;
  wire        _GEN_106974 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1791 & _GEN_106740 : _GEN_1086 ? ~_GEN_1791 & _GEN_106740 : ~(_GEN_106849 & _GEN_1791) & _GEN_106740) : _GEN_106740;
  wire        _GEN_106975 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1792 & _GEN_106741 : _GEN_1086 ? ~_GEN_1792 & _GEN_106741 : ~(_GEN_106849 & _GEN_1792) & _GEN_106741) : _GEN_106741;
  wire        _GEN_106976 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1793 & _GEN_106742 : _GEN_1086 ? ~_GEN_1793 & _GEN_106742 : ~(_GEN_106849 & _GEN_1793) & _GEN_106742) : _GEN_106742;
  wire        _GEN_106977 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1794 & _GEN_106743 : _GEN_1086 ? ~_GEN_1794 & _GEN_106743 : ~(_GEN_106849 & _GEN_1794) & _GEN_106743) : _GEN_106743;
  wire        _GEN_106978 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1795 & _GEN_106744 : _GEN_1086 ? ~_GEN_1795 & _GEN_106744 : ~(_GEN_106849 & _GEN_1795) & _GEN_106744) : _GEN_106744;
  wire        _GEN_106979 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1796 & _GEN_106745 : _GEN_1086 ? ~_GEN_1796 & _GEN_106745 : ~(_GEN_106849 & _GEN_1796) & _GEN_106745) : _GEN_106745;
  wire        _GEN_106980 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1797 & _GEN_106746 : _GEN_1086 ? ~_GEN_1797 & _GEN_106746 : ~(_GEN_106849 & _GEN_1797) & _GEN_106746) : _GEN_106746;
  wire        _GEN_106981 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1798 & _GEN_106747 : _GEN_1086 ? ~_GEN_1798 & _GEN_106747 : ~(_GEN_106849 & _GEN_1798) & _GEN_106747) : _GEN_106747;
  wire        _GEN_106982 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1799 & _GEN_106748 : _GEN_1086 ? ~_GEN_1799 & _GEN_106748 : ~(_GEN_106849 & _GEN_1799) & _GEN_106748) : _GEN_106748;
  wire        _GEN_106983 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1800 & _GEN_106749 : _GEN_1086 ? ~_GEN_1800 & _GEN_106749 : ~(_GEN_106849 & _GEN_1800) & _GEN_106749) : _GEN_106749;
  wire        _GEN_106984 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1801 & _GEN_106750 : _GEN_1086 ? ~_GEN_1801 & _GEN_106750 : ~(_GEN_106849 & _GEN_1801) & _GEN_106750) : _GEN_106750;
  wire        _GEN_106985 = _GEN_1084 ? (_GEN_106918 ? ~_GEN_1802 & _GEN_106751 : _GEN_1086 ? ~_GEN_1802 & _GEN_106751 : ~(_GEN_106849 & _GEN_1802) & _GEN_106751) : _GEN_106751;
  wire        _GEN_106986 = _GEN_1084 ? (_GEN_106918 ? ~(&lcam_ldq_idx_1) & _GEN_106752 : _GEN_1086 ? ~(&lcam_ldq_idx_1) & _GEN_106752 : ~(_GEN_106849 & (&lcam_ldq_idx_1)) & _GEN_106752) : _GEN_106752;
  wire        _GEN_107189 = _GEN_1087 ? (_GEN_107152 ? (|lcam_ldq_idx_0) & _GEN_106955 : _GEN_1089 ? (|lcam_ldq_idx_0) & _GEN_106955 : ~(_GEN_107317 & ~(|lcam_ldq_idx_0)) & _GEN_106955) : _GEN_106955;
  wire        _GEN_107190 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1743 & _GEN_106956 : _GEN_1089 ? ~_GEN_1743 & _GEN_106956 : ~(_GEN_107317 & _GEN_1743) & _GEN_106956) : _GEN_106956;
  wire        _GEN_107191 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1744 & _GEN_106957 : _GEN_1089 ? ~_GEN_1744 & _GEN_106957 : ~(_GEN_107317 & _GEN_1744) & _GEN_106957) : _GEN_106957;
  wire        _GEN_107192 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1745 & _GEN_106958 : _GEN_1089 ? ~_GEN_1745 & _GEN_106958 : ~(_GEN_107317 & _GEN_1745) & _GEN_106958) : _GEN_106958;
  wire        _GEN_107193 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1746 & _GEN_106959 : _GEN_1089 ? ~_GEN_1746 & _GEN_106959 : ~(_GEN_107317 & _GEN_1746) & _GEN_106959) : _GEN_106959;
  wire        _GEN_107194 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1747 & _GEN_106960 : _GEN_1089 ? ~_GEN_1747 & _GEN_106960 : ~(_GEN_107317 & _GEN_1747) & _GEN_106960) : _GEN_106960;
  wire        _GEN_107195 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1748 & _GEN_106961 : _GEN_1089 ? ~_GEN_1748 & _GEN_106961 : ~(_GEN_107317 & _GEN_1748) & _GEN_106961) : _GEN_106961;
  wire        _GEN_107196 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1749 & _GEN_106962 : _GEN_1089 ? ~_GEN_1749 & _GEN_106962 : ~(_GEN_107317 & _GEN_1749) & _GEN_106962) : _GEN_106962;
  wire        _GEN_107197 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1750 & _GEN_106963 : _GEN_1089 ? ~_GEN_1750 & _GEN_106963 : ~(_GEN_107317 & _GEN_1750) & _GEN_106963) : _GEN_106963;
  wire        _GEN_107198 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1751 & _GEN_106964 : _GEN_1089 ? ~_GEN_1751 & _GEN_106964 : ~(_GEN_107317 & _GEN_1751) & _GEN_106964) : _GEN_106964;
  wire        _GEN_107199 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1752 & _GEN_106965 : _GEN_1089 ? ~_GEN_1752 & _GEN_106965 : ~(_GEN_107317 & _GEN_1752) & _GEN_106965) : _GEN_106965;
  wire        _GEN_107200 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1753 & _GEN_106966 : _GEN_1089 ? ~_GEN_1753 & _GEN_106966 : ~(_GEN_107317 & _GEN_1753) & _GEN_106966) : _GEN_106966;
  wire        _GEN_107201 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1754 & _GEN_106967 : _GEN_1089 ? ~_GEN_1754 & _GEN_106967 : ~(_GEN_107317 & _GEN_1754) & _GEN_106967) : _GEN_106967;
  wire        _GEN_107202 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1755 & _GEN_106968 : _GEN_1089 ? ~_GEN_1755 & _GEN_106968 : ~(_GEN_107317 & _GEN_1755) & _GEN_106968) : _GEN_106968;
  wire        _GEN_107203 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1756 & _GEN_106969 : _GEN_1089 ? ~_GEN_1756 & _GEN_106969 : ~(_GEN_107317 & _GEN_1756) & _GEN_106969) : _GEN_106969;
  wire        _GEN_107204 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1757 & _GEN_106970 : _GEN_1089 ? ~_GEN_1757 & _GEN_106970 : ~(_GEN_107317 & _GEN_1757) & _GEN_106970) : _GEN_106970;
  wire        _GEN_107205 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1758 & _GEN_106971 : _GEN_1089 ? ~_GEN_1758 & _GEN_106971 : ~(_GEN_107317 & _GEN_1758) & _GEN_106971) : _GEN_106971;
  wire        _GEN_107206 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1759 & _GEN_106972 : _GEN_1089 ? ~_GEN_1759 & _GEN_106972 : ~(_GEN_107317 & _GEN_1759) & _GEN_106972) : _GEN_106972;
  wire        _GEN_107207 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1760 & _GEN_106973 : _GEN_1089 ? ~_GEN_1760 & _GEN_106973 : ~(_GEN_107317 & _GEN_1760) & _GEN_106973) : _GEN_106973;
  wire        _GEN_107208 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1761 & _GEN_106974 : _GEN_1089 ? ~_GEN_1761 & _GEN_106974 : ~(_GEN_107317 & _GEN_1761) & _GEN_106974) : _GEN_106974;
  wire        _GEN_107209 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1762 & _GEN_106975 : _GEN_1089 ? ~_GEN_1762 & _GEN_106975 : ~(_GEN_107317 & _GEN_1762) & _GEN_106975) : _GEN_106975;
  wire        _GEN_107210 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1763 & _GEN_106976 : _GEN_1089 ? ~_GEN_1763 & _GEN_106976 : ~(_GEN_107317 & _GEN_1763) & _GEN_106976) : _GEN_106976;
  wire        _GEN_107211 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1764 & _GEN_106977 : _GEN_1089 ? ~_GEN_1764 & _GEN_106977 : ~(_GEN_107317 & _GEN_1764) & _GEN_106977) : _GEN_106977;
  wire        _GEN_107212 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1765 & _GEN_106978 : _GEN_1089 ? ~_GEN_1765 & _GEN_106978 : ~(_GEN_107317 & _GEN_1765) & _GEN_106978) : _GEN_106978;
  wire        _GEN_107213 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1766 & _GEN_106979 : _GEN_1089 ? ~_GEN_1766 & _GEN_106979 : ~(_GEN_107317 & _GEN_1766) & _GEN_106979) : _GEN_106979;
  wire        _GEN_107214 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1767 & _GEN_106980 : _GEN_1089 ? ~_GEN_1767 & _GEN_106980 : ~(_GEN_107317 & _GEN_1767) & _GEN_106980) : _GEN_106980;
  wire        _GEN_107215 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1768 & _GEN_106981 : _GEN_1089 ? ~_GEN_1768 & _GEN_106981 : ~(_GEN_107317 & _GEN_1768) & _GEN_106981) : _GEN_106981;
  wire        _GEN_107216 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1769 & _GEN_106982 : _GEN_1089 ? ~_GEN_1769 & _GEN_106982 : ~(_GEN_107317 & _GEN_1769) & _GEN_106982) : _GEN_106982;
  wire        _GEN_107217 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1770 & _GEN_106983 : _GEN_1089 ? ~_GEN_1770 & _GEN_106983 : ~(_GEN_107317 & _GEN_1770) & _GEN_106983) : _GEN_106983;
  wire        _GEN_107218 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1771 & _GEN_106984 : _GEN_1089 ? ~_GEN_1771 & _GEN_106984 : ~(_GEN_107317 & _GEN_1771) & _GEN_106984) : _GEN_106984;
  wire        _GEN_107219 = _GEN_1087 ? (_GEN_107152 ? ~_GEN_1772 & _GEN_106985 : _GEN_1089 ? ~_GEN_1772 & _GEN_106985 : ~(_GEN_107317 & _GEN_1772) & _GEN_106985) : _GEN_106985;
  wire        _GEN_107220 = _GEN_1087 ? (_GEN_107152 ? ~(&lcam_ldq_idx_0) & _GEN_106986 : _GEN_1089 ? ~(&lcam_ldq_idx_0) & _GEN_106986 : ~(_GEN_107317 & (&lcam_ldq_idx_0)) & _GEN_106986) : _GEN_106986;
  wire        _GEN_107423 = _GEN_1090 ? (_GEN_107386 ? (|lcam_ldq_idx_1) & _GEN_107189 : _GEN_1092 ? (|lcam_ldq_idx_1) & _GEN_107189 : ~(_GEN_107317 & ~(|lcam_ldq_idx_1)) & _GEN_107189) : _GEN_107189;
  wire        _GEN_107424 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1773 & _GEN_107190 : _GEN_1092 ? ~_GEN_1773 & _GEN_107190 : ~(_GEN_107317 & _GEN_1773) & _GEN_107190) : _GEN_107190;
  wire        _GEN_107425 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1774 & _GEN_107191 : _GEN_1092 ? ~_GEN_1774 & _GEN_107191 : ~(_GEN_107317 & _GEN_1774) & _GEN_107191) : _GEN_107191;
  wire        _GEN_107426 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1775 & _GEN_107192 : _GEN_1092 ? ~_GEN_1775 & _GEN_107192 : ~(_GEN_107317 & _GEN_1775) & _GEN_107192) : _GEN_107192;
  wire        _GEN_107427 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1776 & _GEN_107193 : _GEN_1092 ? ~_GEN_1776 & _GEN_107193 : ~(_GEN_107317 & _GEN_1776) & _GEN_107193) : _GEN_107193;
  wire        _GEN_107428 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1777 & _GEN_107194 : _GEN_1092 ? ~_GEN_1777 & _GEN_107194 : ~(_GEN_107317 & _GEN_1777) & _GEN_107194) : _GEN_107194;
  wire        _GEN_107429 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1778 & _GEN_107195 : _GEN_1092 ? ~_GEN_1778 & _GEN_107195 : ~(_GEN_107317 & _GEN_1778) & _GEN_107195) : _GEN_107195;
  wire        _GEN_107430 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1779 & _GEN_107196 : _GEN_1092 ? ~_GEN_1779 & _GEN_107196 : ~(_GEN_107317 & _GEN_1779) & _GEN_107196) : _GEN_107196;
  wire        _GEN_107431 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1780 & _GEN_107197 : _GEN_1092 ? ~_GEN_1780 & _GEN_107197 : ~(_GEN_107317 & _GEN_1780) & _GEN_107197) : _GEN_107197;
  wire        _GEN_107432 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1781 & _GEN_107198 : _GEN_1092 ? ~_GEN_1781 & _GEN_107198 : ~(_GEN_107317 & _GEN_1781) & _GEN_107198) : _GEN_107198;
  wire        _GEN_107433 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1782 & _GEN_107199 : _GEN_1092 ? ~_GEN_1782 & _GEN_107199 : ~(_GEN_107317 & _GEN_1782) & _GEN_107199) : _GEN_107199;
  wire        _GEN_107434 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1783 & _GEN_107200 : _GEN_1092 ? ~_GEN_1783 & _GEN_107200 : ~(_GEN_107317 & _GEN_1783) & _GEN_107200) : _GEN_107200;
  wire        _GEN_107435 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1784 & _GEN_107201 : _GEN_1092 ? ~_GEN_1784 & _GEN_107201 : ~(_GEN_107317 & _GEN_1784) & _GEN_107201) : _GEN_107201;
  wire        _GEN_107436 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1785 & _GEN_107202 : _GEN_1092 ? ~_GEN_1785 & _GEN_107202 : ~(_GEN_107317 & _GEN_1785) & _GEN_107202) : _GEN_107202;
  wire        _GEN_107437 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1786 & _GEN_107203 : _GEN_1092 ? ~_GEN_1786 & _GEN_107203 : ~(_GEN_107317 & _GEN_1786) & _GEN_107203) : _GEN_107203;
  wire        _GEN_107438 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1787 & _GEN_107204 : _GEN_1092 ? ~_GEN_1787 & _GEN_107204 : ~(_GEN_107317 & _GEN_1787) & _GEN_107204) : _GEN_107204;
  wire        _GEN_107439 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1788 & _GEN_107205 : _GEN_1092 ? ~_GEN_1788 & _GEN_107205 : ~(_GEN_107317 & _GEN_1788) & _GEN_107205) : _GEN_107205;
  wire        _GEN_107440 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1789 & _GEN_107206 : _GEN_1092 ? ~_GEN_1789 & _GEN_107206 : ~(_GEN_107317 & _GEN_1789) & _GEN_107206) : _GEN_107206;
  wire        _GEN_107441 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1790 & _GEN_107207 : _GEN_1092 ? ~_GEN_1790 & _GEN_107207 : ~(_GEN_107317 & _GEN_1790) & _GEN_107207) : _GEN_107207;
  wire        _GEN_107442 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1791 & _GEN_107208 : _GEN_1092 ? ~_GEN_1791 & _GEN_107208 : ~(_GEN_107317 & _GEN_1791) & _GEN_107208) : _GEN_107208;
  wire        _GEN_107443 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1792 & _GEN_107209 : _GEN_1092 ? ~_GEN_1792 & _GEN_107209 : ~(_GEN_107317 & _GEN_1792) & _GEN_107209) : _GEN_107209;
  wire        _GEN_107444 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1793 & _GEN_107210 : _GEN_1092 ? ~_GEN_1793 & _GEN_107210 : ~(_GEN_107317 & _GEN_1793) & _GEN_107210) : _GEN_107210;
  wire        _GEN_107445 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1794 & _GEN_107211 : _GEN_1092 ? ~_GEN_1794 & _GEN_107211 : ~(_GEN_107317 & _GEN_1794) & _GEN_107211) : _GEN_107211;
  wire        _GEN_107446 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1795 & _GEN_107212 : _GEN_1092 ? ~_GEN_1795 & _GEN_107212 : ~(_GEN_107317 & _GEN_1795) & _GEN_107212) : _GEN_107212;
  wire        _GEN_107447 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1796 & _GEN_107213 : _GEN_1092 ? ~_GEN_1796 & _GEN_107213 : ~(_GEN_107317 & _GEN_1796) & _GEN_107213) : _GEN_107213;
  wire        _GEN_107448 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1797 & _GEN_107214 : _GEN_1092 ? ~_GEN_1797 & _GEN_107214 : ~(_GEN_107317 & _GEN_1797) & _GEN_107214) : _GEN_107214;
  wire        _GEN_107449 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1798 & _GEN_107215 : _GEN_1092 ? ~_GEN_1798 & _GEN_107215 : ~(_GEN_107317 & _GEN_1798) & _GEN_107215) : _GEN_107215;
  wire        _GEN_107450 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1799 & _GEN_107216 : _GEN_1092 ? ~_GEN_1799 & _GEN_107216 : ~(_GEN_107317 & _GEN_1799) & _GEN_107216) : _GEN_107216;
  wire        _GEN_107451 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1800 & _GEN_107217 : _GEN_1092 ? ~_GEN_1800 & _GEN_107217 : ~(_GEN_107317 & _GEN_1800) & _GEN_107217) : _GEN_107217;
  wire        _GEN_107452 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1801 & _GEN_107218 : _GEN_1092 ? ~_GEN_1801 & _GEN_107218 : ~(_GEN_107317 & _GEN_1801) & _GEN_107218) : _GEN_107218;
  wire        _GEN_107453 = _GEN_1090 ? (_GEN_107386 ? ~_GEN_1802 & _GEN_107219 : _GEN_1092 ? ~_GEN_1802 & _GEN_107219 : ~(_GEN_107317 & _GEN_1802) & _GEN_107219) : _GEN_107219;
  wire        _GEN_107454 = _GEN_1090 ? (_GEN_107386 ? ~(&lcam_ldq_idx_1) & _GEN_107220 : _GEN_1092 ? ~(&lcam_ldq_idx_1) & _GEN_107220 : ~(_GEN_107317 & (&lcam_ldq_idx_1)) & _GEN_107220) : _GEN_107220;
  wire        _GEN_107657 = _GEN_1093 ? (_GEN_107620 ? (|lcam_ldq_idx_0) & _GEN_107423 : _GEN_1095 ? (|lcam_ldq_idx_0) & _GEN_107423 : ~(_GEN_107785 & ~(|lcam_ldq_idx_0)) & _GEN_107423) : _GEN_107423;
  wire        _GEN_107658 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1743 & _GEN_107424 : _GEN_1095 ? ~_GEN_1743 & _GEN_107424 : ~(_GEN_107785 & _GEN_1743) & _GEN_107424) : _GEN_107424;
  wire        _GEN_107659 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1744 & _GEN_107425 : _GEN_1095 ? ~_GEN_1744 & _GEN_107425 : ~(_GEN_107785 & _GEN_1744) & _GEN_107425) : _GEN_107425;
  wire        _GEN_107660 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1745 & _GEN_107426 : _GEN_1095 ? ~_GEN_1745 & _GEN_107426 : ~(_GEN_107785 & _GEN_1745) & _GEN_107426) : _GEN_107426;
  wire        _GEN_107661 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1746 & _GEN_107427 : _GEN_1095 ? ~_GEN_1746 & _GEN_107427 : ~(_GEN_107785 & _GEN_1746) & _GEN_107427) : _GEN_107427;
  wire        _GEN_107662 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1747 & _GEN_107428 : _GEN_1095 ? ~_GEN_1747 & _GEN_107428 : ~(_GEN_107785 & _GEN_1747) & _GEN_107428) : _GEN_107428;
  wire        _GEN_107663 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1748 & _GEN_107429 : _GEN_1095 ? ~_GEN_1748 & _GEN_107429 : ~(_GEN_107785 & _GEN_1748) & _GEN_107429) : _GEN_107429;
  wire        _GEN_107664 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1749 & _GEN_107430 : _GEN_1095 ? ~_GEN_1749 & _GEN_107430 : ~(_GEN_107785 & _GEN_1749) & _GEN_107430) : _GEN_107430;
  wire        _GEN_107665 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1750 & _GEN_107431 : _GEN_1095 ? ~_GEN_1750 & _GEN_107431 : ~(_GEN_107785 & _GEN_1750) & _GEN_107431) : _GEN_107431;
  wire        _GEN_107666 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1751 & _GEN_107432 : _GEN_1095 ? ~_GEN_1751 & _GEN_107432 : ~(_GEN_107785 & _GEN_1751) & _GEN_107432) : _GEN_107432;
  wire        _GEN_107667 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1752 & _GEN_107433 : _GEN_1095 ? ~_GEN_1752 & _GEN_107433 : ~(_GEN_107785 & _GEN_1752) & _GEN_107433) : _GEN_107433;
  wire        _GEN_107668 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1753 & _GEN_107434 : _GEN_1095 ? ~_GEN_1753 & _GEN_107434 : ~(_GEN_107785 & _GEN_1753) & _GEN_107434) : _GEN_107434;
  wire        _GEN_107669 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1754 & _GEN_107435 : _GEN_1095 ? ~_GEN_1754 & _GEN_107435 : ~(_GEN_107785 & _GEN_1754) & _GEN_107435) : _GEN_107435;
  wire        _GEN_107670 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1755 & _GEN_107436 : _GEN_1095 ? ~_GEN_1755 & _GEN_107436 : ~(_GEN_107785 & _GEN_1755) & _GEN_107436) : _GEN_107436;
  wire        _GEN_107671 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1756 & _GEN_107437 : _GEN_1095 ? ~_GEN_1756 & _GEN_107437 : ~(_GEN_107785 & _GEN_1756) & _GEN_107437) : _GEN_107437;
  wire        _GEN_107672 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1757 & _GEN_107438 : _GEN_1095 ? ~_GEN_1757 & _GEN_107438 : ~(_GEN_107785 & _GEN_1757) & _GEN_107438) : _GEN_107438;
  wire        _GEN_107673 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1758 & _GEN_107439 : _GEN_1095 ? ~_GEN_1758 & _GEN_107439 : ~(_GEN_107785 & _GEN_1758) & _GEN_107439) : _GEN_107439;
  wire        _GEN_107674 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1759 & _GEN_107440 : _GEN_1095 ? ~_GEN_1759 & _GEN_107440 : ~(_GEN_107785 & _GEN_1759) & _GEN_107440) : _GEN_107440;
  wire        _GEN_107675 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1760 & _GEN_107441 : _GEN_1095 ? ~_GEN_1760 & _GEN_107441 : ~(_GEN_107785 & _GEN_1760) & _GEN_107441) : _GEN_107441;
  wire        _GEN_107676 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1761 & _GEN_107442 : _GEN_1095 ? ~_GEN_1761 & _GEN_107442 : ~(_GEN_107785 & _GEN_1761) & _GEN_107442) : _GEN_107442;
  wire        _GEN_107677 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1762 & _GEN_107443 : _GEN_1095 ? ~_GEN_1762 & _GEN_107443 : ~(_GEN_107785 & _GEN_1762) & _GEN_107443) : _GEN_107443;
  wire        _GEN_107678 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1763 & _GEN_107444 : _GEN_1095 ? ~_GEN_1763 & _GEN_107444 : ~(_GEN_107785 & _GEN_1763) & _GEN_107444) : _GEN_107444;
  wire        _GEN_107679 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1764 & _GEN_107445 : _GEN_1095 ? ~_GEN_1764 & _GEN_107445 : ~(_GEN_107785 & _GEN_1764) & _GEN_107445) : _GEN_107445;
  wire        _GEN_107680 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1765 & _GEN_107446 : _GEN_1095 ? ~_GEN_1765 & _GEN_107446 : ~(_GEN_107785 & _GEN_1765) & _GEN_107446) : _GEN_107446;
  wire        _GEN_107681 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1766 & _GEN_107447 : _GEN_1095 ? ~_GEN_1766 & _GEN_107447 : ~(_GEN_107785 & _GEN_1766) & _GEN_107447) : _GEN_107447;
  wire        _GEN_107682 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1767 & _GEN_107448 : _GEN_1095 ? ~_GEN_1767 & _GEN_107448 : ~(_GEN_107785 & _GEN_1767) & _GEN_107448) : _GEN_107448;
  wire        _GEN_107683 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1768 & _GEN_107449 : _GEN_1095 ? ~_GEN_1768 & _GEN_107449 : ~(_GEN_107785 & _GEN_1768) & _GEN_107449) : _GEN_107449;
  wire        _GEN_107684 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1769 & _GEN_107450 : _GEN_1095 ? ~_GEN_1769 & _GEN_107450 : ~(_GEN_107785 & _GEN_1769) & _GEN_107450) : _GEN_107450;
  wire        _GEN_107685 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1770 & _GEN_107451 : _GEN_1095 ? ~_GEN_1770 & _GEN_107451 : ~(_GEN_107785 & _GEN_1770) & _GEN_107451) : _GEN_107451;
  wire        _GEN_107686 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1771 & _GEN_107452 : _GEN_1095 ? ~_GEN_1771 & _GEN_107452 : ~(_GEN_107785 & _GEN_1771) & _GEN_107452) : _GEN_107452;
  wire        _GEN_107687 = _GEN_1093 ? (_GEN_107620 ? ~_GEN_1772 & _GEN_107453 : _GEN_1095 ? ~_GEN_1772 & _GEN_107453 : ~(_GEN_107785 & _GEN_1772) & _GEN_107453) : _GEN_107453;
  wire        _GEN_107688 = _GEN_1093 ? (_GEN_107620 ? ~(&lcam_ldq_idx_0) & _GEN_107454 : _GEN_1095 ? ~(&lcam_ldq_idx_0) & _GEN_107454 : ~(_GEN_107785 & (&lcam_ldq_idx_0)) & _GEN_107454) : _GEN_107454;
  wire        _GEN_107891 = _GEN_1096 ? (_GEN_107854 ? (|lcam_ldq_idx_1) & _GEN_107657 : _GEN_1098 ? (|lcam_ldq_idx_1) & _GEN_107657 : ~(_GEN_107785 & ~(|lcam_ldq_idx_1)) & _GEN_107657) : _GEN_107657;
  wire        _GEN_107892 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1773 & _GEN_107658 : _GEN_1098 ? ~_GEN_1773 & _GEN_107658 : ~(_GEN_107785 & _GEN_1773) & _GEN_107658) : _GEN_107658;
  wire        _GEN_107893 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1774 & _GEN_107659 : _GEN_1098 ? ~_GEN_1774 & _GEN_107659 : ~(_GEN_107785 & _GEN_1774) & _GEN_107659) : _GEN_107659;
  wire        _GEN_107894 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1775 & _GEN_107660 : _GEN_1098 ? ~_GEN_1775 & _GEN_107660 : ~(_GEN_107785 & _GEN_1775) & _GEN_107660) : _GEN_107660;
  wire        _GEN_107895 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1776 & _GEN_107661 : _GEN_1098 ? ~_GEN_1776 & _GEN_107661 : ~(_GEN_107785 & _GEN_1776) & _GEN_107661) : _GEN_107661;
  wire        _GEN_107896 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1777 & _GEN_107662 : _GEN_1098 ? ~_GEN_1777 & _GEN_107662 : ~(_GEN_107785 & _GEN_1777) & _GEN_107662) : _GEN_107662;
  wire        _GEN_107897 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1778 & _GEN_107663 : _GEN_1098 ? ~_GEN_1778 & _GEN_107663 : ~(_GEN_107785 & _GEN_1778) & _GEN_107663) : _GEN_107663;
  wire        _GEN_107898 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1779 & _GEN_107664 : _GEN_1098 ? ~_GEN_1779 & _GEN_107664 : ~(_GEN_107785 & _GEN_1779) & _GEN_107664) : _GEN_107664;
  wire        _GEN_107899 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1780 & _GEN_107665 : _GEN_1098 ? ~_GEN_1780 & _GEN_107665 : ~(_GEN_107785 & _GEN_1780) & _GEN_107665) : _GEN_107665;
  wire        _GEN_107900 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1781 & _GEN_107666 : _GEN_1098 ? ~_GEN_1781 & _GEN_107666 : ~(_GEN_107785 & _GEN_1781) & _GEN_107666) : _GEN_107666;
  wire        _GEN_107901 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1782 & _GEN_107667 : _GEN_1098 ? ~_GEN_1782 & _GEN_107667 : ~(_GEN_107785 & _GEN_1782) & _GEN_107667) : _GEN_107667;
  wire        _GEN_107902 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1783 & _GEN_107668 : _GEN_1098 ? ~_GEN_1783 & _GEN_107668 : ~(_GEN_107785 & _GEN_1783) & _GEN_107668) : _GEN_107668;
  wire        _GEN_107903 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1784 & _GEN_107669 : _GEN_1098 ? ~_GEN_1784 & _GEN_107669 : ~(_GEN_107785 & _GEN_1784) & _GEN_107669) : _GEN_107669;
  wire        _GEN_107904 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1785 & _GEN_107670 : _GEN_1098 ? ~_GEN_1785 & _GEN_107670 : ~(_GEN_107785 & _GEN_1785) & _GEN_107670) : _GEN_107670;
  wire        _GEN_107905 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1786 & _GEN_107671 : _GEN_1098 ? ~_GEN_1786 & _GEN_107671 : ~(_GEN_107785 & _GEN_1786) & _GEN_107671) : _GEN_107671;
  wire        _GEN_107906 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1787 & _GEN_107672 : _GEN_1098 ? ~_GEN_1787 & _GEN_107672 : ~(_GEN_107785 & _GEN_1787) & _GEN_107672) : _GEN_107672;
  wire        _GEN_107907 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1788 & _GEN_107673 : _GEN_1098 ? ~_GEN_1788 & _GEN_107673 : ~(_GEN_107785 & _GEN_1788) & _GEN_107673) : _GEN_107673;
  wire        _GEN_107908 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1789 & _GEN_107674 : _GEN_1098 ? ~_GEN_1789 & _GEN_107674 : ~(_GEN_107785 & _GEN_1789) & _GEN_107674) : _GEN_107674;
  wire        _GEN_107909 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1790 & _GEN_107675 : _GEN_1098 ? ~_GEN_1790 & _GEN_107675 : ~(_GEN_107785 & _GEN_1790) & _GEN_107675) : _GEN_107675;
  wire        _GEN_107910 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1791 & _GEN_107676 : _GEN_1098 ? ~_GEN_1791 & _GEN_107676 : ~(_GEN_107785 & _GEN_1791) & _GEN_107676) : _GEN_107676;
  wire        _GEN_107911 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1792 & _GEN_107677 : _GEN_1098 ? ~_GEN_1792 & _GEN_107677 : ~(_GEN_107785 & _GEN_1792) & _GEN_107677) : _GEN_107677;
  wire        _GEN_107912 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1793 & _GEN_107678 : _GEN_1098 ? ~_GEN_1793 & _GEN_107678 : ~(_GEN_107785 & _GEN_1793) & _GEN_107678) : _GEN_107678;
  wire        _GEN_107913 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1794 & _GEN_107679 : _GEN_1098 ? ~_GEN_1794 & _GEN_107679 : ~(_GEN_107785 & _GEN_1794) & _GEN_107679) : _GEN_107679;
  wire        _GEN_107914 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1795 & _GEN_107680 : _GEN_1098 ? ~_GEN_1795 & _GEN_107680 : ~(_GEN_107785 & _GEN_1795) & _GEN_107680) : _GEN_107680;
  wire        _GEN_107915 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1796 & _GEN_107681 : _GEN_1098 ? ~_GEN_1796 & _GEN_107681 : ~(_GEN_107785 & _GEN_1796) & _GEN_107681) : _GEN_107681;
  wire        _GEN_107916 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1797 & _GEN_107682 : _GEN_1098 ? ~_GEN_1797 & _GEN_107682 : ~(_GEN_107785 & _GEN_1797) & _GEN_107682) : _GEN_107682;
  wire        _GEN_107917 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1798 & _GEN_107683 : _GEN_1098 ? ~_GEN_1798 & _GEN_107683 : ~(_GEN_107785 & _GEN_1798) & _GEN_107683) : _GEN_107683;
  wire        _GEN_107918 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1799 & _GEN_107684 : _GEN_1098 ? ~_GEN_1799 & _GEN_107684 : ~(_GEN_107785 & _GEN_1799) & _GEN_107684) : _GEN_107684;
  wire        _GEN_107919 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1800 & _GEN_107685 : _GEN_1098 ? ~_GEN_1800 & _GEN_107685 : ~(_GEN_107785 & _GEN_1800) & _GEN_107685) : _GEN_107685;
  wire        _GEN_107920 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1801 & _GEN_107686 : _GEN_1098 ? ~_GEN_1801 & _GEN_107686 : ~(_GEN_107785 & _GEN_1801) & _GEN_107686) : _GEN_107686;
  wire        _GEN_107921 = _GEN_1096 ? (_GEN_107854 ? ~_GEN_1802 & _GEN_107687 : _GEN_1098 ? ~_GEN_1802 & _GEN_107687 : ~(_GEN_107785 & _GEN_1802) & _GEN_107687) : _GEN_107687;
  wire        _GEN_107922 = _GEN_1096 ? (_GEN_107854 ? ~(&lcam_ldq_idx_1) & _GEN_107688 : _GEN_1098 ? ~(&lcam_ldq_idx_1) & _GEN_107688 : ~(_GEN_107785 & (&lcam_ldq_idx_1)) & _GEN_107688) : _GEN_107688;
  wire        _GEN_108125 = _GEN_1099 ? (_GEN_108088 ? (|lcam_ldq_idx_0) & _GEN_107891 : _GEN_1101 ? (|lcam_ldq_idx_0) & _GEN_107891 : ~(_GEN_108253 & ~(|lcam_ldq_idx_0)) & _GEN_107891) : _GEN_107891;
  wire        _GEN_108126 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1743 & _GEN_107892 : _GEN_1101 ? ~_GEN_1743 & _GEN_107892 : ~(_GEN_108253 & _GEN_1743) & _GEN_107892) : _GEN_107892;
  wire        _GEN_108127 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1744 & _GEN_107893 : _GEN_1101 ? ~_GEN_1744 & _GEN_107893 : ~(_GEN_108253 & _GEN_1744) & _GEN_107893) : _GEN_107893;
  wire        _GEN_108128 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1745 & _GEN_107894 : _GEN_1101 ? ~_GEN_1745 & _GEN_107894 : ~(_GEN_108253 & _GEN_1745) & _GEN_107894) : _GEN_107894;
  wire        _GEN_108129 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1746 & _GEN_107895 : _GEN_1101 ? ~_GEN_1746 & _GEN_107895 : ~(_GEN_108253 & _GEN_1746) & _GEN_107895) : _GEN_107895;
  wire        _GEN_108130 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1747 & _GEN_107896 : _GEN_1101 ? ~_GEN_1747 & _GEN_107896 : ~(_GEN_108253 & _GEN_1747) & _GEN_107896) : _GEN_107896;
  wire        _GEN_108131 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1748 & _GEN_107897 : _GEN_1101 ? ~_GEN_1748 & _GEN_107897 : ~(_GEN_108253 & _GEN_1748) & _GEN_107897) : _GEN_107897;
  wire        _GEN_108132 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1749 & _GEN_107898 : _GEN_1101 ? ~_GEN_1749 & _GEN_107898 : ~(_GEN_108253 & _GEN_1749) & _GEN_107898) : _GEN_107898;
  wire        _GEN_108133 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1750 & _GEN_107899 : _GEN_1101 ? ~_GEN_1750 & _GEN_107899 : ~(_GEN_108253 & _GEN_1750) & _GEN_107899) : _GEN_107899;
  wire        _GEN_108134 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1751 & _GEN_107900 : _GEN_1101 ? ~_GEN_1751 & _GEN_107900 : ~(_GEN_108253 & _GEN_1751) & _GEN_107900) : _GEN_107900;
  wire        _GEN_108135 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1752 & _GEN_107901 : _GEN_1101 ? ~_GEN_1752 & _GEN_107901 : ~(_GEN_108253 & _GEN_1752) & _GEN_107901) : _GEN_107901;
  wire        _GEN_108136 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1753 & _GEN_107902 : _GEN_1101 ? ~_GEN_1753 & _GEN_107902 : ~(_GEN_108253 & _GEN_1753) & _GEN_107902) : _GEN_107902;
  wire        _GEN_108137 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1754 & _GEN_107903 : _GEN_1101 ? ~_GEN_1754 & _GEN_107903 : ~(_GEN_108253 & _GEN_1754) & _GEN_107903) : _GEN_107903;
  wire        _GEN_108138 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1755 & _GEN_107904 : _GEN_1101 ? ~_GEN_1755 & _GEN_107904 : ~(_GEN_108253 & _GEN_1755) & _GEN_107904) : _GEN_107904;
  wire        _GEN_108139 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1756 & _GEN_107905 : _GEN_1101 ? ~_GEN_1756 & _GEN_107905 : ~(_GEN_108253 & _GEN_1756) & _GEN_107905) : _GEN_107905;
  wire        _GEN_108140 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1757 & _GEN_107906 : _GEN_1101 ? ~_GEN_1757 & _GEN_107906 : ~(_GEN_108253 & _GEN_1757) & _GEN_107906) : _GEN_107906;
  wire        _GEN_108141 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1758 & _GEN_107907 : _GEN_1101 ? ~_GEN_1758 & _GEN_107907 : ~(_GEN_108253 & _GEN_1758) & _GEN_107907) : _GEN_107907;
  wire        _GEN_108142 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1759 & _GEN_107908 : _GEN_1101 ? ~_GEN_1759 & _GEN_107908 : ~(_GEN_108253 & _GEN_1759) & _GEN_107908) : _GEN_107908;
  wire        _GEN_108143 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1760 & _GEN_107909 : _GEN_1101 ? ~_GEN_1760 & _GEN_107909 : ~(_GEN_108253 & _GEN_1760) & _GEN_107909) : _GEN_107909;
  wire        _GEN_108144 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1761 & _GEN_107910 : _GEN_1101 ? ~_GEN_1761 & _GEN_107910 : ~(_GEN_108253 & _GEN_1761) & _GEN_107910) : _GEN_107910;
  wire        _GEN_108145 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1762 & _GEN_107911 : _GEN_1101 ? ~_GEN_1762 & _GEN_107911 : ~(_GEN_108253 & _GEN_1762) & _GEN_107911) : _GEN_107911;
  wire        _GEN_108146 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1763 & _GEN_107912 : _GEN_1101 ? ~_GEN_1763 & _GEN_107912 : ~(_GEN_108253 & _GEN_1763) & _GEN_107912) : _GEN_107912;
  wire        _GEN_108147 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1764 & _GEN_107913 : _GEN_1101 ? ~_GEN_1764 & _GEN_107913 : ~(_GEN_108253 & _GEN_1764) & _GEN_107913) : _GEN_107913;
  wire        _GEN_108148 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1765 & _GEN_107914 : _GEN_1101 ? ~_GEN_1765 & _GEN_107914 : ~(_GEN_108253 & _GEN_1765) & _GEN_107914) : _GEN_107914;
  wire        _GEN_108149 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1766 & _GEN_107915 : _GEN_1101 ? ~_GEN_1766 & _GEN_107915 : ~(_GEN_108253 & _GEN_1766) & _GEN_107915) : _GEN_107915;
  wire        _GEN_108150 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1767 & _GEN_107916 : _GEN_1101 ? ~_GEN_1767 & _GEN_107916 : ~(_GEN_108253 & _GEN_1767) & _GEN_107916) : _GEN_107916;
  wire        _GEN_108151 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1768 & _GEN_107917 : _GEN_1101 ? ~_GEN_1768 & _GEN_107917 : ~(_GEN_108253 & _GEN_1768) & _GEN_107917) : _GEN_107917;
  wire        _GEN_108152 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1769 & _GEN_107918 : _GEN_1101 ? ~_GEN_1769 & _GEN_107918 : ~(_GEN_108253 & _GEN_1769) & _GEN_107918) : _GEN_107918;
  wire        _GEN_108153 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1770 & _GEN_107919 : _GEN_1101 ? ~_GEN_1770 & _GEN_107919 : ~(_GEN_108253 & _GEN_1770) & _GEN_107919) : _GEN_107919;
  wire        _GEN_108154 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1771 & _GEN_107920 : _GEN_1101 ? ~_GEN_1771 & _GEN_107920 : ~(_GEN_108253 & _GEN_1771) & _GEN_107920) : _GEN_107920;
  wire        _GEN_108155 = _GEN_1099 ? (_GEN_108088 ? ~_GEN_1772 & _GEN_107921 : _GEN_1101 ? ~_GEN_1772 & _GEN_107921 : ~(_GEN_108253 & _GEN_1772) & _GEN_107921) : _GEN_107921;
  wire        _GEN_108156 = _GEN_1099 ? (_GEN_108088 ? ~(&lcam_ldq_idx_0) & _GEN_107922 : _GEN_1101 ? ~(&lcam_ldq_idx_0) & _GEN_107922 : ~(_GEN_108253 & (&lcam_ldq_idx_0)) & _GEN_107922) : _GEN_107922;
  wire        _GEN_108359 = _GEN_1102 ? (_GEN_108322 ? (|lcam_ldq_idx_1) & _GEN_108125 : _GEN_1104 ? (|lcam_ldq_idx_1) & _GEN_108125 : ~(_GEN_108253 & ~(|lcam_ldq_idx_1)) & _GEN_108125) : _GEN_108125;
  wire        _GEN_108360 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1773 & _GEN_108126 : _GEN_1104 ? ~_GEN_1773 & _GEN_108126 : ~(_GEN_108253 & _GEN_1773) & _GEN_108126) : _GEN_108126;
  wire        _GEN_108361 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1774 & _GEN_108127 : _GEN_1104 ? ~_GEN_1774 & _GEN_108127 : ~(_GEN_108253 & _GEN_1774) & _GEN_108127) : _GEN_108127;
  wire        _GEN_108362 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1775 & _GEN_108128 : _GEN_1104 ? ~_GEN_1775 & _GEN_108128 : ~(_GEN_108253 & _GEN_1775) & _GEN_108128) : _GEN_108128;
  wire        _GEN_108363 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1776 & _GEN_108129 : _GEN_1104 ? ~_GEN_1776 & _GEN_108129 : ~(_GEN_108253 & _GEN_1776) & _GEN_108129) : _GEN_108129;
  wire        _GEN_108364 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1777 & _GEN_108130 : _GEN_1104 ? ~_GEN_1777 & _GEN_108130 : ~(_GEN_108253 & _GEN_1777) & _GEN_108130) : _GEN_108130;
  wire        _GEN_108365 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1778 & _GEN_108131 : _GEN_1104 ? ~_GEN_1778 & _GEN_108131 : ~(_GEN_108253 & _GEN_1778) & _GEN_108131) : _GEN_108131;
  wire        _GEN_108366 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1779 & _GEN_108132 : _GEN_1104 ? ~_GEN_1779 & _GEN_108132 : ~(_GEN_108253 & _GEN_1779) & _GEN_108132) : _GEN_108132;
  wire        _GEN_108367 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1780 & _GEN_108133 : _GEN_1104 ? ~_GEN_1780 & _GEN_108133 : ~(_GEN_108253 & _GEN_1780) & _GEN_108133) : _GEN_108133;
  wire        _GEN_108368 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1781 & _GEN_108134 : _GEN_1104 ? ~_GEN_1781 & _GEN_108134 : ~(_GEN_108253 & _GEN_1781) & _GEN_108134) : _GEN_108134;
  wire        _GEN_108369 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1782 & _GEN_108135 : _GEN_1104 ? ~_GEN_1782 & _GEN_108135 : ~(_GEN_108253 & _GEN_1782) & _GEN_108135) : _GEN_108135;
  wire        _GEN_108370 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1783 & _GEN_108136 : _GEN_1104 ? ~_GEN_1783 & _GEN_108136 : ~(_GEN_108253 & _GEN_1783) & _GEN_108136) : _GEN_108136;
  wire        _GEN_108371 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1784 & _GEN_108137 : _GEN_1104 ? ~_GEN_1784 & _GEN_108137 : ~(_GEN_108253 & _GEN_1784) & _GEN_108137) : _GEN_108137;
  wire        _GEN_108372 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1785 & _GEN_108138 : _GEN_1104 ? ~_GEN_1785 & _GEN_108138 : ~(_GEN_108253 & _GEN_1785) & _GEN_108138) : _GEN_108138;
  wire        _GEN_108373 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1786 & _GEN_108139 : _GEN_1104 ? ~_GEN_1786 & _GEN_108139 : ~(_GEN_108253 & _GEN_1786) & _GEN_108139) : _GEN_108139;
  wire        _GEN_108374 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1787 & _GEN_108140 : _GEN_1104 ? ~_GEN_1787 & _GEN_108140 : ~(_GEN_108253 & _GEN_1787) & _GEN_108140) : _GEN_108140;
  wire        _GEN_108375 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1788 & _GEN_108141 : _GEN_1104 ? ~_GEN_1788 & _GEN_108141 : ~(_GEN_108253 & _GEN_1788) & _GEN_108141) : _GEN_108141;
  wire        _GEN_108376 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1789 & _GEN_108142 : _GEN_1104 ? ~_GEN_1789 & _GEN_108142 : ~(_GEN_108253 & _GEN_1789) & _GEN_108142) : _GEN_108142;
  wire        _GEN_108377 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1790 & _GEN_108143 : _GEN_1104 ? ~_GEN_1790 & _GEN_108143 : ~(_GEN_108253 & _GEN_1790) & _GEN_108143) : _GEN_108143;
  wire        _GEN_108378 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1791 & _GEN_108144 : _GEN_1104 ? ~_GEN_1791 & _GEN_108144 : ~(_GEN_108253 & _GEN_1791) & _GEN_108144) : _GEN_108144;
  wire        _GEN_108379 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1792 & _GEN_108145 : _GEN_1104 ? ~_GEN_1792 & _GEN_108145 : ~(_GEN_108253 & _GEN_1792) & _GEN_108145) : _GEN_108145;
  wire        _GEN_108380 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1793 & _GEN_108146 : _GEN_1104 ? ~_GEN_1793 & _GEN_108146 : ~(_GEN_108253 & _GEN_1793) & _GEN_108146) : _GEN_108146;
  wire        _GEN_108381 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1794 & _GEN_108147 : _GEN_1104 ? ~_GEN_1794 & _GEN_108147 : ~(_GEN_108253 & _GEN_1794) & _GEN_108147) : _GEN_108147;
  wire        _GEN_108382 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1795 & _GEN_108148 : _GEN_1104 ? ~_GEN_1795 & _GEN_108148 : ~(_GEN_108253 & _GEN_1795) & _GEN_108148) : _GEN_108148;
  wire        _GEN_108383 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1796 & _GEN_108149 : _GEN_1104 ? ~_GEN_1796 & _GEN_108149 : ~(_GEN_108253 & _GEN_1796) & _GEN_108149) : _GEN_108149;
  wire        _GEN_108384 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1797 & _GEN_108150 : _GEN_1104 ? ~_GEN_1797 & _GEN_108150 : ~(_GEN_108253 & _GEN_1797) & _GEN_108150) : _GEN_108150;
  wire        _GEN_108385 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1798 & _GEN_108151 : _GEN_1104 ? ~_GEN_1798 & _GEN_108151 : ~(_GEN_108253 & _GEN_1798) & _GEN_108151) : _GEN_108151;
  wire        _GEN_108386 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1799 & _GEN_108152 : _GEN_1104 ? ~_GEN_1799 & _GEN_108152 : ~(_GEN_108253 & _GEN_1799) & _GEN_108152) : _GEN_108152;
  wire        _GEN_108387 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1800 & _GEN_108153 : _GEN_1104 ? ~_GEN_1800 & _GEN_108153 : ~(_GEN_108253 & _GEN_1800) & _GEN_108153) : _GEN_108153;
  wire        _GEN_108388 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1801 & _GEN_108154 : _GEN_1104 ? ~_GEN_1801 & _GEN_108154 : ~(_GEN_108253 & _GEN_1801) & _GEN_108154) : _GEN_108154;
  wire        _GEN_108389 = _GEN_1102 ? (_GEN_108322 ? ~_GEN_1802 & _GEN_108155 : _GEN_1104 ? ~_GEN_1802 & _GEN_108155 : ~(_GEN_108253 & _GEN_1802) & _GEN_108155) : _GEN_108155;
  wire        _GEN_108390 = _GEN_1102 ? (_GEN_108322 ? ~(&lcam_ldq_idx_1) & _GEN_108156 : _GEN_1104 ? ~(&lcam_ldq_idx_1) & _GEN_108156 : ~(_GEN_108253 & (&lcam_ldq_idx_1)) & _GEN_108156) : _GEN_108156;
  wire        _GEN_108593 = _GEN_1105 ? (_GEN_108556 ? (|lcam_ldq_idx_0) & _GEN_108359 : _GEN_1107 ? (|lcam_ldq_idx_0) & _GEN_108359 : ~(_GEN_108721 & ~(|lcam_ldq_idx_0)) & _GEN_108359) : _GEN_108359;
  wire        _GEN_108594 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1743 & _GEN_108360 : _GEN_1107 ? ~_GEN_1743 & _GEN_108360 : ~(_GEN_108721 & _GEN_1743) & _GEN_108360) : _GEN_108360;
  wire        _GEN_108595 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1744 & _GEN_108361 : _GEN_1107 ? ~_GEN_1744 & _GEN_108361 : ~(_GEN_108721 & _GEN_1744) & _GEN_108361) : _GEN_108361;
  wire        _GEN_108596 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1745 & _GEN_108362 : _GEN_1107 ? ~_GEN_1745 & _GEN_108362 : ~(_GEN_108721 & _GEN_1745) & _GEN_108362) : _GEN_108362;
  wire        _GEN_108597 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1746 & _GEN_108363 : _GEN_1107 ? ~_GEN_1746 & _GEN_108363 : ~(_GEN_108721 & _GEN_1746) & _GEN_108363) : _GEN_108363;
  wire        _GEN_108598 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1747 & _GEN_108364 : _GEN_1107 ? ~_GEN_1747 & _GEN_108364 : ~(_GEN_108721 & _GEN_1747) & _GEN_108364) : _GEN_108364;
  wire        _GEN_108599 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1748 & _GEN_108365 : _GEN_1107 ? ~_GEN_1748 & _GEN_108365 : ~(_GEN_108721 & _GEN_1748) & _GEN_108365) : _GEN_108365;
  wire        _GEN_108600 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1749 & _GEN_108366 : _GEN_1107 ? ~_GEN_1749 & _GEN_108366 : ~(_GEN_108721 & _GEN_1749) & _GEN_108366) : _GEN_108366;
  wire        _GEN_108601 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1750 & _GEN_108367 : _GEN_1107 ? ~_GEN_1750 & _GEN_108367 : ~(_GEN_108721 & _GEN_1750) & _GEN_108367) : _GEN_108367;
  wire        _GEN_108602 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1751 & _GEN_108368 : _GEN_1107 ? ~_GEN_1751 & _GEN_108368 : ~(_GEN_108721 & _GEN_1751) & _GEN_108368) : _GEN_108368;
  wire        _GEN_108603 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1752 & _GEN_108369 : _GEN_1107 ? ~_GEN_1752 & _GEN_108369 : ~(_GEN_108721 & _GEN_1752) & _GEN_108369) : _GEN_108369;
  wire        _GEN_108604 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1753 & _GEN_108370 : _GEN_1107 ? ~_GEN_1753 & _GEN_108370 : ~(_GEN_108721 & _GEN_1753) & _GEN_108370) : _GEN_108370;
  wire        _GEN_108605 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1754 & _GEN_108371 : _GEN_1107 ? ~_GEN_1754 & _GEN_108371 : ~(_GEN_108721 & _GEN_1754) & _GEN_108371) : _GEN_108371;
  wire        _GEN_108606 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1755 & _GEN_108372 : _GEN_1107 ? ~_GEN_1755 & _GEN_108372 : ~(_GEN_108721 & _GEN_1755) & _GEN_108372) : _GEN_108372;
  wire        _GEN_108607 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1756 & _GEN_108373 : _GEN_1107 ? ~_GEN_1756 & _GEN_108373 : ~(_GEN_108721 & _GEN_1756) & _GEN_108373) : _GEN_108373;
  wire        _GEN_108608 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1757 & _GEN_108374 : _GEN_1107 ? ~_GEN_1757 & _GEN_108374 : ~(_GEN_108721 & _GEN_1757) & _GEN_108374) : _GEN_108374;
  wire        _GEN_108609 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1758 & _GEN_108375 : _GEN_1107 ? ~_GEN_1758 & _GEN_108375 : ~(_GEN_108721 & _GEN_1758) & _GEN_108375) : _GEN_108375;
  wire        _GEN_108610 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1759 & _GEN_108376 : _GEN_1107 ? ~_GEN_1759 & _GEN_108376 : ~(_GEN_108721 & _GEN_1759) & _GEN_108376) : _GEN_108376;
  wire        _GEN_108611 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1760 & _GEN_108377 : _GEN_1107 ? ~_GEN_1760 & _GEN_108377 : ~(_GEN_108721 & _GEN_1760) & _GEN_108377) : _GEN_108377;
  wire        _GEN_108612 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1761 & _GEN_108378 : _GEN_1107 ? ~_GEN_1761 & _GEN_108378 : ~(_GEN_108721 & _GEN_1761) & _GEN_108378) : _GEN_108378;
  wire        _GEN_108613 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1762 & _GEN_108379 : _GEN_1107 ? ~_GEN_1762 & _GEN_108379 : ~(_GEN_108721 & _GEN_1762) & _GEN_108379) : _GEN_108379;
  wire        _GEN_108614 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1763 & _GEN_108380 : _GEN_1107 ? ~_GEN_1763 & _GEN_108380 : ~(_GEN_108721 & _GEN_1763) & _GEN_108380) : _GEN_108380;
  wire        _GEN_108615 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1764 & _GEN_108381 : _GEN_1107 ? ~_GEN_1764 & _GEN_108381 : ~(_GEN_108721 & _GEN_1764) & _GEN_108381) : _GEN_108381;
  wire        _GEN_108616 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1765 & _GEN_108382 : _GEN_1107 ? ~_GEN_1765 & _GEN_108382 : ~(_GEN_108721 & _GEN_1765) & _GEN_108382) : _GEN_108382;
  wire        _GEN_108617 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1766 & _GEN_108383 : _GEN_1107 ? ~_GEN_1766 & _GEN_108383 : ~(_GEN_108721 & _GEN_1766) & _GEN_108383) : _GEN_108383;
  wire        _GEN_108618 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1767 & _GEN_108384 : _GEN_1107 ? ~_GEN_1767 & _GEN_108384 : ~(_GEN_108721 & _GEN_1767) & _GEN_108384) : _GEN_108384;
  wire        _GEN_108619 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1768 & _GEN_108385 : _GEN_1107 ? ~_GEN_1768 & _GEN_108385 : ~(_GEN_108721 & _GEN_1768) & _GEN_108385) : _GEN_108385;
  wire        _GEN_108620 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1769 & _GEN_108386 : _GEN_1107 ? ~_GEN_1769 & _GEN_108386 : ~(_GEN_108721 & _GEN_1769) & _GEN_108386) : _GEN_108386;
  wire        _GEN_108621 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1770 & _GEN_108387 : _GEN_1107 ? ~_GEN_1770 & _GEN_108387 : ~(_GEN_108721 & _GEN_1770) & _GEN_108387) : _GEN_108387;
  wire        _GEN_108622 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1771 & _GEN_108388 : _GEN_1107 ? ~_GEN_1771 & _GEN_108388 : ~(_GEN_108721 & _GEN_1771) & _GEN_108388) : _GEN_108388;
  wire        _GEN_108623 = _GEN_1105 ? (_GEN_108556 ? ~_GEN_1772 & _GEN_108389 : _GEN_1107 ? ~_GEN_1772 & _GEN_108389 : ~(_GEN_108721 & _GEN_1772) & _GEN_108389) : _GEN_108389;
  wire        _GEN_108624 = _GEN_1105 ? (_GEN_108556 ? ~(&lcam_ldq_idx_0) & _GEN_108390 : _GEN_1107 ? ~(&lcam_ldq_idx_0) & _GEN_108390 : ~(_GEN_108721 & (&lcam_ldq_idx_0)) & _GEN_108390) : _GEN_108390;
  wire        _GEN_108827 = _GEN_1108 ? (_GEN_108790 ? (|lcam_ldq_idx_1) & _GEN_108593 : _GEN_1110 ? (|lcam_ldq_idx_1) & _GEN_108593 : ~(_GEN_108721 & ~(|lcam_ldq_idx_1)) & _GEN_108593) : _GEN_108593;
  wire        _GEN_108828 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1773 & _GEN_108594 : _GEN_1110 ? ~_GEN_1773 & _GEN_108594 : ~(_GEN_108721 & _GEN_1773) & _GEN_108594) : _GEN_108594;
  wire        _GEN_108829 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1774 & _GEN_108595 : _GEN_1110 ? ~_GEN_1774 & _GEN_108595 : ~(_GEN_108721 & _GEN_1774) & _GEN_108595) : _GEN_108595;
  wire        _GEN_108830 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1775 & _GEN_108596 : _GEN_1110 ? ~_GEN_1775 & _GEN_108596 : ~(_GEN_108721 & _GEN_1775) & _GEN_108596) : _GEN_108596;
  wire        _GEN_108831 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1776 & _GEN_108597 : _GEN_1110 ? ~_GEN_1776 & _GEN_108597 : ~(_GEN_108721 & _GEN_1776) & _GEN_108597) : _GEN_108597;
  wire        _GEN_108832 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1777 & _GEN_108598 : _GEN_1110 ? ~_GEN_1777 & _GEN_108598 : ~(_GEN_108721 & _GEN_1777) & _GEN_108598) : _GEN_108598;
  wire        _GEN_108833 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1778 & _GEN_108599 : _GEN_1110 ? ~_GEN_1778 & _GEN_108599 : ~(_GEN_108721 & _GEN_1778) & _GEN_108599) : _GEN_108599;
  wire        _GEN_108834 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1779 & _GEN_108600 : _GEN_1110 ? ~_GEN_1779 & _GEN_108600 : ~(_GEN_108721 & _GEN_1779) & _GEN_108600) : _GEN_108600;
  wire        _GEN_108835 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1780 & _GEN_108601 : _GEN_1110 ? ~_GEN_1780 & _GEN_108601 : ~(_GEN_108721 & _GEN_1780) & _GEN_108601) : _GEN_108601;
  wire        _GEN_108836 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1781 & _GEN_108602 : _GEN_1110 ? ~_GEN_1781 & _GEN_108602 : ~(_GEN_108721 & _GEN_1781) & _GEN_108602) : _GEN_108602;
  wire        _GEN_108837 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1782 & _GEN_108603 : _GEN_1110 ? ~_GEN_1782 & _GEN_108603 : ~(_GEN_108721 & _GEN_1782) & _GEN_108603) : _GEN_108603;
  wire        _GEN_108838 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1783 & _GEN_108604 : _GEN_1110 ? ~_GEN_1783 & _GEN_108604 : ~(_GEN_108721 & _GEN_1783) & _GEN_108604) : _GEN_108604;
  wire        _GEN_108839 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1784 & _GEN_108605 : _GEN_1110 ? ~_GEN_1784 & _GEN_108605 : ~(_GEN_108721 & _GEN_1784) & _GEN_108605) : _GEN_108605;
  wire        _GEN_108840 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1785 & _GEN_108606 : _GEN_1110 ? ~_GEN_1785 & _GEN_108606 : ~(_GEN_108721 & _GEN_1785) & _GEN_108606) : _GEN_108606;
  wire        _GEN_108841 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1786 & _GEN_108607 : _GEN_1110 ? ~_GEN_1786 & _GEN_108607 : ~(_GEN_108721 & _GEN_1786) & _GEN_108607) : _GEN_108607;
  wire        _GEN_108842 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1787 & _GEN_108608 : _GEN_1110 ? ~_GEN_1787 & _GEN_108608 : ~(_GEN_108721 & _GEN_1787) & _GEN_108608) : _GEN_108608;
  wire        _GEN_108843 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1788 & _GEN_108609 : _GEN_1110 ? ~_GEN_1788 & _GEN_108609 : ~(_GEN_108721 & _GEN_1788) & _GEN_108609) : _GEN_108609;
  wire        _GEN_108844 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1789 & _GEN_108610 : _GEN_1110 ? ~_GEN_1789 & _GEN_108610 : ~(_GEN_108721 & _GEN_1789) & _GEN_108610) : _GEN_108610;
  wire        _GEN_108845 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1790 & _GEN_108611 : _GEN_1110 ? ~_GEN_1790 & _GEN_108611 : ~(_GEN_108721 & _GEN_1790) & _GEN_108611) : _GEN_108611;
  wire        _GEN_108846 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1791 & _GEN_108612 : _GEN_1110 ? ~_GEN_1791 & _GEN_108612 : ~(_GEN_108721 & _GEN_1791) & _GEN_108612) : _GEN_108612;
  wire        _GEN_108847 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1792 & _GEN_108613 : _GEN_1110 ? ~_GEN_1792 & _GEN_108613 : ~(_GEN_108721 & _GEN_1792) & _GEN_108613) : _GEN_108613;
  wire        _GEN_108848 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1793 & _GEN_108614 : _GEN_1110 ? ~_GEN_1793 & _GEN_108614 : ~(_GEN_108721 & _GEN_1793) & _GEN_108614) : _GEN_108614;
  wire        _GEN_108849 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1794 & _GEN_108615 : _GEN_1110 ? ~_GEN_1794 & _GEN_108615 : ~(_GEN_108721 & _GEN_1794) & _GEN_108615) : _GEN_108615;
  wire        _GEN_108850 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1795 & _GEN_108616 : _GEN_1110 ? ~_GEN_1795 & _GEN_108616 : ~(_GEN_108721 & _GEN_1795) & _GEN_108616) : _GEN_108616;
  wire        _GEN_108851 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1796 & _GEN_108617 : _GEN_1110 ? ~_GEN_1796 & _GEN_108617 : ~(_GEN_108721 & _GEN_1796) & _GEN_108617) : _GEN_108617;
  wire        _GEN_108852 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1797 & _GEN_108618 : _GEN_1110 ? ~_GEN_1797 & _GEN_108618 : ~(_GEN_108721 & _GEN_1797) & _GEN_108618) : _GEN_108618;
  wire        _GEN_108853 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1798 & _GEN_108619 : _GEN_1110 ? ~_GEN_1798 & _GEN_108619 : ~(_GEN_108721 & _GEN_1798) & _GEN_108619) : _GEN_108619;
  wire        _GEN_108854 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1799 & _GEN_108620 : _GEN_1110 ? ~_GEN_1799 & _GEN_108620 : ~(_GEN_108721 & _GEN_1799) & _GEN_108620) : _GEN_108620;
  wire        _GEN_108855 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1800 & _GEN_108621 : _GEN_1110 ? ~_GEN_1800 & _GEN_108621 : ~(_GEN_108721 & _GEN_1800) & _GEN_108621) : _GEN_108621;
  wire        _GEN_108856 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1801 & _GEN_108622 : _GEN_1110 ? ~_GEN_1801 & _GEN_108622 : ~(_GEN_108721 & _GEN_1801) & _GEN_108622) : _GEN_108622;
  wire        _GEN_108857 = _GEN_1108 ? (_GEN_108790 ? ~_GEN_1802 & _GEN_108623 : _GEN_1110 ? ~_GEN_1802 & _GEN_108623 : ~(_GEN_108721 & _GEN_1802) & _GEN_108623) : _GEN_108623;
  wire        _GEN_108858 = _GEN_1108 ? (_GEN_108790 ? ~(&lcam_ldq_idx_1) & _GEN_108624 : _GEN_1110 ? ~(&lcam_ldq_idx_1) & _GEN_108624 : ~(_GEN_108721 & (&lcam_ldq_idx_1)) & _GEN_108624) : _GEN_108624;
  wire        _GEN_109061 = _GEN_1111 ? (_GEN_109024 ? (|lcam_ldq_idx_0) & _GEN_108827 : _GEN_1113 ? (|lcam_ldq_idx_0) & _GEN_108827 : ~(_GEN_109189 & ~(|lcam_ldq_idx_0)) & _GEN_108827) : _GEN_108827;
  wire        _GEN_109062 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1743 & _GEN_108828 : _GEN_1113 ? ~_GEN_1743 & _GEN_108828 : ~(_GEN_109189 & _GEN_1743) & _GEN_108828) : _GEN_108828;
  wire        _GEN_109063 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1744 & _GEN_108829 : _GEN_1113 ? ~_GEN_1744 & _GEN_108829 : ~(_GEN_109189 & _GEN_1744) & _GEN_108829) : _GEN_108829;
  wire        _GEN_109064 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1745 & _GEN_108830 : _GEN_1113 ? ~_GEN_1745 & _GEN_108830 : ~(_GEN_109189 & _GEN_1745) & _GEN_108830) : _GEN_108830;
  wire        _GEN_109065 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1746 & _GEN_108831 : _GEN_1113 ? ~_GEN_1746 & _GEN_108831 : ~(_GEN_109189 & _GEN_1746) & _GEN_108831) : _GEN_108831;
  wire        _GEN_109066 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1747 & _GEN_108832 : _GEN_1113 ? ~_GEN_1747 & _GEN_108832 : ~(_GEN_109189 & _GEN_1747) & _GEN_108832) : _GEN_108832;
  wire        _GEN_109067 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1748 & _GEN_108833 : _GEN_1113 ? ~_GEN_1748 & _GEN_108833 : ~(_GEN_109189 & _GEN_1748) & _GEN_108833) : _GEN_108833;
  wire        _GEN_109068 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1749 & _GEN_108834 : _GEN_1113 ? ~_GEN_1749 & _GEN_108834 : ~(_GEN_109189 & _GEN_1749) & _GEN_108834) : _GEN_108834;
  wire        _GEN_109069 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1750 & _GEN_108835 : _GEN_1113 ? ~_GEN_1750 & _GEN_108835 : ~(_GEN_109189 & _GEN_1750) & _GEN_108835) : _GEN_108835;
  wire        _GEN_109070 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1751 & _GEN_108836 : _GEN_1113 ? ~_GEN_1751 & _GEN_108836 : ~(_GEN_109189 & _GEN_1751) & _GEN_108836) : _GEN_108836;
  wire        _GEN_109071 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1752 & _GEN_108837 : _GEN_1113 ? ~_GEN_1752 & _GEN_108837 : ~(_GEN_109189 & _GEN_1752) & _GEN_108837) : _GEN_108837;
  wire        _GEN_109072 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1753 & _GEN_108838 : _GEN_1113 ? ~_GEN_1753 & _GEN_108838 : ~(_GEN_109189 & _GEN_1753) & _GEN_108838) : _GEN_108838;
  wire        _GEN_109073 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1754 & _GEN_108839 : _GEN_1113 ? ~_GEN_1754 & _GEN_108839 : ~(_GEN_109189 & _GEN_1754) & _GEN_108839) : _GEN_108839;
  wire        _GEN_109074 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1755 & _GEN_108840 : _GEN_1113 ? ~_GEN_1755 & _GEN_108840 : ~(_GEN_109189 & _GEN_1755) & _GEN_108840) : _GEN_108840;
  wire        _GEN_109075 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1756 & _GEN_108841 : _GEN_1113 ? ~_GEN_1756 & _GEN_108841 : ~(_GEN_109189 & _GEN_1756) & _GEN_108841) : _GEN_108841;
  wire        _GEN_109076 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1757 & _GEN_108842 : _GEN_1113 ? ~_GEN_1757 & _GEN_108842 : ~(_GEN_109189 & _GEN_1757) & _GEN_108842) : _GEN_108842;
  wire        _GEN_109077 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1758 & _GEN_108843 : _GEN_1113 ? ~_GEN_1758 & _GEN_108843 : ~(_GEN_109189 & _GEN_1758) & _GEN_108843) : _GEN_108843;
  wire        _GEN_109078 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1759 & _GEN_108844 : _GEN_1113 ? ~_GEN_1759 & _GEN_108844 : ~(_GEN_109189 & _GEN_1759) & _GEN_108844) : _GEN_108844;
  wire        _GEN_109079 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1760 & _GEN_108845 : _GEN_1113 ? ~_GEN_1760 & _GEN_108845 : ~(_GEN_109189 & _GEN_1760) & _GEN_108845) : _GEN_108845;
  wire        _GEN_109080 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1761 & _GEN_108846 : _GEN_1113 ? ~_GEN_1761 & _GEN_108846 : ~(_GEN_109189 & _GEN_1761) & _GEN_108846) : _GEN_108846;
  wire        _GEN_109081 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1762 & _GEN_108847 : _GEN_1113 ? ~_GEN_1762 & _GEN_108847 : ~(_GEN_109189 & _GEN_1762) & _GEN_108847) : _GEN_108847;
  wire        _GEN_109082 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1763 & _GEN_108848 : _GEN_1113 ? ~_GEN_1763 & _GEN_108848 : ~(_GEN_109189 & _GEN_1763) & _GEN_108848) : _GEN_108848;
  wire        _GEN_109083 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1764 & _GEN_108849 : _GEN_1113 ? ~_GEN_1764 & _GEN_108849 : ~(_GEN_109189 & _GEN_1764) & _GEN_108849) : _GEN_108849;
  wire        _GEN_109084 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1765 & _GEN_108850 : _GEN_1113 ? ~_GEN_1765 & _GEN_108850 : ~(_GEN_109189 & _GEN_1765) & _GEN_108850) : _GEN_108850;
  wire        _GEN_109085 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1766 & _GEN_108851 : _GEN_1113 ? ~_GEN_1766 & _GEN_108851 : ~(_GEN_109189 & _GEN_1766) & _GEN_108851) : _GEN_108851;
  wire        _GEN_109086 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1767 & _GEN_108852 : _GEN_1113 ? ~_GEN_1767 & _GEN_108852 : ~(_GEN_109189 & _GEN_1767) & _GEN_108852) : _GEN_108852;
  wire        _GEN_109087 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1768 & _GEN_108853 : _GEN_1113 ? ~_GEN_1768 & _GEN_108853 : ~(_GEN_109189 & _GEN_1768) & _GEN_108853) : _GEN_108853;
  wire        _GEN_109088 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1769 & _GEN_108854 : _GEN_1113 ? ~_GEN_1769 & _GEN_108854 : ~(_GEN_109189 & _GEN_1769) & _GEN_108854) : _GEN_108854;
  wire        _GEN_109089 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1770 & _GEN_108855 : _GEN_1113 ? ~_GEN_1770 & _GEN_108855 : ~(_GEN_109189 & _GEN_1770) & _GEN_108855) : _GEN_108855;
  wire        _GEN_109090 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1771 & _GEN_108856 : _GEN_1113 ? ~_GEN_1771 & _GEN_108856 : ~(_GEN_109189 & _GEN_1771) & _GEN_108856) : _GEN_108856;
  wire        _GEN_109091 = _GEN_1111 ? (_GEN_109024 ? ~_GEN_1772 & _GEN_108857 : _GEN_1113 ? ~_GEN_1772 & _GEN_108857 : ~(_GEN_109189 & _GEN_1772) & _GEN_108857) : _GEN_108857;
  wire        _GEN_109092 = _GEN_1111 ? (_GEN_109024 ? ~(&lcam_ldq_idx_0) & _GEN_108858 : _GEN_1113 ? ~(&lcam_ldq_idx_0) & _GEN_108858 : ~(_GEN_109189 & (&lcam_ldq_idx_0)) & _GEN_108858) : _GEN_108858;
  wire        _GEN_109295 = _GEN_1114 ? (_GEN_109258 ? (|lcam_ldq_idx_1) & _GEN_109061 : _GEN_1116 ? (|lcam_ldq_idx_1) & _GEN_109061 : ~(_GEN_109189 & ~(|lcam_ldq_idx_1)) & _GEN_109061) : _GEN_109061;
  wire        _GEN_109296 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1773 & _GEN_109062 : _GEN_1116 ? ~_GEN_1773 & _GEN_109062 : ~(_GEN_109189 & _GEN_1773) & _GEN_109062) : _GEN_109062;
  wire        _GEN_109297 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1774 & _GEN_109063 : _GEN_1116 ? ~_GEN_1774 & _GEN_109063 : ~(_GEN_109189 & _GEN_1774) & _GEN_109063) : _GEN_109063;
  wire        _GEN_109298 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1775 & _GEN_109064 : _GEN_1116 ? ~_GEN_1775 & _GEN_109064 : ~(_GEN_109189 & _GEN_1775) & _GEN_109064) : _GEN_109064;
  wire        _GEN_109299 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1776 & _GEN_109065 : _GEN_1116 ? ~_GEN_1776 & _GEN_109065 : ~(_GEN_109189 & _GEN_1776) & _GEN_109065) : _GEN_109065;
  wire        _GEN_109300 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1777 & _GEN_109066 : _GEN_1116 ? ~_GEN_1777 & _GEN_109066 : ~(_GEN_109189 & _GEN_1777) & _GEN_109066) : _GEN_109066;
  wire        _GEN_109301 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1778 & _GEN_109067 : _GEN_1116 ? ~_GEN_1778 & _GEN_109067 : ~(_GEN_109189 & _GEN_1778) & _GEN_109067) : _GEN_109067;
  wire        _GEN_109302 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1779 & _GEN_109068 : _GEN_1116 ? ~_GEN_1779 & _GEN_109068 : ~(_GEN_109189 & _GEN_1779) & _GEN_109068) : _GEN_109068;
  wire        _GEN_109303 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1780 & _GEN_109069 : _GEN_1116 ? ~_GEN_1780 & _GEN_109069 : ~(_GEN_109189 & _GEN_1780) & _GEN_109069) : _GEN_109069;
  wire        _GEN_109304 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1781 & _GEN_109070 : _GEN_1116 ? ~_GEN_1781 & _GEN_109070 : ~(_GEN_109189 & _GEN_1781) & _GEN_109070) : _GEN_109070;
  wire        _GEN_109305 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1782 & _GEN_109071 : _GEN_1116 ? ~_GEN_1782 & _GEN_109071 : ~(_GEN_109189 & _GEN_1782) & _GEN_109071) : _GEN_109071;
  wire        _GEN_109306 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1783 & _GEN_109072 : _GEN_1116 ? ~_GEN_1783 & _GEN_109072 : ~(_GEN_109189 & _GEN_1783) & _GEN_109072) : _GEN_109072;
  wire        _GEN_109307 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1784 & _GEN_109073 : _GEN_1116 ? ~_GEN_1784 & _GEN_109073 : ~(_GEN_109189 & _GEN_1784) & _GEN_109073) : _GEN_109073;
  wire        _GEN_109308 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1785 & _GEN_109074 : _GEN_1116 ? ~_GEN_1785 & _GEN_109074 : ~(_GEN_109189 & _GEN_1785) & _GEN_109074) : _GEN_109074;
  wire        _GEN_109309 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1786 & _GEN_109075 : _GEN_1116 ? ~_GEN_1786 & _GEN_109075 : ~(_GEN_109189 & _GEN_1786) & _GEN_109075) : _GEN_109075;
  wire        _GEN_109310 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1787 & _GEN_109076 : _GEN_1116 ? ~_GEN_1787 & _GEN_109076 : ~(_GEN_109189 & _GEN_1787) & _GEN_109076) : _GEN_109076;
  wire        _GEN_109311 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1788 & _GEN_109077 : _GEN_1116 ? ~_GEN_1788 & _GEN_109077 : ~(_GEN_109189 & _GEN_1788) & _GEN_109077) : _GEN_109077;
  wire        _GEN_109312 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1789 & _GEN_109078 : _GEN_1116 ? ~_GEN_1789 & _GEN_109078 : ~(_GEN_109189 & _GEN_1789) & _GEN_109078) : _GEN_109078;
  wire        _GEN_109313 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1790 & _GEN_109079 : _GEN_1116 ? ~_GEN_1790 & _GEN_109079 : ~(_GEN_109189 & _GEN_1790) & _GEN_109079) : _GEN_109079;
  wire        _GEN_109314 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1791 & _GEN_109080 : _GEN_1116 ? ~_GEN_1791 & _GEN_109080 : ~(_GEN_109189 & _GEN_1791) & _GEN_109080) : _GEN_109080;
  wire        _GEN_109315 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1792 & _GEN_109081 : _GEN_1116 ? ~_GEN_1792 & _GEN_109081 : ~(_GEN_109189 & _GEN_1792) & _GEN_109081) : _GEN_109081;
  wire        _GEN_109316 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1793 & _GEN_109082 : _GEN_1116 ? ~_GEN_1793 & _GEN_109082 : ~(_GEN_109189 & _GEN_1793) & _GEN_109082) : _GEN_109082;
  wire        _GEN_109317 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1794 & _GEN_109083 : _GEN_1116 ? ~_GEN_1794 & _GEN_109083 : ~(_GEN_109189 & _GEN_1794) & _GEN_109083) : _GEN_109083;
  wire        _GEN_109318 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1795 & _GEN_109084 : _GEN_1116 ? ~_GEN_1795 & _GEN_109084 : ~(_GEN_109189 & _GEN_1795) & _GEN_109084) : _GEN_109084;
  wire        _GEN_109319 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1796 & _GEN_109085 : _GEN_1116 ? ~_GEN_1796 & _GEN_109085 : ~(_GEN_109189 & _GEN_1796) & _GEN_109085) : _GEN_109085;
  wire        _GEN_109320 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1797 & _GEN_109086 : _GEN_1116 ? ~_GEN_1797 & _GEN_109086 : ~(_GEN_109189 & _GEN_1797) & _GEN_109086) : _GEN_109086;
  wire        _GEN_109321 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1798 & _GEN_109087 : _GEN_1116 ? ~_GEN_1798 & _GEN_109087 : ~(_GEN_109189 & _GEN_1798) & _GEN_109087) : _GEN_109087;
  wire        _GEN_109322 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1799 & _GEN_109088 : _GEN_1116 ? ~_GEN_1799 & _GEN_109088 : ~(_GEN_109189 & _GEN_1799) & _GEN_109088) : _GEN_109088;
  wire        _GEN_109323 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1800 & _GEN_109089 : _GEN_1116 ? ~_GEN_1800 & _GEN_109089 : ~(_GEN_109189 & _GEN_1800) & _GEN_109089) : _GEN_109089;
  wire        _GEN_109324 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1801 & _GEN_109090 : _GEN_1116 ? ~_GEN_1801 & _GEN_109090 : ~(_GEN_109189 & _GEN_1801) & _GEN_109090) : _GEN_109090;
  wire        _GEN_109325 = _GEN_1114 ? (_GEN_109258 ? ~_GEN_1802 & _GEN_109091 : _GEN_1116 ? ~_GEN_1802 & _GEN_109091 : ~(_GEN_109189 & _GEN_1802) & _GEN_109091) : _GEN_109091;
  wire        _GEN_109326 = _GEN_1114 ? (_GEN_109258 ? ~(&lcam_ldq_idx_1) & _GEN_109092 : _GEN_1116 ? ~(&lcam_ldq_idx_1) & _GEN_109092 : ~(_GEN_109189 & (&lcam_ldq_idx_1)) & _GEN_109092) : _GEN_109092;
  wire        _GEN_109529 = _GEN_1117 ? (_GEN_109492 ? (|lcam_ldq_idx_0) & _GEN_109295 : _GEN_1119 ? (|lcam_ldq_idx_0) & _GEN_109295 : ~(_GEN_109657 & ~(|lcam_ldq_idx_0)) & _GEN_109295) : _GEN_109295;
  wire        _GEN_109530 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1743 & _GEN_109296 : _GEN_1119 ? ~_GEN_1743 & _GEN_109296 : ~(_GEN_109657 & _GEN_1743) & _GEN_109296) : _GEN_109296;
  wire        _GEN_109531 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1744 & _GEN_109297 : _GEN_1119 ? ~_GEN_1744 & _GEN_109297 : ~(_GEN_109657 & _GEN_1744) & _GEN_109297) : _GEN_109297;
  wire        _GEN_109532 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1745 & _GEN_109298 : _GEN_1119 ? ~_GEN_1745 & _GEN_109298 : ~(_GEN_109657 & _GEN_1745) & _GEN_109298) : _GEN_109298;
  wire        _GEN_109533 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1746 & _GEN_109299 : _GEN_1119 ? ~_GEN_1746 & _GEN_109299 : ~(_GEN_109657 & _GEN_1746) & _GEN_109299) : _GEN_109299;
  wire        _GEN_109534 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1747 & _GEN_109300 : _GEN_1119 ? ~_GEN_1747 & _GEN_109300 : ~(_GEN_109657 & _GEN_1747) & _GEN_109300) : _GEN_109300;
  wire        _GEN_109535 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1748 & _GEN_109301 : _GEN_1119 ? ~_GEN_1748 & _GEN_109301 : ~(_GEN_109657 & _GEN_1748) & _GEN_109301) : _GEN_109301;
  wire        _GEN_109536 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1749 & _GEN_109302 : _GEN_1119 ? ~_GEN_1749 & _GEN_109302 : ~(_GEN_109657 & _GEN_1749) & _GEN_109302) : _GEN_109302;
  wire        _GEN_109537 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1750 & _GEN_109303 : _GEN_1119 ? ~_GEN_1750 & _GEN_109303 : ~(_GEN_109657 & _GEN_1750) & _GEN_109303) : _GEN_109303;
  wire        _GEN_109538 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1751 & _GEN_109304 : _GEN_1119 ? ~_GEN_1751 & _GEN_109304 : ~(_GEN_109657 & _GEN_1751) & _GEN_109304) : _GEN_109304;
  wire        _GEN_109539 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1752 & _GEN_109305 : _GEN_1119 ? ~_GEN_1752 & _GEN_109305 : ~(_GEN_109657 & _GEN_1752) & _GEN_109305) : _GEN_109305;
  wire        _GEN_109540 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1753 & _GEN_109306 : _GEN_1119 ? ~_GEN_1753 & _GEN_109306 : ~(_GEN_109657 & _GEN_1753) & _GEN_109306) : _GEN_109306;
  wire        _GEN_109541 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1754 & _GEN_109307 : _GEN_1119 ? ~_GEN_1754 & _GEN_109307 : ~(_GEN_109657 & _GEN_1754) & _GEN_109307) : _GEN_109307;
  wire        _GEN_109542 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1755 & _GEN_109308 : _GEN_1119 ? ~_GEN_1755 & _GEN_109308 : ~(_GEN_109657 & _GEN_1755) & _GEN_109308) : _GEN_109308;
  wire        _GEN_109543 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1756 & _GEN_109309 : _GEN_1119 ? ~_GEN_1756 & _GEN_109309 : ~(_GEN_109657 & _GEN_1756) & _GEN_109309) : _GEN_109309;
  wire        _GEN_109544 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1757 & _GEN_109310 : _GEN_1119 ? ~_GEN_1757 & _GEN_109310 : ~(_GEN_109657 & _GEN_1757) & _GEN_109310) : _GEN_109310;
  wire        _GEN_109545 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1758 & _GEN_109311 : _GEN_1119 ? ~_GEN_1758 & _GEN_109311 : ~(_GEN_109657 & _GEN_1758) & _GEN_109311) : _GEN_109311;
  wire        _GEN_109546 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1759 & _GEN_109312 : _GEN_1119 ? ~_GEN_1759 & _GEN_109312 : ~(_GEN_109657 & _GEN_1759) & _GEN_109312) : _GEN_109312;
  wire        _GEN_109547 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1760 & _GEN_109313 : _GEN_1119 ? ~_GEN_1760 & _GEN_109313 : ~(_GEN_109657 & _GEN_1760) & _GEN_109313) : _GEN_109313;
  wire        _GEN_109548 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1761 & _GEN_109314 : _GEN_1119 ? ~_GEN_1761 & _GEN_109314 : ~(_GEN_109657 & _GEN_1761) & _GEN_109314) : _GEN_109314;
  wire        _GEN_109549 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1762 & _GEN_109315 : _GEN_1119 ? ~_GEN_1762 & _GEN_109315 : ~(_GEN_109657 & _GEN_1762) & _GEN_109315) : _GEN_109315;
  wire        _GEN_109550 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1763 & _GEN_109316 : _GEN_1119 ? ~_GEN_1763 & _GEN_109316 : ~(_GEN_109657 & _GEN_1763) & _GEN_109316) : _GEN_109316;
  wire        _GEN_109551 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1764 & _GEN_109317 : _GEN_1119 ? ~_GEN_1764 & _GEN_109317 : ~(_GEN_109657 & _GEN_1764) & _GEN_109317) : _GEN_109317;
  wire        _GEN_109552 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1765 & _GEN_109318 : _GEN_1119 ? ~_GEN_1765 & _GEN_109318 : ~(_GEN_109657 & _GEN_1765) & _GEN_109318) : _GEN_109318;
  wire        _GEN_109553 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1766 & _GEN_109319 : _GEN_1119 ? ~_GEN_1766 & _GEN_109319 : ~(_GEN_109657 & _GEN_1766) & _GEN_109319) : _GEN_109319;
  wire        _GEN_109554 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1767 & _GEN_109320 : _GEN_1119 ? ~_GEN_1767 & _GEN_109320 : ~(_GEN_109657 & _GEN_1767) & _GEN_109320) : _GEN_109320;
  wire        _GEN_109555 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1768 & _GEN_109321 : _GEN_1119 ? ~_GEN_1768 & _GEN_109321 : ~(_GEN_109657 & _GEN_1768) & _GEN_109321) : _GEN_109321;
  wire        _GEN_109556 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1769 & _GEN_109322 : _GEN_1119 ? ~_GEN_1769 & _GEN_109322 : ~(_GEN_109657 & _GEN_1769) & _GEN_109322) : _GEN_109322;
  wire        _GEN_109557 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1770 & _GEN_109323 : _GEN_1119 ? ~_GEN_1770 & _GEN_109323 : ~(_GEN_109657 & _GEN_1770) & _GEN_109323) : _GEN_109323;
  wire        _GEN_109558 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1771 & _GEN_109324 : _GEN_1119 ? ~_GEN_1771 & _GEN_109324 : ~(_GEN_109657 & _GEN_1771) & _GEN_109324) : _GEN_109324;
  wire        _GEN_109559 = _GEN_1117 ? (_GEN_109492 ? ~_GEN_1772 & _GEN_109325 : _GEN_1119 ? ~_GEN_1772 & _GEN_109325 : ~(_GEN_109657 & _GEN_1772) & _GEN_109325) : _GEN_109325;
  wire        _GEN_109560 = _GEN_1117 ? (_GEN_109492 ? ~(&lcam_ldq_idx_0) & _GEN_109326 : _GEN_1119 ? ~(&lcam_ldq_idx_0) & _GEN_109326 : ~(_GEN_109657 & (&lcam_ldq_idx_0)) & _GEN_109326) : _GEN_109326;
  wire        _GEN_109763 = _GEN_1120 ? (_GEN_109726 ? (|lcam_ldq_idx_1) & _GEN_109529 : _GEN_1122 ? (|lcam_ldq_idx_1) & _GEN_109529 : ~(_GEN_109657 & ~(|lcam_ldq_idx_1)) & _GEN_109529) : _GEN_109529;
  wire        _GEN_109764 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1773 & _GEN_109530 : _GEN_1122 ? ~_GEN_1773 & _GEN_109530 : ~(_GEN_109657 & _GEN_1773) & _GEN_109530) : _GEN_109530;
  wire        _GEN_109765 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1774 & _GEN_109531 : _GEN_1122 ? ~_GEN_1774 & _GEN_109531 : ~(_GEN_109657 & _GEN_1774) & _GEN_109531) : _GEN_109531;
  wire        _GEN_109766 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1775 & _GEN_109532 : _GEN_1122 ? ~_GEN_1775 & _GEN_109532 : ~(_GEN_109657 & _GEN_1775) & _GEN_109532) : _GEN_109532;
  wire        _GEN_109767 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1776 & _GEN_109533 : _GEN_1122 ? ~_GEN_1776 & _GEN_109533 : ~(_GEN_109657 & _GEN_1776) & _GEN_109533) : _GEN_109533;
  wire        _GEN_109768 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1777 & _GEN_109534 : _GEN_1122 ? ~_GEN_1777 & _GEN_109534 : ~(_GEN_109657 & _GEN_1777) & _GEN_109534) : _GEN_109534;
  wire        _GEN_109769 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1778 & _GEN_109535 : _GEN_1122 ? ~_GEN_1778 & _GEN_109535 : ~(_GEN_109657 & _GEN_1778) & _GEN_109535) : _GEN_109535;
  wire        _GEN_109770 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1779 & _GEN_109536 : _GEN_1122 ? ~_GEN_1779 & _GEN_109536 : ~(_GEN_109657 & _GEN_1779) & _GEN_109536) : _GEN_109536;
  wire        _GEN_109771 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1780 & _GEN_109537 : _GEN_1122 ? ~_GEN_1780 & _GEN_109537 : ~(_GEN_109657 & _GEN_1780) & _GEN_109537) : _GEN_109537;
  wire        _GEN_109772 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1781 & _GEN_109538 : _GEN_1122 ? ~_GEN_1781 & _GEN_109538 : ~(_GEN_109657 & _GEN_1781) & _GEN_109538) : _GEN_109538;
  wire        _GEN_109773 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1782 & _GEN_109539 : _GEN_1122 ? ~_GEN_1782 & _GEN_109539 : ~(_GEN_109657 & _GEN_1782) & _GEN_109539) : _GEN_109539;
  wire        _GEN_109774 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1783 & _GEN_109540 : _GEN_1122 ? ~_GEN_1783 & _GEN_109540 : ~(_GEN_109657 & _GEN_1783) & _GEN_109540) : _GEN_109540;
  wire        _GEN_109775 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1784 & _GEN_109541 : _GEN_1122 ? ~_GEN_1784 & _GEN_109541 : ~(_GEN_109657 & _GEN_1784) & _GEN_109541) : _GEN_109541;
  wire        _GEN_109776 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1785 & _GEN_109542 : _GEN_1122 ? ~_GEN_1785 & _GEN_109542 : ~(_GEN_109657 & _GEN_1785) & _GEN_109542) : _GEN_109542;
  wire        _GEN_109777 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1786 & _GEN_109543 : _GEN_1122 ? ~_GEN_1786 & _GEN_109543 : ~(_GEN_109657 & _GEN_1786) & _GEN_109543) : _GEN_109543;
  wire        _GEN_109778 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1787 & _GEN_109544 : _GEN_1122 ? ~_GEN_1787 & _GEN_109544 : ~(_GEN_109657 & _GEN_1787) & _GEN_109544) : _GEN_109544;
  wire        _GEN_109779 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1788 & _GEN_109545 : _GEN_1122 ? ~_GEN_1788 & _GEN_109545 : ~(_GEN_109657 & _GEN_1788) & _GEN_109545) : _GEN_109545;
  wire        _GEN_109780 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1789 & _GEN_109546 : _GEN_1122 ? ~_GEN_1789 & _GEN_109546 : ~(_GEN_109657 & _GEN_1789) & _GEN_109546) : _GEN_109546;
  wire        _GEN_109781 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1790 & _GEN_109547 : _GEN_1122 ? ~_GEN_1790 & _GEN_109547 : ~(_GEN_109657 & _GEN_1790) & _GEN_109547) : _GEN_109547;
  wire        _GEN_109782 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1791 & _GEN_109548 : _GEN_1122 ? ~_GEN_1791 & _GEN_109548 : ~(_GEN_109657 & _GEN_1791) & _GEN_109548) : _GEN_109548;
  wire        _GEN_109783 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1792 & _GEN_109549 : _GEN_1122 ? ~_GEN_1792 & _GEN_109549 : ~(_GEN_109657 & _GEN_1792) & _GEN_109549) : _GEN_109549;
  wire        _GEN_109784 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1793 & _GEN_109550 : _GEN_1122 ? ~_GEN_1793 & _GEN_109550 : ~(_GEN_109657 & _GEN_1793) & _GEN_109550) : _GEN_109550;
  wire        _GEN_109785 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1794 & _GEN_109551 : _GEN_1122 ? ~_GEN_1794 & _GEN_109551 : ~(_GEN_109657 & _GEN_1794) & _GEN_109551) : _GEN_109551;
  wire        _GEN_109786 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1795 & _GEN_109552 : _GEN_1122 ? ~_GEN_1795 & _GEN_109552 : ~(_GEN_109657 & _GEN_1795) & _GEN_109552) : _GEN_109552;
  wire        _GEN_109787 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1796 & _GEN_109553 : _GEN_1122 ? ~_GEN_1796 & _GEN_109553 : ~(_GEN_109657 & _GEN_1796) & _GEN_109553) : _GEN_109553;
  wire        _GEN_109788 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1797 & _GEN_109554 : _GEN_1122 ? ~_GEN_1797 & _GEN_109554 : ~(_GEN_109657 & _GEN_1797) & _GEN_109554) : _GEN_109554;
  wire        _GEN_109789 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1798 & _GEN_109555 : _GEN_1122 ? ~_GEN_1798 & _GEN_109555 : ~(_GEN_109657 & _GEN_1798) & _GEN_109555) : _GEN_109555;
  wire        _GEN_109790 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1799 & _GEN_109556 : _GEN_1122 ? ~_GEN_1799 & _GEN_109556 : ~(_GEN_109657 & _GEN_1799) & _GEN_109556) : _GEN_109556;
  wire        _GEN_109791 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1800 & _GEN_109557 : _GEN_1122 ? ~_GEN_1800 & _GEN_109557 : ~(_GEN_109657 & _GEN_1800) & _GEN_109557) : _GEN_109557;
  wire        _GEN_109792 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1801 & _GEN_109558 : _GEN_1122 ? ~_GEN_1801 & _GEN_109558 : ~(_GEN_109657 & _GEN_1801) & _GEN_109558) : _GEN_109558;
  wire        _GEN_109793 = _GEN_1120 ? (_GEN_109726 ? ~_GEN_1802 & _GEN_109559 : _GEN_1122 ? ~_GEN_1802 & _GEN_109559 : ~(_GEN_109657 & _GEN_1802) & _GEN_109559) : _GEN_109559;
  wire        _GEN_109794 = _GEN_1120 ? (_GEN_109726 ? ~(&lcam_ldq_idx_1) & _GEN_109560 : _GEN_1122 ? ~(&lcam_ldq_idx_1) & _GEN_109560 : ~(_GEN_109657 & (&lcam_ldq_idx_1)) & _GEN_109560) : _GEN_109560;
  wire        _GEN_109997 = _GEN_1123 ? (_GEN_109960 ? (|lcam_ldq_idx_0) & _GEN_109763 : _GEN_1125 ? (|lcam_ldq_idx_0) & _GEN_109763 : ~(_GEN_110125 & ~(|lcam_ldq_idx_0)) & _GEN_109763) : _GEN_109763;
  wire        _GEN_109998 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1743 & _GEN_109764 : _GEN_1125 ? ~_GEN_1743 & _GEN_109764 : ~(_GEN_110125 & _GEN_1743) & _GEN_109764) : _GEN_109764;
  wire        _GEN_109999 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1744 & _GEN_109765 : _GEN_1125 ? ~_GEN_1744 & _GEN_109765 : ~(_GEN_110125 & _GEN_1744) & _GEN_109765) : _GEN_109765;
  wire        _GEN_110000 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1745 & _GEN_109766 : _GEN_1125 ? ~_GEN_1745 & _GEN_109766 : ~(_GEN_110125 & _GEN_1745) & _GEN_109766) : _GEN_109766;
  wire        _GEN_110001 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1746 & _GEN_109767 : _GEN_1125 ? ~_GEN_1746 & _GEN_109767 : ~(_GEN_110125 & _GEN_1746) & _GEN_109767) : _GEN_109767;
  wire        _GEN_110002 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1747 & _GEN_109768 : _GEN_1125 ? ~_GEN_1747 & _GEN_109768 : ~(_GEN_110125 & _GEN_1747) & _GEN_109768) : _GEN_109768;
  wire        _GEN_110003 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1748 & _GEN_109769 : _GEN_1125 ? ~_GEN_1748 & _GEN_109769 : ~(_GEN_110125 & _GEN_1748) & _GEN_109769) : _GEN_109769;
  wire        _GEN_110004 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1749 & _GEN_109770 : _GEN_1125 ? ~_GEN_1749 & _GEN_109770 : ~(_GEN_110125 & _GEN_1749) & _GEN_109770) : _GEN_109770;
  wire        _GEN_110005 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1750 & _GEN_109771 : _GEN_1125 ? ~_GEN_1750 & _GEN_109771 : ~(_GEN_110125 & _GEN_1750) & _GEN_109771) : _GEN_109771;
  wire        _GEN_110006 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1751 & _GEN_109772 : _GEN_1125 ? ~_GEN_1751 & _GEN_109772 : ~(_GEN_110125 & _GEN_1751) & _GEN_109772) : _GEN_109772;
  wire        _GEN_110007 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1752 & _GEN_109773 : _GEN_1125 ? ~_GEN_1752 & _GEN_109773 : ~(_GEN_110125 & _GEN_1752) & _GEN_109773) : _GEN_109773;
  wire        _GEN_110008 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1753 & _GEN_109774 : _GEN_1125 ? ~_GEN_1753 & _GEN_109774 : ~(_GEN_110125 & _GEN_1753) & _GEN_109774) : _GEN_109774;
  wire        _GEN_110009 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1754 & _GEN_109775 : _GEN_1125 ? ~_GEN_1754 & _GEN_109775 : ~(_GEN_110125 & _GEN_1754) & _GEN_109775) : _GEN_109775;
  wire        _GEN_110010 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1755 & _GEN_109776 : _GEN_1125 ? ~_GEN_1755 & _GEN_109776 : ~(_GEN_110125 & _GEN_1755) & _GEN_109776) : _GEN_109776;
  wire        _GEN_110011 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1756 & _GEN_109777 : _GEN_1125 ? ~_GEN_1756 & _GEN_109777 : ~(_GEN_110125 & _GEN_1756) & _GEN_109777) : _GEN_109777;
  wire        _GEN_110012 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1757 & _GEN_109778 : _GEN_1125 ? ~_GEN_1757 & _GEN_109778 : ~(_GEN_110125 & _GEN_1757) & _GEN_109778) : _GEN_109778;
  wire        _GEN_110013 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1758 & _GEN_109779 : _GEN_1125 ? ~_GEN_1758 & _GEN_109779 : ~(_GEN_110125 & _GEN_1758) & _GEN_109779) : _GEN_109779;
  wire        _GEN_110014 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1759 & _GEN_109780 : _GEN_1125 ? ~_GEN_1759 & _GEN_109780 : ~(_GEN_110125 & _GEN_1759) & _GEN_109780) : _GEN_109780;
  wire        _GEN_110015 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1760 & _GEN_109781 : _GEN_1125 ? ~_GEN_1760 & _GEN_109781 : ~(_GEN_110125 & _GEN_1760) & _GEN_109781) : _GEN_109781;
  wire        _GEN_110016 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1761 & _GEN_109782 : _GEN_1125 ? ~_GEN_1761 & _GEN_109782 : ~(_GEN_110125 & _GEN_1761) & _GEN_109782) : _GEN_109782;
  wire        _GEN_110017 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1762 & _GEN_109783 : _GEN_1125 ? ~_GEN_1762 & _GEN_109783 : ~(_GEN_110125 & _GEN_1762) & _GEN_109783) : _GEN_109783;
  wire        _GEN_110018 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1763 & _GEN_109784 : _GEN_1125 ? ~_GEN_1763 & _GEN_109784 : ~(_GEN_110125 & _GEN_1763) & _GEN_109784) : _GEN_109784;
  wire        _GEN_110019 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1764 & _GEN_109785 : _GEN_1125 ? ~_GEN_1764 & _GEN_109785 : ~(_GEN_110125 & _GEN_1764) & _GEN_109785) : _GEN_109785;
  wire        _GEN_110020 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1765 & _GEN_109786 : _GEN_1125 ? ~_GEN_1765 & _GEN_109786 : ~(_GEN_110125 & _GEN_1765) & _GEN_109786) : _GEN_109786;
  wire        _GEN_110021 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1766 & _GEN_109787 : _GEN_1125 ? ~_GEN_1766 & _GEN_109787 : ~(_GEN_110125 & _GEN_1766) & _GEN_109787) : _GEN_109787;
  wire        _GEN_110022 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1767 & _GEN_109788 : _GEN_1125 ? ~_GEN_1767 & _GEN_109788 : ~(_GEN_110125 & _GEN_1767) & _GEN_109788) : _GEN_109788;
  wire        _GEN_110023 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1768 & _GEN_109789 : _GEN_1125 ? ~_GEN_1768 & _GEN_109789 : ~(_GEN_110125 & _GEN_1768) & _GEN_109789) : _GEN_109789;
  wire        _GEN_110024 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1769 & _GEN_109790 : _GEN_1125 ? ~_GEN_1769 & _GEN_109790 : ~(_GEN_110125 & _GEN_1769) & _GEN_109790) : _GEN_109790;
  wire        _GEN_110025 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1770 & _GEN_109791 : _GEN_1125 ? ~_GEN_1770 & _GEN_109791 : ~(_GEN_110125 & _GEN_1770) & _GEN_109791) : _GEN_109791;
  wire        _GEN_110026 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1771 & _GEN_109792 : _GEN_1125 ? ~_GEN_1771 & _GEN_109792 : ~(_GEN_110125 & _GEN_1771) & _GEN_109792) : _GEN_109792;
  wire        _GEN_110027 = _GEN_1123 ? (_GEN_109960 ? ~_GEN_1772 & _GEN_109793 : _GEN_1125 ? ~_GEN_1772 & _GEN_109793 : ~(_GEN_110125 & _GEN_1772) & _GEN_109793) : _GEN_109793;
  wire        _GEN_110028 = _GEN_1123 ? (_GEN_109960 ? ~(&lcam_ldq_idx_0) & _GEN_109794 : _GEN_1125 ? ~(&lcam_ldq_idx_0) & _GEN_109794 : ~(_GEN_110125 & (&lcam_ldq_idx_0)) & _GEN_109794) : _GEN_109794;
  wire        _GEN_110231 = _GEN_1126 ? (_GEN_110194 ? (|lcam_ldq_idx_1) & _GEN_109997 : _GEN_1128 ? (|lcam_ldq_idx_1) & _GEN_109997 : ~(_GEN_110125 & ~(|lcam_ldq_idx_1)) & _GEN_109997) : _GEN_109997;
  wire        _GEN_110232 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1773 & _GEN_109998 : _GEN_1128 ? ~_GEN_1773 & _GEN_109998 : ~(_GEN_110125 & _GEN_1773) & _GEN_109998) : _GEN_109998;
  wire        _GEN_110233 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1774 & _GEN_109999 : _GEN_1128 ? ~_GEN_1774 & _GEN_109999 : ~(_GEN_110125 & _GEN_1774) & _GEN_109999) : _GEN_109999;
  wire        _GEN_110234 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1775 & _GEN_110000 : _GEN_1128 ? ~_GEN_1775 & _GEN_110000 : ~(_GEN_110125 & _GEN_1775) & _GEN_110000) : _GEN_110000;
  wire        _GEN_110235 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1776 & _GEN_110001 : _GEN_1128 ? ~_GEN_1776 & _GEN_110001 : ~(_GEN_110125 & _GEN_1776) & _GEN_110001) : _GEN_110001;
  wire        _GEN_110236 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1777 & _GEN_110002 : _GEN_1128 ? ~_GEN_1777 & _GEN_110002 : ~(_GEN_110125 & _GEN_1777) & _GEN_110002) : _GEN_110002;
  wire        _GEN_110237 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1778 & _GEN_110003 : _GEN_1128 ? ~_GEN_1778 & _GEN_110003 : ~(_GEN_110125 & _GEN_1778) & _GEN_110003) : _GEN_110003;
  wire        _GEN_110238 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1779 & _GEN_110004 : _GEN_1128 ? ~_GEN_1779 & _GEN_110004 : ~(_GEN_110125 & _GEN_1779) & _GEN_110004) : _GEN_110004;
  wire        _GEN_110239 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1780 & _GEN_110005 : _GEN_1128 ? ~_GEN_1780 & _GEN_110005 : ~(_GEN_110125 & _GEN_1780) & _GEN_110005) : _GEN_110005;
  wire        _GEN_110240 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1781 & _GEN_110006 : _GEN_1128 ? ~_GEN_1781 & _GEN_110006 : ~(_GEN_110125 & _GEN_1781) & _GEN_110006) : _GEN_110006;
  wire        _GEN_110241 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1782 & _GEN_110007 : _GEN_1128 ? ~_GEN_1782 & _GEN_110007 : ~(_GEN_110125 & _GEN_1782) & _GEN_110007) : _GEN_110007;
  wire        _GEN_110242 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1783 & _GEN_110008 : _GEN_1128 ? ~_GEN_1783 & _GEN_110008 : ~(_GEN_110125 & _GEN_1783) & _GEN_110008) : _GEN_110008;
  wire        _GEN_110243 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1784 & _GEN_110009 : _GEN_1128 ? ~_GEN_1784 & _GEN_110009 : ~(_GEN_110125 & _GEN_1784) & _GEN_110009) : _GEN_110009;
  wire        _GEN_110244 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1785 & _GEN_110010 : _GEN_1128 ? ~_GEN_1785 & _GEN_110010 : ~(_GEN_110125 & _GEN_1785) & _GEN_110010) : _GEN_110010;
  wire        _GEN_110245 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1786 & _GEN_110011 : _GEN_1128 ? ~_GEN_1786 & _GEN_110011 : ~(_GEN_110125 & _GEN_1786) & _GEN_110011) : _GEN_110011;
  wire        _GEN_110246 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1787 & _GEN_110012 : _GEN_1128 ? ~_GEN_1787 & _GEN_110012 : ~(_GEN_110125 & _GEN_1787) & _GEN_110012) : _GEN_110012;
  wire        _GEN_110247 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1788 & _GEN_110013 : _GEN_1128 ? ~_GEN_1788 & _GEN_110013 : ~(_GEN_110125 & _GEN_1788) & _GEN_110013) : _GEN_110013;
  wire        _GEN_110248 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1789 & _GEN_110014 : _GEN_1128 ? ~_GEN_1789 & _GEN_110014 : ~(_GEN_110125 & _GEN_1789) & _GEN_110014) : _GEN_110014;
  wire        _GEN_110249 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1790 & _GEN_110015 : _GEN_1128 ? ~_GEN_1790 & _GEN_110015 : ~(_GEN_110125 & _GEN_1790) & _GEN_110015) : _GEN_110015;
  wire        _GEN_110250 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1791 & _GEN_110016 : _GEN_1128 ? ~_GEN_1791 & _GEN_110016 : ~(_GEN_110125 & _GEN_1791) & _GEN_110016) : _GEN_110016;
  wire        _GEN_110251 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1792 & _GEN_110017 : _GEN_1128 ? ~_GEN_1792 & _GEN_110017 : ~(_GEN_110125 & _GEN_1792) & _GEN_110017) : _GEN_110017;
  wire        _GEN_110252 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1793 & _GEN_110018 : _GEN_1128 ? ~_GEN_1793 & _GEN_110018 : ~(_GEN_110125 & _GEN_1793) & _GEN_110018) : _GEN_110018;
  wire        _GEN_110253 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1794 & _GEN_110019 : _GEN_1128 ? ~_GEN_1794 & _GEN_110019 : ~(_GEN_110125 & _GEN_1794) & _GEN_110019) : _GEN_110019;
  wire        _GEN_110254 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1795 & _GEN_110020 : _GEN_1128 ? ~_GEN_1795 & _GEN_110020 : ~(_GEN_110125 & _GEN_1795) & _GEN_110020) : _GEN_110020;
  wire        _GEN_110255 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1796 & _GEN_110021 : _GEN_1128 ? ~_GEN_1796 & _GEN_110021 : ~(_GEN_110125 & _GEN_1796) & _GEN_110021) : _GEN_110021;
  wire        _GEN_110256 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1797 & _GEN_110022 : _GEN_1128 ? ~_GEN_1797 & _GEN_110022 : ~(_GEN_110125 & _GEN_1797) & _GEN_110022) : _GEN_110022;
  wire        _GEN_110257 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1798 & _GEN_110023 : _GEN_1128 ? ~_GEN_1798 & _GEN_110023 : ~(_GEN_110125 & _GEN_1798) & _GEN_110023) : _GEN_110023;
  wire        _GEN_110258 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1799 & _GEN_110024 : _GEN_1128 ? ~_GEN_1799 & _GEN_110024 : ~(_GEN_110125 & _GEN_1799) & _GEN_110024) : _GEN_110024;
  wire        _GEN_110259 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1800 & _GEN_110025 : _GEN_1128 ? ~_GEN_1800 & _GEN_110025 : ~(_GEN_110125 & _GEN_1800) & _GEN_110025) : _GEN_110025;
  wire        _GEN_110260 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1801 & _GEN_110026 : _GEN_1128 ? ~_GEN_1801 & _GEN_110026 : ~(_GEN_110125 & _GEN_1801) & _GEN_110026) : _GEN_110026;
  wire        _GEN_110261 = _GEN_1126 ? (_GEN_110194 ? ~_GEN_1802 & _GEN_110027 : _GEN_1128 ? ~_GEN_1802 & _GEN_110027 : ~(_GEN_110125 & _GEN_1802) & _GEN_110027) : _GEN_110027;
  wire        _GEN_110262 = _GEN_1126 ? (_GEN_110194 ? ~(&lcam_ldq_idx_1) & _GEN_110028 : _GEN_1128 ? ~(&lcam_ldq_idx_1) & _GEN_110028 : ~(_GEN_110125 & (&lcam_ldq_idx_1)) & _GEN_110028) : _GEN_110028;
  wire        _GEN_110465 = _GEN_1129 ? (_GEN_110428 ? (|lcam_ldq_idx_0) & _GEN_110231 : _GEN_1131 ? (|lcam_ldq_idx_0) & _GEN_110231 : ~(_GEN_110593 & ~(|lcam_ldq_idx_0)) & _GEN_110231) : _GEN_110231;
  wire        _GEN_110466 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1743 & _GEN_110232 : _GEN_1131 ? ~_GEN_1743 & _GEN_110232 : ~(_GEN_110593 & _GEN_1743) & _GEN_110232) : _GEN_110232;
  wire        _GEN_110467 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1744 & _GEN_110233 : _GEN_1131 ? ~_GEN_1744 & _GEN_110233 : ~(_GEN_110593 & _GEN_1744) & _GEN_110233) : _GEN_110233;
  wire        _GEN_110468 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1745 & _GEN_110234 : _GEN_1131 ? ~_GEN_1745 & _GEN_110234 : ~(_GEN_110593 & _GEN_1745) & _GEN_110234) : _GEN_110234;
  wire        _GEN_110469 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1746 & _GEN_110235 : _GEN_1131 ? ~_GEN_1746 & _GEN_110235 : ~(_GEN_110593 & _GEN_1746) & _GEN_110235) : _GEN_110235;
  wire        _GEN_110470 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1747 & _GEN_110236 : _GEN_1131 ? ~_GEN_1747 & _GEN_110236 : ~(_GEN_110593 & _GEN_1747) & _GEN_110236) : _GEN_110236;
  wire        _GEN_110471 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1748 & _GEN_110237 : _GEN_1131 ? ~_GEN_1748 & _GEN_110237 : ~(_GEN_110593 & _GEN_1748) & _GEN_110237) : _GEN_110237;
  wire        _GEN_110472 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1749 & _GEN_110238 : _GEN_1131 ? ~_GEN_1749 & _GEN_110238 : ~(_GEN_110593 & _GEN_1749) & _GEN_110238) : _GEN_110238;
  wire        _GEN_110473 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1750 & _GEN_110239 : _GEN_1131 ? ~_GEN_1750 & _GEN_110239 : ~(_GEN_110593 & _GEN_1750) & _GEN_110239) : _GEN_110239;
  wire        _GEN_110474 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1751 & _GEN_110240 : _GEN_1131 ? ~_GEN_1751 & _GEN_110240 : ~(_GEN_110593 & _GEN_1751) & _GEN_110240) : _GEN_110240;
  wire        _GEN_110475 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1752 & _GEN_110241 : _GEN_1131 ? ~_GEN_1752 & _GEN_110241 : ~(_GEN_110593 & _GEN_1752) & _GEN_110241) : _GEN_110241;
  wire        _GEN_110476 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1753 & _GEN_110242 : _GEN_1131 ? ~_GEN_1753 & _GEN_110242 : ~(_GEN_110593 & _GEN_1753) & _GEN_110242) : _GEN_110242;
  wire        _GEN_110477 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1754 & _GEN_110243 : _GEN_1131 ? ~_GEN_1754 & _GEN_110243 : ~(_GEN_110593 & _GEN_1754) & _GEN_110243) : _GEN_110243;
  wire        _GEN_110478 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1755 & _GEN_110244 : _GEN_1131 ? ~_GEN_1755 & _GEN_110244 : ~(_GEN_110593 & _GEN_1755) & _GEN_110244) : _GEN_110244;
  wire        _GEN_110479 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1756 & _GEN_110245 : _GEN_1131 ? ~_GEN_1756 & _GEN_110245 : ~(_GEN_110593 & _GEN_1756) & _GEN_110245) : _GEN_110245;
  wire        _GEN_110480 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1757 & _GEN_110246 : _GEN_1131 ? ~_GEN_1757 & _GEN_110246 : ~(_GEN_110593 & _GEN_1757) & _GEN_110246) : _GEN_110246;
  wire        _GEN_110481 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1758 & _GEN_110247 : _GEN_1131 ? ~_GEN_1758 & _GEN_110247 : ~(_GEN_110593 & _GEN_1758) & _GEN_110247) : _GEN_110247;
  wire        _GEN_110482 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1759 & _GEN_110248 : _GEN_1131 ? ~_GEN_1759 & _GEN_110248 : ~(_GEN_110593 & _GEN_1759) & _GEN_110248) : _GEN_110248;
  wire        _GEN_110483 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1760 & _GEN_110249 : _GEN_1131 ? ~_GEN_1760 & _GEN_110249 : ~(_GEN_110593 & _GEN_1760) & _GEN_110249) : _GEN_110249;
  wire        _GEN_110484 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1761 & _GEN_110250 : _GEN_1131 ? ~_GEN_1761 & _GEN_110250 : ~(_GEN_110593 & _GEN_1761) & _GEN_110250) : _GEN_110250;
  wire        _GEN_110485 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1762 & _GEN_110251 : _GEN_1131 ? ~_GEN_1762 & _GEN_110251 : ~(_GEN_110593 & _GEN_1762) & _GEN_110251) : _GEN_110251;
  wire        _GEN_110486 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1763 & _GEN_110252 : _GEN_1131 ? ~_GEN_1763 & _GEN_110252 : ~(_GEN_110593 & _GEN_1763) & _GEN_110252) : _GEN_110252;
  wire        _GEN_110487 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1764 & _GEN_110253 : _GEN_1131 ? ~_GEN_1764 & _GEN_110253 : ~(_GEN_110593 & _GEN_1764) & _GEN_110253) : _GEN_110253;
  wire        _GEN_110488 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1765 & _GEN_110254 : _GEN_1131 ? ~_GEN_1765 & _GEN_110254 : ~(_GEN_110593 & _GEN_1765) & _GEN_110254) : _GEN_110254;
  wire        _GEN_110489 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1766 & _GEN_110255 : _GEN_1131 ? ~_GEN_1766 & _GEN_110255 : ~(_GEN_110593 & _GEN_1766) & _GEN_110255) : _GEN_110255;
  wire        _GEN_110490 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1767 & _GEN_110256 : _GEN_1131 ? ~_GEN_1767 & _GEN_110256 : ~(_GEN_110593 & _GEN_1767) & _GEN_110256) : _GEN_110256;
  wire        _GEN_110491 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1768 & _GEN_110257 : _GEN_1131 ? ~_GEN_1768 & _GEN_110257 : ~(_GEN_110593 & _GEN_1768) & _GEN_110257) : _GEN_110257;
  wire        _GEN_110492 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1769 & _GEN_110258 : _GEN_1131 ? ~_GEN_1769 & _GEN_110258 : ~(_GEN_110593 & _GEN_1769) & _GEN_110258) : _GEN_110258;
  wire        _GEN_110493 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1770 & _GEN_110259 : _GEN_1131 ? ~_GEN_1770 & _GEN_110259 : ~(_GEN_110593 & _GEN_1770) & _GEN_110259) : _GEN_110259;
  wire        _GEN_110494 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1771 & _GEN_110260 : _GEN_1131 ? ~_GEN_1771 & _GEN_110260 : ~(_GEN_110593 & _GEN_1771) & _GEN_110260) : _GEN_110260;
  wire        _GEN_110495 = _GEN_1129 ? (_GEN_110428 ? ~_GEN_1772 & _GEN_110261 : _GEN_1131 ? ~_GEN_1772 & _GEN_110261 : ~(_GEN_110593 & _GEN_1772) & _GEN_110261) : _GEN_110261;
  wire        _GEN_110496 = _GEN_1129 ? (_GEN_110428 ? ~(&lcam_ldq_idx_0) & _GEN_110262 : _GEN_1131 ? ~(&lcam_ldq_idx_0) & _GEN_110262 : ~(_GEN_110593 & (&lcam_ldq_idx_0)) & _GEN_110262) : _GEN_110262;
  wire        _GEN_110699 = _GEN_1132 ? (_GEN_110662 ? (|lcam_ldq_idx_1) & _GEN_110465 : _GEN_1134 ? (|lcam_ldq_idx_1) & _GEN_110465 : ~(_GEN_110593 & ~(|lcam_ldq_idx_1)) & _GEN_110465) : _GEN_110465;
  wire        _GEN_110700 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1773 & _GEN_110466 : _GEN_1134 ? ~_GEN_1773 & _GEN_110466 : ~(_GEN_110593 & _GEN_1773) & _GEN_110466) : _GEN_110466;
  wire        _GEN_110701 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1774 & _GEN_110467 : _GEN_1134 ? ~_GEN_1774 & _GEN_110467 : ~(_GEN_110593 & _GEN_1774) & _GEN_110467) : _GEN_110467;
  wire        _GEN_110702 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1775 & _GEN_110468 : _GEN_1134 ? ~_GEN_1775 & _GEN_110468 : ~(_GEN_110593 & _GEN_1775) & _GEN_110468) : _GEN_110468;
  wire        _GEN_110703 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1776 & _GEN_110469 : _GEN_1134 ? ~_GEN_1776 & _GEN_110469 : ~(_GEN_110593 & _GEN_1776) & _GEN_110469) : _GEN_110469;
  wire        _GEN_110704 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1777 & _GEN_110470 : _GEN_1134 ? ~_GEN_1777 & _GEN_110470 : ~(_GEN_110593 & _GEN_1777) & _GEN_110470) : _GEN_110470;
  wire        _GEN_110705 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1778 & _GEN_110471 : _GEN_1134 ? ~_GEN_1778 & _GEN_110471 : ~(_GEN_110593 & _GEN_1778) & _GEN_110471) : _GEN_110471;
  wire        _GEN_110706 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1779 & _GEN_110472 : _GEN_1134 ? ~_GEN_1779 & _GEN_110472 : ~(_GEN_110593 & _GEN_1779) & _GEN_110472) : _GEN_110472;
  wire        _GEN_110707 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1780 & _GEN_110473 : _GEN_1134 ? ~_GEN_1780 & _GEN_110473 : ~(_GEN_110593 & _GEN_1780) & _GEN_110473) : _GEN_110473;
  wire        _GEN_110708 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1781 & _GEN_110474 : _GEN_1134 ? ~_GEN_1781 & _GEN_110474 : ~(_GEN_110593 & _GEN_1781) & _GEN_110474) : _GEN_110474;
  wire        _GEN_110709 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1782 & _GEN_110475 : _GEN_1134 ? ~_GEN_1782 & _GEN_110475 : ~(_GEN_110593 & _GEN_1782) & _GEN_110475) : _GEN_110475;
  wire        _GEN_110710 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1783 & _GEN_110476 : _GEN_1134 ? ~_GEN_1783 & _GEN_110476 : ~(_GEN_110593 & _GEN_1783) & _GEN_110476) : _GEN_110476;
  wire        _GEN_110711 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1784 & _GEN_110477 : _GEN_1134 ? ~_GEN_1784 & _GEN_110477 : ~(_GEN_110593 & _GEN_1784) & _GEN_110477) : _GEN_110477;
  wire        _GEN_110712 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1785 & _GEN_110478 : _GEN_1134 ? ~_GEN_1785 & _GEN_110478 : ~(_GEN_110593 & _GEN_1785) & _GEN_110478) : _GEN_110478;
  wire        _GEN_110713 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1786 & _GEN_110479 : _GEN_1134 ? ~_GEN_1786 & _GEN_110479 : ~(_GEN_110593 & _GEN_1786) & _GEN_110479) : _GEN_110479;
  wire        _GEN_110714 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1787 & _GEN_110480 : _GEN_1134 ? ~_GEN_1787 & _GEN_110480 : ~(_GEN_110593 & _GEN_1787) & _GEN_110480) : _GEN_110480;
  wire        _GEN_110715 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1788 & _GEN_110481 : _GEN_1134 ? ~_GEN_1788 & _GEN_110481 : ~(_GEN_110593 & _GEN_1788) & _GEN_110481) : _GEN_110481;
  wire        _GEN_110716 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1789 & _GEN_110482 : _GEN_1134 ? ~_GEN_1789 & _GEN_110482 : ~(_GEN_110593 & _GEN_1789) & _GEN_110482) : _GEN_110482;
  wire        _GEN_110717 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1790 & _GEN_110483 : _GEN_1134 ? ~_GEN_1790 & _GEN_110483 : ~(_GEN_110593 & _GEN_1790) & _GEN_110483) : _GEN_110483;
  wire        _GEN_110718 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1791 & _GEN_110484 : _GEN_1134 ? ~_GEN_1791 & _GEN_110484 : ~(_GEN_110593 & _GEN_1791) & _GEN_110484) : _GEN_110484;
  wire        _GEN_110719 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1792 & _GEN_110485 : _GEN_1134 ? ~_GEN_1792 & _GEN_110485 : ~(_GEN_110593 & _GEN_1792) & _GEN_110485) : _GEN_110485;
  wire        _GEN_110720 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1793 & _GEN_110486 : _GEN_1134 ? ~_GEN_1793 & _GEN_110486 : ~(_GEN_110593 & _GEN_1793) & _GEN_110486) : _GEN_110486;
  wire        _GEN_110721 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1794 & _GEN_110487 : _GEN_1134 ? ~_GEN_1794 & _GEN_110487 : ~(_GEN_110593 & _GEN_1794) & _GEN_110487) : _GEN_110487;
  wire        _GEN_110722 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1795 & _GEN_110488 : _GEN_1134 ? ~_GEN_1795 & _GEN_110488 : ~(_GEN_110593 & _GEN_1795) & _GEN_110488) : _GEN_110488;
  wire        _GEN_110723 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1796 & _GEN_110489 : _GEN_1134 ? ~_GEN_1796 & _GEN_110489 : ~(_GEN_110593 & _GEN_1796) & _GEN_110489) : _GEN_110489;
  wire        _GEN_110724 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1797 & _GEN_110490 : _GEN_1134 ? ~_GEN_1797 & _GEN_110490 : ~(_GEN_110593 & _GEN_1797) & _GEN_110490) : _GEN_110490;
  wire        _GEN_110725 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1798 & _GEN_110491 : _GEN_1134 ? ~_GEN_1798 & _GEN_110491 : ~(_GEN_110593 & _GEN_1798) & _GEN_110491) : _GEN_110491;
  wire        _GEN_110726 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1799 & _GEN_110492 : _GEN_1134 ? ~_GEN_1799 & _GEN_110492 : ~(_GEN_110593 & _GEN_1799) & _GEN_110492) : _GEN_110492;
  wire        _GEN_110727 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1800 & _GEN_110493 : _GEN_1134 ? ~_GEN_1800 & _GEN_110493 : ~(_GEN_110593 & _GEN_1800) & _GEN_110493) : _GEN_110493;
  wire        _GEN_110728 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1801 & _GEN_110494 : _GEN_1134 ? ~_GEN_1801 & _GEN_110494 : ~(_GEN_110593 & _GEN_1801) & _GEN_110494) : _GEN_110494;
  wire        _GEN_110729 = _GEN_1132 ? (_GEN_110662 ? ~_GEN_1802 & _GEN_110495 : _GEN_1134 ? ~_GEN_1802 & _GEN_110495 : ~(_GEN_110593 & _GEN_1802) & _GEN_110495) : _GEN_110495;
  wire        _GEN_110730 = _GEN_1132 ? (_GEN_110662 ? ~(&lcam_ldq_idx_1) & _GEN_110496 : _GEN_1134 ? ~(&lcam_ldq_idx_1) & _GEN_110496 : ~(_GEN_110593 & (&lcam_ldq_idx_1)) & _GEN_110496) : _GEN_110496;
  wire        _GEN_110933 = _GEN_1135 ? (_GEN_110896 ? (|lcam_ldq_idx_0) & _GEN_110699 : _GEN_1137 ? (|lcam_ldq_idx_0) & _GEN_110699 : ~(_GEN_111061 & ~(|lcam_ldq_idx_0)) & _GEN_110699) : _GEN_110699;
  wire        _GEN_110934 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1743 & _GEN_110700 : _GEN_1137 ? ~_GEN_1743 & _GEN_110700 : ~(_GEN_111061 & _GEN_1743) & _GEN_110700) : _GEN_110700;
  wire        _GEN_110935 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1744 & _GEN_110701 : _GEN_1137 ? ~_GEN_1744 & _GEN_110701 : ~(_GEN_111061 & _GEN_1744) & _GEN_110701) : _GEN_110701;
  wire        _GEN_110936 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1745 & _GEN_110702 : _GEN_1137 ? ~_GEN_1745 & _GEN_110702 : ~(_GEN_111061 & _GEN_1745) & _GEN_110702) : _GEN_110702;
  wire        _GEN_110937 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1746 & _GEN_110703 : _GEN_1137 ? ~_GEN_1746 & _GEN_110703 : ~(_GEN_111061 & _GEN_1746) & _GEN_110703) : _GEN_110703;
  wire        _GEN_110938 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1747 & _GEN_110704 : _GEN_1137 ? ~_GEN_1747 & _GEN_110704 : ~(_GEN_111061 & _GEN_1747) & _GEN_110704) : _GEN_110704;
  wire        _GEN_110939 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1748 & _GEN_110705 : _GEN_1137 ? ~_GEN_1748 & _GEN_110705 : ~(_GEN_111061 & _GEN_1748) & _GEN_110705) : _GEN_110705;
  wire        _GEN_110940 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1749 & _GEN_110706 : _GEN_1137 ? ~_GEN_1749 & _GEN_110706 : ~(_GEN_111061 & _GEN_1749) & _GEN_110706) : _GEN_110706;
  wire        _GEN_110941 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1750 & _GEN_110707 : _GEN_1137 ? ~_GEN_1750 & _GEN_110707 : ~(_GEN_111061 & _GEN_1750) & _GEN_110707) : _GEN_110707;
  wire        _GEN_110942 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1751 & _GEN_110708 : _GEN_1137 ? ~_GEN_1751 & _GEN_110708 : ~(_GEN_111061 & _GEN_1751) & _GEN_110708) : _GEN_110708;
  wire        _GEN_110943 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1752 & _GEN_110709 : _GEN_1137 ? ~_GEN_1752 & _GEN_110709 : ~(_GEN_111061 & _GEN_1752) & _GEN_110709) : _GEN_110709;
  wire        _GEN_110944 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1753 & _GEN_110710 : _GEN_1137 ? ~_GEN_1753 & _GEN_110710 : ~(_GEN_111061 & _GEN_1753) & _GEN_110710) : _GEN_110710;
  wire        _GEN_110945 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1754 & _GEN_110711 : _GEN_1137 ? ~_GEN_1754 & _GEN_110711 : ~(_GEN_111061 & _GEN_1754) & _GEN_110711) : _GEN_110711;
  wire        _GEN_110946 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1755 & _GEN_110712 : _GEN_1137 ? ~_GEN_1755 & _GEN_110712 : ~(_GEN_111061 & _GEN_1755) & _GEN_110712) : _GEN_110712;
  wire        _GEN_110947 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1756 & _GEN_110713 : _GEN_1137 ? ~_GEN_1756 & _GEN_110713 : ~(_GEN_111061 & _GEN_1756) & _GEN_110713) : _GEN_110713;
  wire        _GEN_110948 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1757 & _GEN_110714 : _GEN_1137 ? ~_GEN_1757 & _GEN_110714 : ~(_GEN_111061 & _GEN_1757) & _GEN_110714) : _GEN_110714;
  wire        _GEN_110949 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1758 & _GEN_110715 : _GEN_1137 ? ~_GEN_1758 & _GEN_110715 : ~(_GEN_111061 & _GEN_1758) & _GEN_110715) : _GEN_110715;
  wire        _GEN_110950 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1759 & _GEN_110716 : _GEN_1137 ? ~_GEN_1759 & _GEN_110716 : ~(_GEN_111061 & _GEN_1759) & _GEN_110716) : _GEN_110716;
  wire        _GEN_110951 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1760 & _GEN_110717 : _GEN_1137 ? ~_GEN_1760 & _GEN_110717 : ~(_GEN_111061 & _GEN_1760) & _GEN_110717) : _GEN_110717;
  wire        _GEN_110952 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1761 & _GEN_110718 : _GEN_1137 ? ~_GEN_1761 & _GEN_110718 : ~(_GEN_111061 & _GEN_1761) & _GEN_110718) : _GEN_110718;
  wire        _GEN_110953 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1762 & _GEN_110719 : _GEN_1137 ? ~_GEN_1762 & _GEN_110719 : ~(_GEN_111061 & _GEN_1762) & _GEN_110719) : _GEN_110719;
  wire        _GEN_110954 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1763 & _GEN_110720 : _GEN_1137 ? ~_GEN_1763 & _GEN_110720 : ~(_GEN_111061 & _GEN_1763) & _GEN_110720) : _GEN_110720;
  wire        _GEN_110955 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1764 & _GEN_110721 : _GEN_1137 ? ~_GEN_1764 & _GEN_110721 : ~(_GEN_111061 & _GEN_1764) & _GEN_110721) : _GEN_110721;
  wire        _GEN_110956 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1765 & _GEN_110722 : _GEN_1137 ? ~_GEN_1765 & _GEN_110722 : ~(_GEN_111061 & _GEN_1765) & _GEN_110722) : _GEN_110722;
  wire        _GEN_110957 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1766 & _GEN_110723 : _GEN_1137 ? ~_GEN_1766 & _GEN_110723 : ~(_GEN_111061 & _GEN_1766) & _GEN_110723) : _GEN_110723;
  wire        _GEN_110958 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1767 & _GEN_110724 : _GEN_1137 ? ~_GEN_1767 & _GEN_110724 : ~(_GEN_111061 & _GEN_1767) & _GEN_110724) : _GEN_110724;
  wire        _GEN_110959 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1768 & _GEN_110725 : _GEN_1137 ? ~_GEN_1768 & _GEN_110725 : ~(_GEN_111061 & _GEN_1768) & _GEN_110725) : _GEN_110725;
  wire        _GEN_110960 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1769 & _GEN_110726 : _GEN_1137 ? ~_GEN_1769 & _GEN_110726 : ~(_GEN_111061 & _GEN_1769) & _GEN_110726) : _GEN_110726;
  wire        _GEN_110961 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1770 & _GEN_110727 : _GEN_1137 ? ~_GEN_1770 & _GEN_110727 : ~(_GEN_111061 & _GEN_1770) & _GEN_110727) : _GEN_110727;
  wire        _GEN_110962 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1771 & _GEN_110728 : _GEN_1137 ? ~_GEN_1771 & _GEN_110728 : ~(_GEN_111061 & _GEN_1771) & _GEN_110728) : _GEN_110728;
  wire        _GEN_110963 = _GEN_1135 ? (_GEN_110896 ? ~_GEN_1772 & _GEN_110729 : _GEN_1137 ? ~_GEN_1772 & _GEN_110729 : ~(_GEN_111061 & _GEN_1772) & _GEN_110729) : _GEN_110729;
  wire        _GEN_110964 = _GEN_1135 ? (_GEN_110896 ? ~(&lcam_ldq_idx_0) & _GEN_110730 : _GEN_1137 ? ~(&lcam_ldq_idx_0) & _GEN_110730 : ~(_GEN_111061 & (&lcam_ldq_idx_0)) & _GEN_110730) : _GEN_110730;
  wire        _GEN_111167 = _GEN_1138 ? (_GEN_111130 ? (|lcam_ldq_idx_1) & _GEN_110933 : _GEN_1140 ? (|lcam_ldq_idx_1) & _GEN_110933 : ~(_GEN_111061 & ~(|lcam_ldq_idx_1)) & _GEN_110933) : _GEN_110933;
  wire        _GEN_111168 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1773 & _GEN_110934 : _GEN_1140 ? ~_GEN_1773 & _GEN_110934 : ~(_GEN_111061 & _GEN_1773) & _GEN_110934) : _GEN_110934;
  wire        _GEN_111169 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1774 & _GEN_110935 : _GEN_1140 ? ~_GEN_1774 & _GEN_110935 : ~(_GEN_111061 & _GEN_1774) & _GEN_110935) : _GEN_110935;
  wire        _GEN_111170 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1775 & _GEN_110936 : _GEN_1140 ? ~_GEN_1775 & _GEN_110936 : ~(_GEN_111061 & _GEN_1775) & _GEN_110936) : _GEN_110936;
  wire        _GEN_111171 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1776 & _GEN_110937 : _GEN_1140 ? ~_GEN_1776 & _GEN_110937 : ~(_GEN_111061 & _GEN_1776) & _GEN_110937) : _GEN_110937;
  wire        _GEN_111172 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1777 & _GEN_110938 : _GEN_1140 ? ~_GEN_1777 & _GEN_110938 : ~(_GEN_111061 & _GEN_1777) & _GEN_110938) : _GEN_110938;
  wire        _GEN_111173 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1778 & _GEN_110939 : _GEN_1140 ? ~_GEN_1778 & _GEN_110939 : ~(_GEN_111061 & _GEN_1778) & _GEN_110939) : _GEN_110939;
  wire        _GEN_111174 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1779 & _GEN_110940 : _GEN_1140 ? ~_GEN_1779 & _GEN_110940 : ~(_GEN_111061 & _GEN_1779) & _GEN_110940) : _GEN_110940;
  wire        _GEN_111175 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1780 & _GEN_110941 : _GEN_1140 ? ~_GEN_1780 & _GEN_110941 : ~(_GEN_111061 & _GEN_1780) & _GEN_110941) : _GEN_110941;
  wire        _GEN_111176 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1781 & _GEN_110942 : _GEN_1140 ? ~_GEN_1781 & _GEN_110942 : ~(_GEN_111061 & _GEN_1781) & _GEN_110942) : _GEN_110942;
  wire        _GEN_111177 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1782 & _GEN_110943 : _GEN_1140 ? ~_GEN_1782 & _GEN_110943 : ~(_GEN_111061 & _GEN_1782) & _GEN_110943) : _GEN_110943;
  wire        _GEN_111178 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1783 & _GEN_110944 : _GEN_1140 ? ~_GEN_1783 & _GEN_110944 : ~(_GEN_111061 & _GEN_1783) & _GEN_110944) : _GEN_110944;
  wire        _GEN_111179 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1784 & _GEN_110945 : _GEN_1140 ? ~_GEN_1784 & _GEN_110945 : ~(_GEN_111061 & _GEN_1784) & _GEN_110945) : _GEN_110945;
  wire        _GEN_111180 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1785 & _GEN_110946 : _GEN_1140 ? ~_GEN_1785 & _GEN_110946 : ~(_GEN_111061 & _GEN_1785) & _GEN_110946) : _GEN_110946;
  wire        _GEN_111181 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1786 & _GEN_110947 : _GEN_1140 ? ~_GEN_1786 & _GEN_110947 : ~(_GEN_111061 & _GEN_1786) & _GEN_110947) : _GEN_110947;
  wire        _GEN_111182 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1787 & _GEN_110948 : _GEN_1140 ? ~_GEN_1787 & _GEN_110948 : ~(_GEN_111061 & _GEN_1787) & _GEN_110948) : _GEN_110948;
  wire        _GEN_111183 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1788 & _GEN_110949 : _GEN_1140 ? ~_GEN_1788 & _GEN_110949 : ~(_GEN_111061 & _GEN_1788) & _GEN_110949) : _GEN_110949;
  wire        _GEN_111184 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1789 & _GEN_110950 : _GEN_1140 ? ~_GEN_1789 & _GEN_110950 : ~(_GEN_111061 & _GEN_1789) & _GEN_110950) : _GEN_110950;
  wire        _GEN_111185 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1790 & _GEN_110951 : _GEN_1140 ? ~_GEN_1790 & _GEN_110951 : ~(_GEN_111061 & _GEN_1790) & _GEN_110951) : _GEN_110951;
  wire        _GEN_111186 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1791 & _GEN_110952 : _GEN_1140 ? ~_GEN_1791 & _GEN_110952 : ~(_GEN_111061 & _GEN_1791) & _GEN_110952) : _GEN_110952;
  wire        _GEN_111187 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1792 & _GEN_110953 : _GEN_1140 ? ~_GEN_1792 & _GEN_110953 : ~(_GEN_111061 & _GEN_1792) & _GEN_110953) : _GEN_110953;
  wire        _GEN_111188 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1793 & _GEN_110954 : _GEN_1140 ? ~_GEN_1793 & _GEN_110954 : ~(_GEN_111061 & _GEN_1793) & _GEN_110954) : _GEN_110954;
  wire        _GEN_111189 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1794 & _GEN_110955 : _GEN_1140 ? ~_GEN_1794 & _GEN_110955 : ~(_GEN_111061 & _GEN_1794) & _GEN_110955) : _GEN_110955;
  wire        _GEN_111190 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1795 & _GEN_110956 : _GEN_1140 ? ~_GEN_1795 & _GEN_110956 : ~(_GEN_111061 & _GEN_1795) & _GEN_110956) : _GEN_110956;
  wire        _GEN_111191 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1796 & _GEN_110957 : _GEN_1140 ? ~_GEN_1796 & _GEN_110957 : ~(_GEN_111061 & _GEN_1796) & _GEN_110957) : _GEN_110957;
  wire        _GEN_111192 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1797 & _GEN_110958 : _GEN_1140 ? ~_GEN_1797 & _GEN_110958 : ~(_GEN_111061 & _GEN_1797) & _GEN_110958) : _GEN_110958;
  wire        _GEN_111193 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1798 & _GEN_110959 : _GEN_1140 ? ~_GEN_1798 & _GEN_110959 : ~(_GEN_111061 & _GEN_1798) & _GEN_110959) : _GEN_110959;
  wire        _GEN_111194 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1799 & _GEN_110960 : _GEN_1140 ? ~_GEN_1799 & _GEN_110960 : ~(_GEN_111061 & _GEN_1799) & _GEN_110960) : _GEN_110960;
  wire        _GEN_111195 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1800 & _GEN_110961 : _GEN_1140 ? ~_GEN_1800 & _GEN_110961 : ~(_GEN_111061 & _GEN_1800) & _GEN_110961) : _GEN_110961;
  wire        _GEN_111196 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1801 & _GEN_110962 : _GEN_1140 ? ~_GEN_1801 & _GEN_110962 : ~(_GEN_111061 & _GEN_1801) & _GEN_110962) : _GEN_110962;
  wire        _GEN_111197 = _GEN_1138 ? (_GEN_111130 ? ~_GEN_1802 & _GEN_110963 : _GEN_1140 ? ~_GEN_1802 & _GEN_110963 : ~(_GEN_111061 & _GEN_1802) & _GEN_110963) : _GEN_110963;
  wire        _GEN_111198 = _GEN_1138 ? (_GEN_111130 ? ~(&lcam_ldq_idx_1) & _GEN_110964 : _GEN_1140 ? ~(&lcam_ldq_idx_1) & _GEN_110964 : ~(_GEN_111061 & (&lcam_ldq_idx_1)) & _GEN_110964) : _GEN_110964;
  wire        _GEN_111401 = _GEN_1141 ? (_GEN_111364 ? (|lcam_ldq_idx_0) & _GEN_111167 : _GEN_1143 ? (|lcam_ldq_idx_0) & _GEN_111167 : ~(_GEN_111529 & ~(|lcam_ldq_idx_0)) & _GEN_111167) : _GEN_111167;
  wire        _GEN_111402 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1743 & _GEN_111168 : _GEN_1143 ? ~_GEN_1743 & _GEN_111168 : ~(_GEN_111529 & _GEN_1743) & _GEN_111168) : _GEN_111168;
  wire        _GEN_111403 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1744 & _GEN_111169 : _GEN_1143 ? ~_GEN_1744 & _GEN_111169 : ~(_GEN_111529 & _GEN_1744) & _GEN_111169) : _GEN_111169;
  wire        _GEN_111404 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1745 & _GEN_111170 : _GEN_1143 ? ~_GEN_1745 & _GEN_111170 : ~(_GEN_111529 & _GEN_1745) & _GEN_111170) : _GEN_111170;
  wire        _GEN_111405 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1746 & _GEN_111171 : _GEN_1143 ? ~_GEN_1746 & _GEN_111171 : ~(_GEN_111529 & _GEN_1746) & _GEN_111171) : _GEN_111171;
  wire        _GEN_111406 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1747 & _GEN_111172 : _GEN_1143 ? ~_GEN_1747 & _GEN_111172 : ~(_GEN_111529 & _GEN_1747) & _GEN_111172) : _GEN_111172;
  wire        _GEN_111407 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1748 & _GEN_111173 : _GEN_1143 ? ~_GEN_1748 & _GEN_111173 : ~(_GEN_111529 & _GEN_1748) & _GEN_111173) : _GEN_111173;
  wire        _GEN_111408 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1749 & _GEN_111174 : _GEN_1143 ? ~_GEN_1749 & _GEN_111174 : ~(_GEN_111529 & _GEN_1749) & _GEN_111174) : _GEN_111174;
  wire        _GEN_111409 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1750 & _GEN_111175 : _GEN_1143 ? ~_GEN_1750 & _GEN_111175 : ~(_GEN_111529 & _GEN_1750) & _GEN_111175) : _GEN_111175;
  wire        _GEN_111410 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1751 & _GEN_111176 : _GEN_1143 ? ~_GEN_1751 & _GEN_111176 : ~(_GEN_111529 & _GEN_1751) & _GEN_111176) : _GEN_111176;
  wire        _GEN_111411 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1752 & _GEN_111177 : _GEN_1143 ? ~_GEN_1752 & _GEN_111177 : ~(_GEN_111529 & _GEN_1752) & _GEN_111177) : _GEN_111177;
  wire        _GEN_111412 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1753 & _GEN_111178 : _GEN_1143 ? ~_GEN_1753 & _GEN_111178 : ~(_GEN_111529 & _GEN_1753) & _GEN_111178) : _GEN_111178;
  wire        _GEN_111413 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1754 & _GEN_111179 : _GEN_1143 ? ~_GEN_1754 & _GEN_111179 : ~(_GEN_111529 & _GEN_1754) & _GEN_111179) : _GEN_111179;
  wire        _GEN_111414 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1755 & _GEN_111180 : _GEN_1143 ? ~_GEN_1755 & _GEN_111180 : ~(_GEN_111529 & _GEN_1755) & _GEN_111180) : _GEN_111180;
  wire        _GEN_111415 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1756 & _GEN_111181 : _GEN_1143 ? ~_GEN_1756 & _GEN_111181 : ~(_GEN_111529 & _GEN_1756) & _GEN_111181) : _GEN_111181;
  wire        _GEN_111416 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1757 & _GEN_111182 : _GEN_1143 ? ~_GEN_1757 & _GEN_111182 : ~(_GEN_111529 & _GEN_1757) & _GEN_111182) : _GEN_111182;
  wire        _GEN_111417 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1758 & _GEN_111183 : _GEN_1143 ? ~_GEN_1758 & _GEN_111183 : ~(_GEN_111529 & _GEN_1758) & _GEN_111183) : _GEN_111183;
  wire        _GEN_111418 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1759 & _GEN_111184 : _GEN_1143 ? ~_GEN_1759 & _GEN_111184 : ~(_GEN_111529 & _GEN_1759) & _GEN_111184) : _GEN_111184;
  wire        _GEN_111419 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1760 & _GEN_111185 : _GEN_1143 ? ~_GEN_1760 & _GEN_111185 : ~(_GEN_111529 & _GEN_1760) & _GEN_111185) : _GEN_111185;
  wire        _GEN_111420 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1761 & _GEN_111186 : _GEN_1143 ? ~_GEN_1761 & _GEN_111186 : ~(_GEN_111529 & _GEN_1761) & _GEN_111186) : _GEN_111186;
  wire        _GEN_111421 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1762 & _GEN_111187 : _GEN_1143 ? ~_GEN_1762 & _GEN_111187 : ~(_GEN_111529 & _GEN_1762) & _GEN_111187) : _GEN_111187;
  wire        _GEN_111422 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1763 & _GEN_111188 : _GEN_1143 ? ~_GEN_1763 & _GEN_111188 : ~(_GEN_111529 & _GEN_1763) & _GEN_111188) : _GEN_111188;
  wire        _GEN_111423 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1764 & _GEN_111189 : _GEN_1143 ? ~_GEN_1764 & _GEN_111189 : ~(_GEN_111529 & _GEN_1764) & _GEN_111189) : _GEN_111189;
  wire        _GEN_111424 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1765 & _GEN_111190 : _GEN_1143 ? ~_GEN_1765 & _GEN_111190 : ~(_GEN_111529 & _GEN_1765) & _GEN_111190) : _GEN_111190;
  wire        _GEN_111425 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1766 & _GEN_111191 : _GEN_1143 ? ~_GEN_1766 & _GEN_111191 : ~(_GEN_111529 & _GEN_1766) & _GEN_111191) : _GEN_111191;
  wire        _GEN_111426 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1767 & _GEN_111192 : _GEN_1143 ? ~_GEN_1767 & _GEN_111192 : ~(_GEN_111529 & _GEN_1767) & _GEN_111192) : _GEN_111192;
  wire        _GEN_111427 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1768 & _GEN_111193 : _GEN_1143 ? ~_GEN_1768 & _GEN_111193 : ~(_GEN_111529 & _GEN_1768) & _GEN_111193) : _GEN_111193;
  wire        _GEN_111428 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1769 & _GEN_111194 : _GEN_1143 ? ~_GEN_1769 & _GEN_111194 : ~(_GEN_111529 & _GEN_1769) & _GEN_111194) : _GEN_111194;
  wire        _GEN_111429 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1770 & _GEN_111195 : _GEN_1143 ? ~_GEN_1770 & _GEN_111195 : ~(_GEN_111529 & _GEN_1770) & _GEN_111195) : _GEN_111195;
  wire        _GEN_111430 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1771 & _GEN_111196 : _GEN_1143 ? ~_GEN_1771 & _GEN_111196 : ~(_GEN_111529 & _GEN_1771) & _GEN_111196) : _GEN_111196;
  wire        _GEN_111431 = _GEN_1141 ? (_GEN_111364 ? ~_GEN_1772 & _GEN_111197 : _GEN_1143 ? ~_GEN_1772 & _GEN_111197 : ~(_GEN_111529 & _GEN_1772) & _GEN_111197) : _GEN_111197;
  wire        _GEN_111432 = _GEN_1141 ? (_GEN_111364 ? ~(&lcam_ldq_idx_0) & _GEN_111198 : _GEN_1143 ? ~(&lcam_ldq_idx_0) & _GEN_111198 : ~(_GEN_111529 & (&lcam_ldq_idx_0)) & _GEN_111198) : _GEN_111198;
  wire        _GEN_111635 = _GEN_1144 ? (_GEN_111598 ? (|lcam_ldq_idx_1) & _GEN_111401 : _GEN_1146 ? (|lcam_ldq_idx_1) & _GEN_111401 : ~(_GEN_111529 & ~(|lcam_ldq_idx_1)) & _GEN_111401) : _GEN_111401;
  wire        _GEN_111636 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1773 & _GEN_111402 : _GEN_1146 ? ~_GEN_1773 & _GEN_111402 : ~(_GEN_111529 & _GEN_1773) & _GEN_111402) : _GEN_111402;
  wire        _GEN_111637 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1774 & _GEN_111403 : _GEN_1146 ? ~_GEN_1774 & _GEN_111403 : ~(_GEN_111529 & _GEN_1774) & _GEN_111403) : _GEN_111403;
  wire        _GEN_111638 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1775 & _GEN_111404 : _GEN_1146 ? ~_GEN_1775 & _GEN_111404 : ~(_GEN_111529 & _GEN_1775) & _GEN_111404) : _GEN_111404;
  wire        _GEN_111639 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1776 & _GEN_111405 : _GEN_1146 ? ~_GEN_1776 & _GEN_111405 : ~(_GEN_111529 & _GEN_1776) & _GEN_111405) : _GEN_111405;
  wire        _GEN_111640 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1777 & _GEN_111406 : _GEN_1146 ? ~_GEN_1777 & _GEN_111406 : ~(_GEN_111529 & _GEN_1777) & _GEN_111406) : _GEN_111406;
  wire        _GEN_111641 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1778 & _GEN_111407 : _GEN_1146 ? ~_GEN_1778 & _GEN_111407 : ~(_GEN_111529 & _GEN_1778) & _GEN_111407) : _GEN_111407;
  wire        _GEN_111642 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1779 & _GEN_111408 : _GEN_1146 ? ~_GEN_1779 & _GEN_111408 : ~(_GEN_111529 & _GEN_1779) & _GEN_111408) : _GEN_111408;
  wire        _GEN_111643 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1780 & _GEN_111409 : _GEN_1146 ? ~_GEN_1780 & _GEN_111409 : ~(_GEN_111529 & _GEN_1780) & _GEN_111409) : _GEN_111409;
  wire        _GEN_111644 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1781 & _GEN_111410 : _GEN_1146 ? ~_GEN_1781 & _GEN_111410 : ~(_GEN_111529 & _GEN_1781) & _GEN_111410) : _GEN_111410;
  wire        _GEN_111645 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1782 & _GEN_111411 : _GEN_1146 ? ~_GEN_1782 & _GEN_111411 : ~(_GEN_111529 & _GEN_1782) & _GEN_111411) : _GEN_111411;
  wire        _GEN_111646 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1783 & _GEN_111412 : _GEN_1146 ? ~_GEN_1783 & _GEN_111412 : ~(_GEN_111529 & _GEN_1783) & _GEN_111412) : _GEN_111412;
  wire        _GEN_111647 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1784 & _GEN_111413 : _GEN_1146 ? ~_GEN_1784 & _GEN_111413 : ~(_GEN_111529 & _GEN_1784) & _GEN_111413) : _GEN_111413;
  wire        _GEN_111648 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1785 & _GEN_111414 : _GEN_1146 ? ~_GEN_1785 & _GEN_111414 : ~(_GEN_111529 & _GEN_1785) & _GEN_111414) : _GEN_111414;
  wire        _GEN_111649 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1786 & _GEN_111415 : _GEN_1146 ? ~_GEN_1786 & _GEN_111415 : ~(_GEN_111529 & _GEN_1786) & _GEN_111415) : _GEN_111415;
  wire        _GEN_111650 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1787 & _GEN_111416 : _GEN_1146 ? ~_GEN_1787 & _GEN_111416 : ~(_GEN_111529 & _GEN_1787) & _GEN_111416) : _GEN_111416;
  wire        _GEN_111651 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1788 & _GEN_111417 : _GEN_1146 ? ~_GEN_1788 & _GEN_111417 : ~(_GEN_111529 & _GEN_1788) & _GEN_111417) : _GEN_111417;
  wire        _GEN_111652 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1789 & _GEN_111418 : _GEN_1146 ? ~_GEN_1789 & _GEN_111418 : ~(_GEN_111529 & _GEN_1789) & _GEN_111418) : _GEN_111418;
  wire        _GEN_111653 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1790 & _GEN_111419 : _GEN_1146 ? ~_GEN_1790 & _GEN_111419 : ~(_GEN_111529 & _GEN_1790) & _GEN_111419) : _GEN_111419;
  wire        _GEN_111654 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1791 & _GEN_111420 : _GEN_1146 ? ~_GEN_1791 & _GEN_111420 : ~(_GEN_111529 & _GEN_1791) & _GEN_111420) : _GEN_111420;
  wire        _GEN_111655 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1792 & _GEN_111421 : _GEN_1146 ? ~_GEN_1792 & _GEN_111421 : ~(_GEN_111529 & _GEN_1792) & _GEN_111421) : _GEN_111421;
  wire        _GEN_111656 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1793 & _GEN_111422 : _GEN_1146 ? ~_GEN_1793 & _GEN_111422 : ~(_GEN_111529 & _GEN_1793) & _GEN_111422) : _GEN_111422;
  wire        _GEN_111657 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1794 & _GEN_111423 : _GEN_1146 ? ~_GEN_1794 & _GEN_111423 : ~(_GEN_111529 & _GEN_1794) & _GEN_111423) : _GEN_111423;
  wire        _GEN_111658 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1795 & _GEN_111424 : _GEN_1146 ? ~_GEN_1795 & _GEN_111424 : ~(_GEN_111529 & _GEN_1795) & _GEN_111424) : _GEN_111424;
  wire        _GEN_111659 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1796 & _GEN_111425 : _GEN_1146 ? ~_GEN_1796 & _GEN_111425 : ~(_GEN_111529 & _GEN_1796) & _GEN_111425) : _GEN_111425;
  wire        _GEN_111660 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1797 & _GEN_111426 : _GEN_1146 ? ~_GEN_1797 & _GEN_111426 : ~(_GEN_111529 & _GEN_1797) & _GEN_111426) : _GEN_111426;
  wire        _GEN_111661 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1798 & _GEN_111427 : _GEN_1146 ? ~_GEN_1798 & _GEN_111427 : ~(_GEN_111529 & _GEN_1798) & _GEN_111427) : _GEN_111427;
  wire        _GEN_111662 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1799 & _GEN_111428 : _GEN_1146 ? ~_GEN_1799 & _GEN_111428 : ~(_GEN_111529 & _GEN_1799) & _GEN_111428) : _GEN_111428;
  wire        _GEN_111663 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1800 & _GEN_111429 : _GEN_1146 ? ~_GEN_1800 & _GEN_111429 : ~(_GEN_111529 & _GEN_1800) & _GEN_111429) : _GEN_111429;
  wire        _GEN_111664 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1801 & _GEN_111430 : _GEN_1146 ? ~_GEN_1801 & _GEN_111430 : ~(_GEN_111529 & _GEN_1801) & _GEN_111430) : _GEN_111430;
  wire        _GEN_111665 = _GEN_1144 ? (_GEN_111598 ? ~_GEN_1802 & _GEN_111431 : _GEN_1146 ? ~_GEN_1802 & _GEN_111431 : ~(_GEN_111529 & _GEN_1802) & _GEN_111431) : _GEN_111431;
  wire        _GEN_111666 = _GEN_1144 ? (_GEN_111598 ? ~(&lcam_ldq_idx_1) & _GEN_111432 : _GEN_1146 ? ~(&lcam_ldq_idx_1) & _GEN_111432 : ~(_GEN_111529 & (&lcam_ldq_idx_1)) & _GEN_111432) : _GEN_111432;
  wire        _GEN_111869 = _GEN_1147 ? (_GEN_111832 ? (|lcam_ldq_idx_0) & _GEN_111635 : _GEN_1149 ? (|lcam_ldq_idx_0) & _GEN_111635 : ~(_GEN_111997 & ~(|lcam_ldq_idx_0)) & _GEN_111635) : _GEN_111635;
  wire        _GEN_111870 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1743 & _GEN_111636 : _GEN_1149 ? ~_GEN_1743 & _GEN_111636 : ~(_GEN_111997 & _GEN_1743) & _GEN_111636) : _GEN_111636;
  wire        _GEN_111871 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1744 & _GEN_111637 : _GEN_1149 ? ~_GEN_1744 & _GEN_111637 : ~(_GEN_111997 & _GEN_1744) & _GEN_111637) : _GEN_111637;
  wire        _GEN_111872 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1745 & _GEN_111638 : _GEN_1149 ? ~_GEN_1745 & _GEN_111638 : ~(_GEN_111997 & _GEN_1745) & _GEN_111638) : _GEN_111638;
  wire        _GEN_111873 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1746 & _GEN_111639 : _GEN_1149 ? ~_GEN_1746 & _GEN_111639 : ~(_GEN_111997 & _GEN_1746) & _GEN_111639) : _GEN_111639;
  wire        _GEN_111874 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1747 & _GEN_111640 : _GEN_1149 ? ~_GEN_1747 & _GEN_111640 : ~(_GEN_111997 & _GEN_1747) & _GEN_111640) : _GEN_111640;
  wire        _GEN_111875 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1748 & _GEN_111641 : _GEN_1149 ? ~_GEN_1748 & _GEN_111641 : ~(_GEN_111997 & _GEN_1748) & _GEN_111641) : _GEN_111641;
  wire        _GEN_111876 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1749 & _GEN_111642 : _GEN_1149 ? ~_GEN_1749 & _GEN_111642 : ~(_GEN_111997 & _GEN_1749) & _GEN_111642) : _GEN_111642;
  wire        _GEN_111877 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1750 & _GEN_111643 : _GEN_1149 ? ~_GEN_1750 & _GEN_111643 : ~(_GEN_111997 & _GEN_1750) & _GEN_111643) : _GEN_111643;
  wire        _GEN_111878 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1751 & _GEN_111644 : _GEN_1149 ? ~_GEN_1751 & _GEN_111644 : ~(_GEN_111997 & _GEN_1751) & _GEN_111644) : _GEN_111644;
  wire        _GEN_111879 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1752 & _GEN_111645 : _GEN_1149 ? ~_GEN_1752 & _GEN_111645 : ~(_GEN_111997 & _GEN_1752) & _GEN_111645) : _GEN_111645;
  wire        _GEN_111880 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1753 & _GEN_111646 : _GEN_1149 ? ~_GEN_1753 & _GEN_111646 : ~(_GEN_111997 & _GEN_1753) & _GEN_111646) : _GEN_111646;
  wire        _GEN_111881 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1754 & _GEN_111647 : _GEN_1149 ? ~_GEN_1754 & _GEN_111647 : ~(_GEN_111997 & _GEN_1754) & _GEN_111647) : _GEN_111647;
  wire        _GEN_111882 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1755 & _GEN_111648 : _GEN_1149 ? ~_GEN_1755 & _GEN_111648 : ~(_GEN_111997 & _GEN_1755) & _GEN_111648) : _GEN_111648;
  wire        _GEN_111883 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1756 & _GEN_111649 : _GEN_1149 ? ~_GEN_1756 & _GEN_111649 : ~(_GEN_111997 & _GEN_1756) & _GEN_111649) : _GEN_111649;
  wire        _GEN_111884 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1757 & _GEN_111650 : _GEN_1149 ? ~_GEN_1757 & _GEN_111650 : ~(_GEN_111997 & _GEN_1757) & _GEN_111650) : _GEN_111650;
  wire        _GEN_111885 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1758 & _GEN_111651 : _GEN_1149 ? ~_GEN_1758 & _GEN_111651 : ~(_GEN_111997 & _GEN_1758) & _GEN_111651) : _GEN_111651;
  wire        _GEN_111886 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1759 & _GEN_111652 : _GEN_1149 ? ~_GEN_1759 & _GEN_111652 : ~(_GEN_111997 & _GEN_1759) & _GEN_111652) : _GEN_111652;
  wire        _GEN_111887 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1760 & _GEN_111653 : _GEN_1149 ? ~_GEN_1760 & _GEN_111653 : ~(_GEN_111997 & _GEN_1760) & _GEN_111653) : _GEN_111653;
  wire        _GEN_111888 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1761 & _GEN_111654 : _GEN_1149 ? ~_GEN_1761 & _GEN_111654 : ~(_GEN_111997 & _GEN_1761) & _GEN_111654) : _GEN_111654;
  wire        _GEN_111889 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1762 & _GEN_111655 : _GEN_1149 ? ~_GEN_1762 & _GEN_111655 : ~(_GEN_111997 & _GEN_1762) & _GEN_111655) : _GEN_111655;
  wire        _GEN_111890 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1763 & _GEN_111656 : _GEN_1149 ? ~_GEN_1763 & _GEN_111656 : ~(_GEN_111997 & _GEN_1763) & _GEN_111656) : _GEN_111656;
  wire        _GEN_111891 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1764 & _GEN_111657 : _GEN_1149 ? ~_GEN_1764 & _GEN_111657 : ~(_GEN_111997 & _GEN_1764) & _GEN_111657) : _GEN_111657;
  wire        _GEN_111892 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1765 & _GEN_111658 : _GEN_1149 ? ~_GEN_1765 & _GEN_111658 : ~(_GEN_111997 & _GEN_1765) & _GEN_111658) : _GEN_111658;
  wire        _GEN_111893 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1766 & _GEN_111659 : _GEN_1149 ? ~_GEN_1766 & _GEN_111659 : ~(_GEN_111997 & _GEN_1766) & _GEN_111659) : _GEN_111659;
  wire        _GEN_111894 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1767 & _GEN_111660 : _GEN_1149 ? ~_GEN_1767 & _GEN_111660 : ~(_GEN_111997 & _GEN_1767) & _GEN_111660) : _GEN_111660;
  wire        _GEN_111895 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1768 & _GEN_111661 : _GEN_1149 ? ~_GEN_1768 & _GEN_111661 : ~(_GEN_111997 & _GEN_1768) & _GEN_111661) : _GEN_111661;
  wire        _GEN_111896 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1769 & _GEN_111662 : _GEN_1149 ? ~_GEN_1769 & _GEN_111662 : ~(_GEN_111997 & _GEN_1769) & _GEN_111662) : _GEN_111662;
  wire        _GEN_111897 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1770 & _GEN_111663 : _GEN_1149 ? ~_GEN_1770 & _GEN_111663 : ~(_GEN_111997 & _GEN_1770) & _GEN_111663) : _GEN_111663;
  wire        _GEN_111898 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1771 & _GEN_111664 : _GEN_1149 ? ~_GEN_1771 & _GEN_111664 : ~(_GEN_111997 & _GEN_1771) & _GEN_111664) : _GEN_111664;
  wire        _GEN_111899 = _GEN_1147 ? (_GEN_111832 ? ~_GEN_1772 & _GEN_111665 : _GEN_1149 ? ~_GEN_1772 & _GEN_111665 : ~(_GEN_111997 & _GEN_1772) & _GEN_111665) : _GEN_111665;
  wire        _GEN_111900 = _GEN_1147 ? (_GEN_111832 ? ~(&lcam_ldq_idx_0) & _GEN_111666 : _GEN_1149 ? ~(&lcam_ldq_idx_0) & _GEN_111666 : ~(_GEN_111997 & (&lcam_ldq_idx_0)) & _GEN_111666) : _GEN_111666;
  wire        _GEN_112103 = _GEN_1150 ? (_GEN_112066 ? (|lcam_ldq_idx_1) & _GEN_111869 : _GEN_1152 ? (|lcam_ldq_idx_1) & _GEN_111869 : ~(_GEN_111997 & ~(|lcam_ldq_idx_1)) & _GEN_111869) : _GEN_111869;
  wire        _GEN_112104 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1773 & _GEN_111870 : _GEN_1152 ? ~_GEN_1773 & _GEN_111870 : ~(_GEN_111997 & _GEN_1773) & _GEN_111870) : _GEN_111870;
  wire        _GEN_112105 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1774 & _GEN_111871 : _GEN_1152 ? ~_GEN_1774 & _GEN_111871 : ~(_GEN_111997 & _GEN_1774) & _GEN_111871) : _GEN_111871;
  wire        _GEN_112106 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1775 & _GEN_111872 : _GEN_1152 ? ~_GEN_1775 & _GEN_111872 : ~(_GEN_111997 & _GEN_1775) & _GEN_111872) : _GEN_111872;
  wire        _GEN_112107 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1776 & _GEN_111873 : _GEN_1152 ? ~_GEN_1776 & _GEN_111873 : ~(_GEN_111997 & _GEN_1776) & _GEN_111873) : _GEN_111873;
  wire        _GEN_112108 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1777 & _GEN_111874 : _GEN_1152 ? ~_GEN_1777 & _GEN_111874 : ~(_GEN_111997 & _GEN_1777) & _GEN_111874) : _GEN_111874;
  wire        _GEN_112109 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1778 & _GEN_111875 : _GEN_1152 ? ~_GEN_1778 & _GEN_111875 : ~(_GEN_111997 & _GEN_1778) & _GEN_111875) : _GEN_111875;
  wire        _GEN_112110 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1779 & _GEN_111876 : _GEN_1152 ? ~_GEN_1779 & _GEN_111876 : ~(_GEN_111997 & _GEN_1779) & _GEN_111876) : _GEN_111876;
  wire        _GEN_112111 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1780 & _GEN_111877 : _GEN_1152 ? ~_GEN_1780 & _GEN_111877 : ~(_GEN_111997 & _GEN_1780) & _GEN_111877) : _GEN_111877;
  wire        _GEN_112112 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1781 & _GEN_111878 : _GEN_1152 ? ~_GEN_1781 & _GEN_111878 : ~(_GEN_111997 & _GEN_1781) & _GEN_111878) : _GEN_111878;
  wire        _GEN_112113 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1782 & _GEN_111879 : _GEN_1152 ? ~_GEN_1782 & _GEN_111879 : ~(_GEN_111997 & _GEN_1782) & _GEN_111879) : _GEN_111879;
  wire        _GEN_112114 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1783 & _GEN_111880 : _GEN_1152 ? ~_GEN_1783 & _GEN_111880 : ~(_GEN_111997 & _GEN_1783) & _GEN_111880) : _GEN_111880;
  wire        _GEN_112115 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1784 & _GEN_111881 : _GEN_1152 ? ~_GEN_1784 & _GEN_111881 : ~(_GEN_111997 & _GEN_1784) & _GEN_111881) : _GEN_111881;
  wire        _GEN_112116 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1785 & _GEN_111882 : _GEN_1152 ? ~_GEN_1785 & _GEN_111882 : ~(_GEN_111997 & _GEN_1785) & _GEN_111882) : _GEN_111882;
  wire        _GEN_112117 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1786 & _GEN_111883 : _GEN_1152 ? ~_GEN_1786 & _GEN_111883 : ~(_GEN_111997 & _GEN_1786) & _GEN_111883) : _GEN_111883;
  wire        _GEN_112118 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1787 & _GEN_111884 : _GEN_1152 ? ~_GEN_1787 & _GEN_111884 : ~(_GEN_111997 & _GEN_1787) & _GEN_111884) : _GEN_111884;
  wire        _GEN_112119 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1788 & _GEN_111885 : _GEN_1152 ? ~_GEN_1788 & _GEN_111885 : ~(_GEN_111997 & _GEN_1788) & _GEN_111885) : _GEN_111885;
  wire        _GEN_112120 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1789 & _GEN_111886 : _GEN_1152 ? ~_GEN_1789 & _GEN_111886 : ~(_GEN_111997 & _GEN_1789) & _GEN_111886) : _GEN_111886;
  wire        _GEN_112121 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1790 & _GEN_111887 : _GEN_1152 ? ~_GEN_1790 & _GEN_111887 : ~(_GEN_111997 & _GEN_1790) & _GEN_111887) : _GEN_111887;
  wire        _GEN_112122 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1791 & _GEN_111888 : _GEN_1152 ? ~_GEN_1791 & _GEN_111888 : ~(_GEN_111997 & _GEN_1791) & _GEN_111888) : _GEN_111888;
  wire        _GEN_112123 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1792 & _GEN_111889 : _GEN_1152 ? ~_GEN_1792 & _GEN_111889 : ~(_GEN_111997 & _GEN_1792) & _GEN_111889) : _GEN_111889;
  wire        _GEN_112124 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1793 & _GEN_111890 : _GEN_1152 ? ~_GEN_1793 & _GEN_111890 : ~(_GEN_111997 & _GEN_1793) & _GEN_111890) : _GEN_111890;
  wire        _GEN_112125 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1794 & _GEN_111891 : _GEN_1152 ? ~_GEN_1794 & _GEN_111891 : ~(_GEN_111997 & _GEN_1794) & _GEN_111891) : _GEN_111891;
  wire        _GEN_112126 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1795 & _GEN_111892 : _GEN_1152 ? ~_GEN_1795 & _GEN_111892 : ~(_GEN_111997 & _GEN_1795) & _GEN_111892) : _GEN_111892;
  wire        _GEN_112127 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1796 & _GEN_111893 : _GEN_1152 ? ~_GEN_1796 & _GEN_111893 : ~(_GEN_111997 & _GEN_1796) & _GEN_111893) : _GEN_111893;
  wire        _GEN_112128 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1797 & _GEN_111894 : _GEN_1152 ? ~_GEN_1797 & _GEN_111894 : ~(_GEN_111997 & _GEN_1797) & _GEN_111894) : _GEN_111894;
  wire        _GEN_112129 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1798 & _GEN_111895 : _GEN_1152 ? ~_GEN_1798 & _GEN_111895 : ~(_GEN_111997 & _GEN_1798) & _GEN_111895) : _GEN_111895;
  wire        _GEN_112130 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1799 & _GEN_111896 : _GEN_1152 ? ~_GEN_1799 & _GEN_111896 : ~(_GEN_111997 & _GEN_1799) & _GEN_111896) : _GEN_111896;
  wire        _GEN_112131 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1800 & _GEN_111897 : _GEN_1152 ? ~_GEN_1800 & _GEN_111897 : ~(_GEN_111997 & _GEN_1800) & _GEN_111897) : _GEN_111897;
  wire        _GEN_112132 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1801 & _GEN_111898 : _GEN_1152 ? ~_GEN_1801 & _GEN_111898 : ~(_GEN_111997 & _GEN_1801) & _GEN_111898) : _GEN_111898;
  wire        _GEN_112133 = _GEN_1150 ? (_GEN_112066 ? ~_GEN_1802 & _GEN_111899 : _GEN_1152 ? ~_GEN_1802 & _GEN_111899 : ~(_GEN_111997 & _GEN_1802) & _GEN_111899) : _GEN_111899;
  wire        _GEN_112134 = _GEN_1150 ? (_GEN_112066 ? ~(&lcam_ldq_idx_1) & _GEN_111900 : _GEN_1152 ? ~(&lcam_ldq_idx_1) & _GEN_111900 : ~(_GEN_111997 & (&lcam_ldq_idx_1)) & _GEN_111900) : _GEN_111900;
  wire        _GEN_112337 = _GEN_1153 ? (_GEN_112300 ? (|lcam_ldq_idx_0) & _GEN_112103 : _GEN_1155 ? (|lcam_ldq_idx_0) & _GEN_112103 : ~(_GEN_112465 & ~(|lcam_ldq_idx_0)) & _GEN_112103) : _GEN_112103;
  wire        _GEN_112338 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1743 & _GEN_112104 : _GEN_1155 ? ~_GEN_1743 & _GEN_112104 : ~(_GEN_112465 & _GEN_1743) & _GEN_112104) : _GEN_112104;
  wire        _GEN_112339 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1744 & _GEN_112105 : _GEN_1155 ? ~_GEN_1744 & _GEN_112105 : ~(_GEN_112465 & _GEN_1744) & _GEN_112105) : _GEN_112105;
  wire        _GEN_112340 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1745 & _GEN_112106 : _GEN_1155 ? ~_GEN_1745 & _GEN_112106 : ~(_GEN_112465 & _GEN_1745) & _GEN_112106) : _GEN_112106;
  wire        _GEN_112341 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1746 & _GEN_112107 : _GEN_1155 ? ~_GEN_1746 & _GEN_112107 : ~(_GEN_112465 & _GEN_1746) & _GEN_112107) : _GEN_112107;
  wire        _GEN_112342 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1747 & _GEN_112108 : _GEN_1155 ? ~_GEN_1747 & _GEN_112108 : ~(_GEN_112465 & _GEN_1747) & _GEN_112108) : _GEN_112108;
  wire        _GEN_112343 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1748 & _GEN_112109 : _GEN_1155 ? ~_GEN_1748 & _GEN_112109 : ~(_GEN_112465 & _GEN_1748) & _GEN_112109) : _GEN_112109;
  wire        _GEN_112344 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1749 & _GEN_112110 : _GEN_1155 ? ~_GEN_1749 & _GEN_112110 : ~(_GEN_112465 & _GEN_1749) & _GEN_112110) : _GEN_112110;
  wire        _GEN_112345 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1750 & _GEN_112111 : _GEN_1155 ? ~_GEN_1750 & _GEN_112111 : ~(_GEN_112465 & _GEN_1750) & _GEN_112111) : _GEN_112111;
  wire        _GEN_112346 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1751 & _GEN_112112 : _GEN_1155 ? ~_GEN_1751 & _GEN_112112 : ~(_GEN_112465 & _GEN_1751) & _GEN_112112) : _GEN_112112;
  wire        _GEN_112347 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1752 & _GEN_112113 : _GEN_1155 ? ~_GEN_1752 & _GEN_112113 : ~(_GEN_112465 & _GEN_1752) & _GEN_112113) : _GEN_112113;
  wire        _GEN_112348 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1753 & _GEN_112114 : _GEN_1155 ? ~_GEN_1753 & _GEN_112114 : ~(_GEN_112465 & _GEN_1753) & _GEN_112114) : _GEN_112114;
  wire        _GEN_112349 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1754 & _GEN_112115 : _GEN_1155 ? ~_GEN_1754 & _GEN_112115 : ~(_GEN_112465 & _GEN_1754) & _GEN_112115) : _GEN_112115;
  wire        _GEN_112350 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1755 & _GEN_112116 : _GEN_1155 ? ~_GEN_1755 & _GEN_112116 : ~(_GEN_112465 & _GEN_1755) & _GEN_112116) : _GEN_112116;
  wire        _GEN_112351 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1756 & _GEN_112117 : _GEN_1155 ? ~_GEN_1756 & _GEN_112117 : ~(_GEN_112465 & _GEN_1756) & _GEN_112117) : _GEN_112117;
  wire        _GEN_112352 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1757 & _GEN_112118 : _GEN_1155 ? ~_GEN_1757 & _GEN_112118 : ~(_GEN_112465 & _GEN_1757) & _GEN_112118) : _GEN_112118;
  wire        _GEN_112353 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1758 & _GEN_112119 : _GEN_1155 ? ~_GEN_1758 & _GEN_112119 : ~(_GEN_112465 & _GEN_1758) & _GEN_112119) : _GEN_112119;
  wire        _GEN_112354 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1759 & _GEN_112120 : _GEN_1155 ? ~_GEN_1759 & _GEN_112120 : ~(_GEN_112465 & _GEN_1759) & _GEN_112120) : _GEN_112120;
  wire        _GEN_112355 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1760 & _GEN_112121 : _GEN_1155 ? ~_GEN_1760 & _GEN_112121 : ~(_GEN_112465 & _GEN_1760) & _GEN_112121) : _GEN_112121;
  wire        _GEN_112356 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1761 & _GEN_112122 : _GEN_1155 ? ~_GEN_1761 & _GEN_112122 : ~(_GEN_112465 & _GEN_1761) & _GEN_112122) : _GEN_112122;
  wire        _GEN_112357 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1762 & _GEN_112123 : _GEN_1155 ? ~_GEN_1762 & _GEN_112123 : ~(_GEN_112465 & _GEN_1762) & _GEN_112123) : _GEN_112123;
  wire        _GEN_112358 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1763 & _GEN_112124 : _GEN_1155 ? ~_GEN_1763 & _GEN_112124 : ~(_GEN_112465 & _GEN_1763) & _GEN_112124) : _GEN_112124;
  wire        _GEN_112359 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1764 & _GEN_112125 : _GEN_1155 ? ~_GEN_1764 & _GEN_112125 : ~(_GEN_112465 & _GEN_1764) & _GEN_112125) : _GEN_112125;
  wire        _GEN_112360 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1765 & _GEN_112126 : _GEN_1155 ? ~_GEN_1765 & _GEN_112126 : ~(_GEN_112465 & _GEN_1765) & _GEN_112126) : _GEN_112126;
  wire        _GEN_112361 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1766 & _GEN_112127 : _GEN_1155 ? ~_GEN_1766 & _GEN_112127 : ~(_GEN_112465 & _GEN_1766) & _GEN_112127) : _GEN_112127;
  wire        _GEN_112362 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1767 & _GEN_112128 : _GEN_1155 ? ~_GEN_1767 & _GEN_112128 : ~(_GEN_112465 & _GEN_1767) & _GEN_112128) : _GEN_112128;
  wire        _GEN_112363 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1768 & _GEN_112129 : _GEN_1155 ? ~_GEN_1768 & _GEN_112129 : ~(_GEN_112465 & _GEN_1768) & _GEN_112129) : _GEN_112129;
  wire        _GEN_112364 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1769 & _GEN_112130 : _GEN_1155 ? ~_GEN_1769 & _GEN_112130 : ~(_GEN_112465 & _GEN_1769) & _GEN_112130) : _GEN_112130;
  wire        _GEN_112365 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1770 & _GEN_112131 : _GEN_1155 ? ~_GEN_1770 & _GEN_112131 : ~(_GEN_112465 & _GEN_1770) & _GEN_112131) : _GEN_112131;
  wire        _GEN_112366 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1771 & _GEN_112132 : _GEN_1155 ? ~_GEN_1771 & _GEN_112132 : ~(_GEN_112465 & _GEN_1771) & _GEN_112132) : _GEN_112132;
  wire        _GEN_112367 = _GEN_1153 ? (_GEN_112300 ? ~_GEN_1772 & _GEN_112133 : _GEN_1155 ? ~_GEN_1772 & _GEN_112133 : ~(_GEN_112465 & _GEN_1772) & _GEN_112133) : _GEN_112133;
  wire        _GEN_112368 = _GEN_1153 ? (_GEN_112300 ? ~(&lcam_ldq_idx_0) & _GEN_112134 : _GEN_1155 ? ~(&lcam_ldq_idx_0) & _GEN_112134 : ~(_GEN_112465 & (&lcam_ldq_idx_0)) & _GEN_112134) : _GEN_112134;
  wire        _GEN_112571 = _GEN_1156 ? (_GEN_112534 ? (|lcam_ldq_idx_1) & _GEN_112337 : _GEN_1158 ? (|lcam_ldq_idx_1) & _GEN_112337 : ~(_GEN_112465 & ~(|lcam_ldq_idx_1)) & _GEN_112337) : _GEN_112337;
  wire        _GEN_112572 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1773 & _GEN_112338 : _GEN_1158 ? ~_GEN_1773 & _GEN_112338 : ~(_GEN_112465 & _GEN_1773) & _GEN_112338) : _GEN_112338;
  wire        _GEN_112573 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1774 & _GEN_112339 : _GEN_1158 ? ~_GEN_1774 & _GEN_112339 : ~(_GEN_112465 & _GEN_1774) & _GEN_112339) : _GEN_112339;
  wire        _GEN_112574 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1775 & _GEN_112340 : _GEN_1158 ? ~_GEN_1775 & _GEN_112340 : ~(_GEN_112465 & _GEN_1775) & _GEN_112340) : _GEN_112340;
  wire        _GEN_112575 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1776 & _GEN_112341 : _GEN_1158 ? ~_GEN_1776 & _GEN_112341 : ~(_GEN_112465 & _GEN_1776) & _GEN_112341) : _GEN_112341;
  wire        _GEN_112576 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1777 & _GEN_112342 : _GEN_1158 ? ~_GEN_1777 & _GEN_112342 : ~(_GEN_112465 & _GEN_1777) & _GEN_112342) : _GEN_112342;
  wire        _GEN_112577 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1778 & _GEN_112343 : _GEN_1158 ? ~_GEN_1778 & _GEN_112343 : ~(_GEN_112465 & _GEN_1778) & _GEN_112343) : _GEN_112343;
  wire        _GEN_112578 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1779 & _GEN_112344 : _GEN_1158 ? ~_GEN_1779 & _GEN_112344 : ~(_GEN_112465 & _GEN_1779) & _GEN_112344) : _GEN_112344;
  wire        _GEN_112579 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1780 & _GEN_112345 : _GEN_1158 ? ~_GEN_1780 & _GEN_112345 : ~(_GEN_112465 & _GEN_1780) & _GEN_112345) : _GEN_112345;
  wire        _GEN_112580 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1781 & _GEN_112346 : _GEN_1158 ? ~_GEN_1781 & _GEN_112346 : ~(_GEN_112465 & _GEN_1781) & _GEN_112346) : _GEN_112346;
  wire        _GEN_112581 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1782 & _GEN_112347 : _GEN_1158 ? ~_GEN_1782 & _GEN_112347 : ~(_GEN_112465 & _GEN_1782) & _GEN_112347) : _GEN_112347;
  wire        _GEN_112582 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1783 & _GEN_112348 : _GEN_1158 ? ~_GEN_1783 & _GEN_112348 : ~(_GEN_112465 & _GEN_1783) & _GEN_112348) : _GEN_112348;
  wire        _GEN_112583 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1784 & _GEN_112349 : _GEN_1158 ? ~_GEN_1784 & _GEN_112349 : ~(_GEN_112465 & _GEN_1784) & _GEN_112349) : _GEN_112349;
  wire        _GEN_112584 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1785 & _GEN_112350 : _GEN_1158 ? ~_GEN_1785 & _GEN_112350 : ~(_GEN_112465 & _GEN_1785) & _GEN_112350) : _GEN_112350;
  wire        _GEN_112585 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1786 & _GEN_112351 : _GEN_1158 ? ~_GEN_1786 & _GEN_112351 : ~(_GEN_112465 & _GEN_1786) & _GEN_112351) : _GEN_112351;
  wire        _GEN_112586 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1787 & _GEN_112352 : _GEN_1158 ? ~_GEN_1787 & _GEN_112352 : ~(_GEN_112465 & _GEN_1787) & _GEN_112352) : _GEN_112352;
  wire        _GEN_112587 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1788 & _GEN_112353 : _GEN_1158 ? ~_GEN_1788 & _GEN_112353 : ~(_GEN_112465 & _GEN_1788) & _GEN_112353) : _GEN_112353;
  wire        _GEN_112588 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1789 & _GEN_112354 : _GEN_1158 ? ~_GEN_1789 & _GEN_112354 : ~(_GEN_112465 & _GEN_1789) & _GEN_112354) : _GEN_112354;
  wire        _GEN_112589 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1790 & _GEN_112355 : _GEN_1158 ? ~_GEN_1790 & _GEN_112355 : ~(_GEN_112465 & _GEN_1790) & _GEN_112355) : _GEN_112355;
  wire        _GEN_112590 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1791 & _GEN_112356 : _GEN_1158 ? ~_GEN_1791 & _GEN_112356 : ~(_GEN_112465 & _GEN_1791) & _GEN_112356) : _GEN_112356;
  wire        _GEN_112591 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1792 & _GEN_112357 : _GEN_1158 ? ~_GEN_1792 & _GEN_112357 : ~(_GEN_112465 & _GEN_1792) & _GEN_112357) : _GEN_112357;
  wire        _GEN_112592 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1793 & _GEN_112358 : _GEN_1158 ? ~_GEN_1793 & _GEN_112358 : ~(_GEN_112465 & _GEN_1793) & _GEN_112358) : _GEN_112358;
  wire        _GEN_112593 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1794 & _GEN_112359 : _GEN_1158 ? ~_GEN_1794 & _GEN_112359 : ~(_GEN_112465 & _GEN_1794) & _GEN_112359) : _GEN_112359;
  wire        _GEN_112594 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1795 & _GEN_112360 : _GEN_1158 ? ~_GEN_1795 & _GEN_112360 : ~(_GEN_112465 & _GEN_1795) & _GEN_112360) : _GEN_112360;
  wire        _GEN_112595 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1796 & _GEN_112361 : _GEN_1158 ? ~_GEN_1796 & _GEN_112361 : ~(_GEN_112465 & _GEN_1796) & _GEN_112361) : _GEN_112361;
  wire        _GEN_112596 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1797 & _GEN_112362 : _GEN_1158 ? ~_GEN_1797 & _GEN_112362 : ~(_GEN_112465 & _GEN_1797) & _GEN_112362) : _GEN_112362;
  wire        _GEN_112597 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1798 & _GEN_112363 : _GEN_1158 ? ~_GEN_1798 & _GEN_112363 : ~(_GEN_112465 & _GEN_1798) & _GEN_112363) : _GEN_112363;
  wire        _GEN_112598 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1799 & _GEN_112364 : _GEN_1158 ? ~_GEN_1799 & _GEN_112364 : ~(_GEN_112465 & _GEN_1799) & _GEN_112364) : _GEN_112364;
  wire        _GEN_112599 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1800 & _GEN_112365 : _GEN_1158 ? ~_GEN_1800 & _GEN_112365 : ~(_GEN_112465 & _GEN_1800) & _GEN_112365) : _GEN_112365;
  wire        _GEN_112600 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1801 & _GEN_112366 : _GEN_1158 ? ~_GEN_1801 & _GEN_112366 : ~(_GEN_112465 & _GEN_1801) & _GEN_112366) : _GEN_112366;
  wire        _GEN_112601 = _GEN_1156 ? (_GEN_112534 ? ~_GEN_1802 & _GEN_112367 : _GEN_1158 ? ~_GEN_1802 & _GEN_112367 : ~(_GEN_112465 & _GEN_1802) & _GEN_112367) : _GEN_112367;
  wire        _GEN_112602 = _GEN_1156 ? (_GEN_112534 ? ~(&lcam_ldq_idx_1) & _GEN_112368 : _GEN_1158 ? ~(&lcam_ldq_idx_1) & _GEN_112368 : ~(_GEN_112465 & (&lcam_ldq_idx_1)) & _GEN_112368) : _GEN_112368;
  wire        _GEN_112805 = _GEN_1159 ? (_GEN_112768 ? (|lcam_ldq_idx_0) & _GEN_112571 : _GEN_1161 ? (|lcam_ldq_idx_0) & _GEN_112571 : ~(_GEN_112933 & ~(|lcam_ldq_idx_0)) & _GEN_112571) : _GEN_112571;
  wire        _GEN_112806 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1743 & _GEN_112572 : _GEN_1161 ? ~_GEN_1743 & _GEN_112572 : ~(_GEN_112933 & _GEN_1743) & _GEN_112572) : _GEN_112572;
  wire        _GEN_112807 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1744 & _GEN_112573 : _GEN_1161 ? ~_GEN_1744 & _GEN_112573 : ~(_GEN_112933 & _GEN_1744) & _GEN_112573) : _GEN_112573;
  wire        _GEN_112808 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1745 & _GEN_112574 : _GEN_1161 ? ~_GEN_1745 & _GEN_112574 : ~(_GEN_112933 & _GEN_1745) & _GEN_112574) : _GEN_112574;
  wire        _GEN_112809 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1746 & _GEN_112575 : _GEN_1161 ? ~_GEN_1746 & _GEN_112575 : ~(_GEN_112933 & _GEN_1746) & _GEN_112575) : _GEN_112575;
  wire        _GEN_112810 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1747 & _GEN_112576 : _GEN_1161 ? ~_GEN_1747 & _GEN_112576 : ~(_GEN_112933 & _GEN_1747) & _GEN_112576) : _GEN_112576;
  wire        _GEN_112811 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1748 & _GEN_112577 : _GEN_1161 ? ~_GEN_1748 & _GEN_112577 : ~(_GEN_112933 & _GEN_1748) & _GEN_112577) : _GEN_112577;
  wire        _GEN_112812 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1749 & _GEN_112578 : _GEN_1161 ? ~_GEN_1749 & _GEN_112578 : ~(_GEN_112933 & _GEN_1749) & _GEN_112578) : _GEN_112578;
  wire        _GEN_112813 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1750 & _GEN_112579 : _GEN_1161 ? ~_GEN_1750 & _GEN_112579 : ~(_GEN_112933 & _GEN_1750) & _GEN_112579) : _GEN_112579;
  wire        _GEN_112814 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1751 & _GEN_112580 : _GEN_1161 ? ~_GEN_1751 & _GEN_112580 : ~(_GEN_112933 & _GEN_1751) & _GEN_112580) : _GEN_112580;
  wire        _GEN_112815 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1752 & _GEN_112581 : _GEN_1161 ? ~_GEN_1752 & _GEN_112581 : ~(_GEN_112933 & _GEN_1752) & _GEN_112581) : _GEN_112581;
  wire        _GEN_112816 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1753 & _GEN_112582 : _GEN_1161 ? ~_GEN_1753 & _GEN_112582 : ~(_GEN_112933 & _GEN_1753) & _GEN_112582) : _GEN_112582;
  wire        _GEN_112817 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1754 & _GEN_112583 : _GEN_1161 ? ~_GEN_1754 & _GEN_112583 : ~(_GEN_112933 & _GEN_1754) & _GEN_112583) : _GEN_112583;
  wire        _GEN_112818 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1755 & _GEN_112584 : _GEN_1161 ? ~_GEN_1755 & _GEN_112584 : ~(_GEN_112933 & _GEN_1755) & _GEN_112584) : _GEN_112584;
  wire        _GEN_112819 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1756 & _GEN_112585 : _GEN_1161 ? ~_GEN_1756 & _GEN_112585 : ~(_GEN_112933 & _GEN_1756) & _GEN_112585) : _GEN_112585;
  wire        _GEN_112820 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1757 & _GEN_112586 : _GEN_1161 ? ~_GEN_1757 & _GEN_112586 : ~(_GEN_112933 & _GEN_1757) & _GEN_112586) : _GEN_112586;
  wire        _GEN_112821 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1758 & _GEN_112587 : _GEN_1161 ? ~_GEN_1758 & _GEN_112587 : ~(_GEN_112933 & _GEN_1758) & _GEN_112587) : _GEN_112587;
  wire        _GEN_112822 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1759 & _GEN_112588 : _GEN_1161 ? ~_GEN_1759 & _GEN_112588 : ~(_GEN_112933 & _GEN_1759) & _GEN_112588) : _GEN_112588;
  wire        _GEN_112823 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1760 & _GEN_112589 : _GEN_1161 ? ~_GEN_1760 & _GEN_112589 : ~(_GEN_112933 & _GEN_1760) & _GEN_112589) : _GEN_112589;
  wire        _GEN_112824 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1761 & _GEN_112590 : _GEN_1161 ? ~_GEN_1761 & _GEN_112590 : ~(_GEN_112933 & _GEN_1761) & _GEN_112590) : _GEN_112590;
  wire        _GEN_112825 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1762 & _GEN_112591 : _GEN_1161 ? ~_GEN_1762 & _GEN_112591 : ~(_GEN_112933 & _GEN_1762) & _GEN_112591) : _GEN_112591;
  wire        _GEN_112826 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1763 & _GEN_112592 : _GEN_1161 ? ~_GEN_1763 & _GEN_112592 : ~(_GEN_112933 & _GEN_1763) & _GEN_112592) : _GEN_112592;
  wire        _GEN_112827 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1764 & _GEN_112593 : _GEN_1161 ? ~_GEN_1764 & _GEN_112593 : ~(_GEN_112933 & _GEN_1764) & _GEN_112593) : _GEN_112593;
  wire        _GEN_112828 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1765 & _GEN_112594 : _GEN_1161 ? ~_GEN_1765 & _GEN_112594 : ~(_GEN_112933 & _GEN_1765) & _GEN_112594) : _GEN_112594;
  wire        _GEN_112829 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1766 & _GEN_112595 : _GEN_1161 ? ~_GEN_1766 & _GEN_112595 : ~(_GEN_112933 & _GEN_1766) & _GEN_112595) : _GEN_112595;
  wire        _GEN_112830 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1767 & _GEN_112596 : _GEN_1161 ? ~_GEN_1767 & _GEN_112596 : ~(_GEN_112933 & _GEN_1767) & _GEN_112596) : _GEN_112596;
  wire        _GEN_112831 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1768 & _GEN_112597 : _GEN_1161 ? ~_GEN_1768 & _GEN_112597 : ~(_GEN_112933 & _GEN_1768) & _GEN_112597) : _GEN_112597;
  wire        _GEN_112832 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1769 & _GEN_112598 : _GEN_1161 ? ~_GEN_1769 & _GEN_112598 : ~(_GEN_112933 & _GEN_1769) & _GEN_112598) : _GEN_112598;
  wire        _GEN_112833 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1770 & _GEN_112599 : _GEN_1161 ? ~_GEN_1770 & _GEN_112599 : ~(_GEN_112933 & _GEN_1770) & _GEN_112599) : _GEN_112599;
  wire        _GEN_112834 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1771 & _GEN_112600 : _GEN_1161 ? ~_GEN_1771 & _GEN_112600 : ~(_GEN_112933 & _GEN_1771) & _GEN_112600) : _GEN_112600;
  wire        _GEN_112835 = _GEN_1159 ? (_GEN_112768 ? ~_GEN_1772 & _GEN_112601 : _GEN_1161 ? ~_GEN_1772 & _GEN_112601 : ~(_GEN_112933 & _GEN_1772) & _GEN_112601) : _GEN_112601;
  wire        _GEN_112836 = _GEN_1159 ? (_GEN_112768 ? ~(&lcam_ldq_idx_0) & _GEN_112602 : _GEN_1161 ? ~(&lcam_ldq_idx_0) & _GEN_112602 : ~(_GEN_112933 & (&lcam_ldq_idx_0)) & _GEN_112602) : _GEN_112602;
  wire        _GEN_113039 = _GEN_1162 ? (_GEN_113002 ? (|lcam_ldq_idx_1) & _GEN_112805 : _GEN_1164 ? (|lcam_ldq_idx_1) & _GEN_112805 : ~(_GEN_112933 & ~(|lcam_ldq_idx_1)) & _GEN_112805) : _GEN_112805;
  wire        _GEN_113040 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1773 & _GEN_112806 : _GEN_1164 ? ~_GEN_1773 & _GEN_112806 : ~(_GEN_112933 & _GEN_1773) & _GEN_112806) : _GEN_112806;
  wire        _GEN_113041 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1774 & _GEN_112807 : _GEN_1164 ? ~_GEN_1774 & _GEN_112807 : ~(_GEN_112933 & _GEN_1774) & _GEN_112807) : _GEN_112807;
  wire        _GEN_113042 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1775 & _GEN_112808 : _GEN_1164 ? ~_GEN_1775 & _GEN_112808 : ~(_GEN_112933 & _GEN_1775) & _GEN_112808) : _GEN_112808;
  wire        _GEN_113043 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1776 & _GEN_112809 : _GEN_1164 ? ~_GEN_1776 & _GEN_112809 : ~(_GEN_112933 & _GEN_1776) & _GEN_112809) : _GEN_112809;
  wire        _GEN_113044 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1777 & _GEN_112810 : _GEN_1164 ? ~_GEN_1777 & _GEN_112810 : ~(_GEN_112933 & _GEN_1777) & _GEN_112810) : _GEN_112810;
  wire        _GEN_113045 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1778 & _GEN_112811 : _GEN_1164 ? ~_GEN_1778 & _GEN_112811 : ~(_GEN_112933 & _GEN_1778) & _GEN_112811) : _GEN_112811;
  wire        _GEN_113046 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1779 & _GEN_112812 : _GEN_1164 ? ~_GEN_1779 & _GEN_112812 : ~(_GEN_112933 & _GEN_1779) & _GEN_112812) : _GEN_112812;
  wire        _GEN_113047 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1780 & _GEN_112813 : _GEN_1164 ? ~_GEN_1780 & _GEN_112813 : ~(_GEN_112933 & _GEN_1780) & _GEN_112813) : _GEN_112813;
  wire        _GEN_113048 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1781 & _GEN_112814 : _GEN_1164 ? ~_GEN_1781 & _GEN_112814 : ~(_GEN_112933 & _GEN_1781) & _GEN_112814) : _GEN_112814;
  wire        _GEN_113049 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1782 & _GEN_112815 : _GEN_1164 ? ~_GEN_1782 & _GEN_112815 : ~(_GEN_112933 & _GEN_1782) & _GEN_112815) : _GEN_112815;
  wire        _GEN_113050 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1783 & _GEN_112816 : _GEN_1164 ? ~_GEN_1783 & _GEN_112816 : ~(_GEN_112933 & _GEN_1783) & _GEN_112816) : _GEN_112816;
  wire        _GEN_113051 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1784 & _GEN_112817 : _GEN_1164 ? ~_GEN_1784 & _GEN_112817 : ~(_GEN_112933 & _GEN_1784) & _GEN_112817) : _GEN_112817;
  wire        _GEN_113052 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1785 & _GEN_112818 : _GEN_1164 ? ~_GEN_1785 & _GEN_112818 : ~(_GEN_112933 & _GEN_1785) & _GEN_112818) : _GEN_112818;
  wire        _GEN_113053 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1786 & _GEN_112819 : _GEN_1164 ? ~_GEN_1786 & _GEN_112819 : ~(_GEN_112933 & _GEN_1786) & _GEN_112819) : _GEN_112819;
  wire        _GEN_113054 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1787 & _GEN_112820 : _GEN_1164 ? ~_GEN_1787 & _GEN_112820 : ~(_GEN_112933 & _GEN_1787) & _GEN_112820) : _GEN_112820;
  wire        _GEN_113055 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1788 & _GEN_112821 : _GEN_1164 ? ~_GEN_1788 & _GEN_112821 : ~(_GEN_112933 & _GEN_1788) & _GEN_112821) : _GEN_112821;
  wire        _GEN_113056 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1789 & _GEN_112822 : _GEN_1164 ? ~_GEN_1789 & _GEN_112822 : ~(_GEN_112933 & _GEN_1789) & _GEN_112822) : _GEN_112822;
  wire        _GEN_113057 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1790 & _GEN_112823 : _GEN_1164 ? ~_GEN_1790 & _GEN_112823 : ~(_GEN_112933 & _GEN_1790) & _GEN_112823) : _GEN_112823;
  wire        _GEN_113058 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1791 & _GEN_112824 : _GEN_1164 ? ~_GEN_1791 & _GEN_112824 : ~(_GEN_112933 & _GEN_1791) & _GEN_112824) : _GEN_112824;
  wire        _GEN_113059 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1792 & _GEN_112825 : _GEN_1164 ? ~_GEN_1792 & _GEN_112825 : ~(_GEN_112933 & _GEN_1792) & _GEN_112825) : _GEN_112825;
  wire        _GEN_113060 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1793 & _GEN_112826 : _GEN_1164 ? ~_GEN_1793 & _GEN_112826 : ~(_GEN_112933 & _GEN_1793) & _GEN_112826) : _GEN_112826;
  wire        _GEN_113061 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1794 & _GEN_112827 : _GEN_1164 ? ~_GEN_1794 & _GEN_112827 : ~(_GEN_112933 & _GEN_1794) & _GEN_112827) : _GEN_112827;
  wire        _GEN_113062 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1795 & _GEN_112828 : _GEN_1164 ? ~_GEN_1795 & _GEN_112828 : ~(_GEN_112933 & _GEN_1795) & _GEN_112828) : _GEN_112828;
  wire        _GEN_113063 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1796 & _GEN_112829 : _GEN_1164 ? ~_GEN_1796 & _GEN_112829 : ~(_GEN_112933 & _GEN_1796) & _GEN_112829) : _GEN_112829;
  wire        _GEN_113064 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1797 & _GEN_112830 : _GEN_1164 ? ~_GEN_1797 & _GEN_112830 : ~(_GEN_112933 & _GEN_1797) & _GEN_112830) : _GEN_112830;
  wire        _GEN_113065 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1798 & _GEN_112831 : _GEN_1164 ? ~_GEN_1798 & _GEN_112831 : ~(_GEN_112933 & _GEN_1798) & _GEN_112831) : _GEN_112831;
  wire        _GEN_113066 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1799 & _GEN_112832 : _GEN_1164 ? ~_GEN_1799 & _GEN_112832 : ~(_GEN_112933 & _GEN_1799) & _GEN_112832) : _GEN_112832;
  wire        _GEN_113067 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1800 & _GEN_112833 : _GEN_1164 ? ~_GEN_1800 & _GEN_112833 : ~(_GEN_112933 & _GEN_1800) & _GEN_112833) : _GEN_112833;
  wire        _GEN_113068 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1801 & _GEN_112834 : _GEN_1164 ? ~_GEN_1801 & _GEN_112834 : ~(_GEN_112933 & _GEN_1801) & _GEN_112834) : _GEN_112834;
  wire        _GEN_113069 = _GEN_1162 ? (_GEN_113002 ? ~_GEN_1802 & _GEN_112835 : _GEN_1164 ? ~_GEN_1802 & _GEN_112835 : ~(_GEN_112933 & _GEN_1802) & _GEN_112835) : _GEN_112835;
  wire        _GEN_113070 = _GEN_1162 ? (_GEN_113002 ? ~(&lcam_ldq_idx_1) & _GEN_112836 : _GEN_1164 ? ~(&lcam_ldq_idx_1) & _GEN_112836 : ~(_GEN_112933 & (&lcam_ldq_idx_1)) & _GEN_112836) : _GEN_112836;
  wire        _GEN_113273 = _GEN_1165 ? (_GEN_113236 ? (|lcam_ldq_idx_0) & _GEN_113039 : _GEN_1167 ? (|lcam_ldq_idx_0) & _GEN_113039 : ~(_GEN_113401 & ~(|lcam_ldq_idx_0)) & _GEN_113039) : _GEN_113039;
  wire        _GEN_113274 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1743 & _GEN_113040 : _GEN_1167 ? ~_GEN_1743 & _GEN_113040 : ~(_GEN_113401 & _GEN_1743) & _GEN_113040) : _GEN_113040;
  wire        _GEN_113275 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1744 & _GEN_113041 : _GEN_1167 ? ~_GEN_1744 & _GEN_113041 : ~(_GEN_113401 & _GEN_1744) & _GEN_113041) : _GEN_113041;
  wire        _GEN_113276 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1745 & _GEN_113042 : _GEN_1167 ? ~_GEN_1745 & _GEN_113042 : ~(_GEN_113401 & _GEN_1745) & _GEN_113042) : _GEN_113042;
  wire        _GEN_113277 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1746 & _GEN_113043 : _GEN_1167 ? ~_GEN_1746 & _GEN_113043 : ~(_GEN_113401 & _GEN_1746) & _GEN_113043) : _GEN_113043;
  wire        _GEN_113278 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1747 & _GEN_113044 : _GEN_1167 ? ~_GEN_1747 & _GEN_113044 : ~(_GEN_113401 & _GEN_1747) & _GEN_113044) : _GEN_113044;
  wire        _GEN_113279 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1748 & _GEN_113045 : _GEN_1167 ? ~_GEN_1748 & _GEN_113045 : ~(_GEN_113401 & _GEN_1748) & _GEN_113045) : _GEN_113045;
  wire        _GEN_113280 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1749 & _GEN_113046 : _GEN_1167 ? ~_GEN_1749 & _GEN_113046 : ~(_GEN_113401 & _GEN_1749) & _GEN_113046) : _GEN_113046;
  wire        _GEN_113281 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1750 & _GEN_113047 : _GEN_1167 ? ~_GEN_1750 & _GEN_113047 : ~(_GEN_113401 & _GEN_1750) & _GEN_113047) : _GEN_113047;
  wire        _GEN_113282 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1751 & _GEN_113048 : _GEN_1167 ? ~_GEN_1751 & _GEN_113048 : ~(_GEN_113401 & _GEN_1751) & _GEN_113048) : _GEN_113048;
  wire        _GEN_113283 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1752 & _GEN_113049 : _GEN_1167 ? ~_GEN_1752 & _GEN_113049 : ~(_GEN_113401 & _GEN_1752) & _GEN_113049) : _GEN_113049;
  wire        _GEN_113284 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1753 & _GEN_113050 : _GEN_1167 ? ~_GEN_1753 & _GEN_113050 : ~(_GEN_113401 & _GEN_1753) & _GEN_113050) : _GEN_113050;
  wire        _GEN_113285 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1754 & _GEN_113051 : _GEN_1167 ? ~_GEN_1754 & _GEN_113051 : ~(_GEN_113401 & _GEN_1754) & _GEN_113051) : _GEN_113051;
  wire        _GEN_113286 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1755 & _GEN_113052 : _GEN_1167 ? ~_GEN_1755 & _GEN_113052 : ~(_GEN_113401 & _GEN_1755) & _GEN_113052) : _GEN_113052;
  wire        _GEN_113287 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1756 & _GEN_113053 : _GEN_1167 ? ~_GEN_1756 & _GEN_113053 : ~(_GEN_113401 & _GEN_1756) & _GEN_113053) : _GEN_113053;
  wire        _GEN_113288 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1757 & _GEN_113054 : _GEN_1167 ? ~_GEN_1757 & _GEN_113054 : ~(_GEN_113401 & _GEN_1757) & _GEN_113054) : _GEN_113054;
  wire        _GEN_113289 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1758 & _GEN_113055 : _GEN_1167 ? ~_GEN_1758 & _GEN_113055 : ~(_GEN_113401 & _GEN_1758) & _GEN_113055) : _GEN_113055;
  wire        _GEN_113290 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1759 & _GEN_113056 : _GEN_1167 ? ~_GEN_1759 & _GEN_113056 : ~(_GEN_113401 & _GEN_1759) & _GEN_113056) : _GEN_113056;
  wire        _GEN_113291 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1760 & _GEN_113057 : _GEN_1167 ? ~_GEN_1760 & _GEN_113057 : ~(_GEN_113401 & _GEN_1760) & _GEN_113057) : _GEN_113057;
  wire        _GEN_113292 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1761 & _GEN_113058 : _GEN_1167 ? ~_GEN_1761 & _GEN_113058 : ~(_GEN_113401 & _GEN_1761) & _GEN_113058) : _GEN_113058;
  wire        _GEN_113293 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1762 & _GEN_113059 : _GEN_1167 ? ~_GEN_1762 & _GEN_113059 : ~(_GEN_113401 & _GEN_1762) & _GEN_113059) : _GEN_113059;
  wire        _GEN_113294 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1763 & _GEN_113060 : _GEN_1167 ? ~_GEN_1763 & _GEN_113060 : ~(_GEN_113401 & _GEN_1763) & _GEN_113060) : _GEN_113060;
  wire        _GEN_113295 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1764 & _GEN_113061 : _GEN_1167 ? ~_GEN_1764 & _GEN_113061 : ~(_GEN_113401 & _GEN_1764) & _GEN_113061) : _GEN_113061;
  wire        _GEN_113296 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1765 & _GEN_113062 : _GEN_1167 ? ~_GEN_1765 & _GEN_113062 : ~(_GEN_113401 & _GEN_1765) & _GEN_113062) : _GEN_113062;
  wire        _GEN_113297 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1766 & _GEN_113063 : _GEN_1167 ? ~_GEN_1766 & _GEN_113063 : ~(_GEN_113401 & _GEN_1766) & _GEN_113063) : _GEN_113063;
  wire        _GEN_113298 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1767 & _GEN_113064 : _GEN_1167 ? ~_GEN_1767 & _GEN_113064 : ~(_GEN_113401 & _GEN_1767) & _GEN_113064) : _GEN_113064;
  wire        _GEN_113299 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1768 & _GEN_113065 : _GEN_1167 ? ~_GEN_1768 & _GEN_113065 : ~(_GEN_113401 & _GEN_1768) & _GEN_113065) : _GEN_113065;
  wire        _GEN_113300 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1769 & _GEN_113066 : _GEN_1167 ? ~_GEN_1769 & _GEN_113066 : ~(_GEN_113401 & _GEN_1769) & _GEN_113066) : _GEN_113066;
  wire        _GEN_113301 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1770 & _GEN_113067 : _GEN_1167 ? ~_GEN_1770 & _GEN_113067 : ~(_GEN_113401 & _GEN_1770) & _GEN_113067) : _GEN_113067;
  wire        _GEN_113302 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1771 & _GEN_113068 : _GEN_1167 ? ~_GEN_1771 & _GEN_113068 : ~(_GEN_113401 & _GEN_1771) & _GEN_113068) : _GEN_113068;
  wire        _GEN_113303 = _GEN_1165 ? (_GEN_113236 ? ~_GEN_1772 & _GEN_113069 : _GEN_1167 ? ~_GEN_1772 & _GEN_113069 : ~(_GEN_113401 & _GEN_1772) & _GEN_113069) : _GEN_113069;
  wire        _GEN_113304 = _GEN_1165 ? (_GEN_113236 ? ~(&lcam_ldq_idx_0) & _GEN_113070 : _GEN_1167 ? ~(&lcam_ldq_idx_0) & _GEN_113070 : ~(_GEN_113401 & (&lcam_ldq_idx_0)) & _GEN_113070) : _GEN_113070;
  wire        _GEN_113507 = _GEN_1168 ? (_GEN_113470 ? (|lcam_ldq_idx_1) & _GEN_113273 : _GEN_1170 ? (|lcam_ldq_idx_1) & _GEN_113273 : ~(_GEN_113401 & ~(|lcam_ldq_idx_1)) & _GEN_113273) : _GEN_113273;
  wire        _GEN_113508 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1773 & _GEN_113274 : _GEN_1170 ? ~_GEN_1773 & _GEN_113274 : ~(_GEN_113401 & _GEN_1773) & _GEN_113274) : _GEN_113274;
  wire        _GEN_113509 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1774 & _GEN_113275 : _GEN_1170 ? ~_GEN_1774 & _GEN_113275 : ~(_GEN_113401 & _GEN_1774) & _GEN_113275) : _GEN_113275;
  wire        _GEN_113510 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1775 & _GEN_113276 : _GEN_1170 ? ~_GEN_1775 & _GEN_113276 : ~(_GEN_113401 & _GEN_1775) & _GEN_113276) : _GEN_113276;
  wire        _GEN_113511 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1776 & _GEN_113277 : _GEN_1170 ? ~_GEN_1776 & _GEN_113277 : ~(_GEN_113401 & _GEN_1776) & _GEN_113277) : _GEN_113277;
  wire        _GEN_113512 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1777 & _GEN_113278 : _GEN_1170 ? ~_GEN_1777 & _GEN_113278 : ~(_GEN_113401 & _GEN_1777) & _GEN_113278) : _GEN_113278;
  wire        _GEN_113513 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1778 & _GEN_113279 : _GEN_1170 ? ~_GEN_1778 & _GEN_113279 : ~(_GEN_113401 & _GEN_1778) & _GEN_113279) : _GEN_113279;
  wire        _GEN_113514 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1779 & _GEN_113280 : _GEN_1170 ? ~_GEN_1779 & _GEN_113280 : ~(_GEN_113401 & _GEN_1779) & _GEN_113280) : _GEN_113280;
  wire        _GEN_113515 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1780 & _GEN_113281 : _GEN_1170 ? ~_GEN_1780 & _GEN_113281 : ~(_GEN_113401 & _GEN_1780) & _GEN_113281) : _GEN_113281;
  wire        _GEN_113516 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1781 & _GEN_113282 : _GEN_1170 ? ~_GEN_1781 & _GEN_113282 : ~(_GEN_113401 & _GEN_1781) & _GEN_113282) : _GEN_113282;
  wire        _GEN_113517 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1782 & _GEN_113283 : _GEN_1170 ? ~_GEN_1782 & _GEN_113283 : ~(_GEN_113401 & _GEN_1782) & _GEN_113283) : _GEN_113283;
  wire        _GEN_113518 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1783 & _GEN_113284 : _GEN_1170 ? ~_GEN_1783 & _GEN_113284 : ~(_GEN_113401 & _GEN_1783) & _GEN_113284) : _GEN_113284;
  wire        _GEN_113519 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1784 & _GEN_113285 : _GEN_1170 ? ~_GEN_1784 & _GEN_113285 : ~(_GEN_113401 & _GEN_1784) & _GEN_113285) : _GEN_113285;
  wire        _GEN_113520 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1785 & _GEN_113286 : _GEN_1170 ? ~_GEN_1785 & _GEN_113286 : ~(_GEN_113401 & _GEN_1785) & _GEN_113286) : _GEN_113286;
  wire        _GEN_113521 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1786 & _GEN_113287 : _GEN_1170 ? ~_GEN_1786 & _GEN_113287 : ~(_GEN_113401 & _GEN_1786) & _GEN_113287) : _GEN_113287;
  wire        _GEN_113522 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1787 & _GEN_113288 : _GEN_1170 ? ~_GEN_1787 & _GEN_113288 : ~(_GEN_113401 & _GEN_1787) & _GEN_113288) : _GEN_113288;
  wire        _GEN_113523 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1788 & _GEN_113289 : _GEN_1170 ? ~_GEN_1788 & _GEN_113289 : ~(_GEN_113401 & _GEN_1788) & _GEN_113289) : _GEN_113289;
  wire        _GEN_113524 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1789 & _GEN_113290 : _GEN_1170 ? ~_GEN_1789 & _GEN_113290 : ~(_GEN_113401 & _GEN_1789) & _GEN_113290) : _GEN_113290;
  wire        _GEN_113525 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1790 & _GEN_113291 : _GEN_1170 ? ~_GEN_1790 & _GEN_113291 : ~(_GEN_113401 & _GEN_1790) & _GEN_113291) : _GEN_113291;
  wire        _GEN_113526 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1791 & _GEN_113292 : _GEN_1170 ? ~_GEN_1791 & _GEN_113292 : ~(_GEN_113401 & _GEN_1791) & _GEN_113292) : _GEN_113292;
  wire        _GEN_113527 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1792 & _GEN_113293 : _GEN_1170 ? ~_GEN_1792 & _GEN_113293 : ~(_GEN_113401 & _GEN_1792) & _GEN_113293) : _GEN_113293;
  wire        _GEN_113528 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1793 & _GEN_113294 : _GEN_1170 ? ~_GEN_1793 & _GEN_113294 : ~(_GEN_113401 & _GEN_1793) & _GEN_113294) : _GEN_113294;
  wire        _GEN_113529 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1794 & _GEN_113295 : _GEN_1170 ? ~_GEN_1794 & _GEN_113295 : ~(_GEN_113401 & _GEN_1794) & _GEN_113295) : _GEN_113295;
  wire        _GEN_113530 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1795 & _GEN_113296 : _GEN_1170 ? ~_GEN_1795 & _GEN_113296 : ~(_GEN_113401 & _GEN_1795) & _GEN_113296) : _GEN_113296;
  wire        _GEN_113531 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1796 & _GEN_113297 : _GEN_1170 ? ~_GEN_1796 & _GEN_113297 : ~(_GEN_113401 & _GEN_1796) & _GEN_113297) : _GEN_113297;
  wire        _GEN_113532 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1797 & _GEN_113298 : _GEN_1170 ? ~_GEN_1797 & _GEN_113298 : ~(_GEN_113401 & _GEN_1797) & _GEN_113298) : _GEN_113298;
  wire        _GEN_113533 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1798 & _GEN_113299 : _GEN_1170 ? ~_GEN_1798 & _GEN_113299 : ~(_GEN_113401 & _GEN_1798) & _GEN_113299) : _GEN_113299;
  wire        _GEN_113534 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1799 & _GEN_113300 : _GEN_1170 ? ~_GEN_1799 & _GEN_113300 : ~(_GEN_113401 & _GEN_1799) & _GEN_113300) : _GEN_113300;
  wire        _GEN_113535 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1800 & _GEN_113301 : _GEN_1170 ? ~_GEN_1800 & _GEN_113301 : ~(_GEN_113401 & _GEN_1800) & _GEN_113301) : _GEN_113301;
  wire        _GEN_113536 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1801 & _GEN_113302 : _GEN_1170 ? ~_GEN_1801 & _GEN_113302 : ~(_GEN_113401 & _GEN_1801) & _GEN_113302) : _GEN_113302;
  wire        _GEN_113537 = _GEN_1168 ? (_GEN_113470 ? ~_GEN_1802 & _GEN_113303 : _GEN_1170 ? ~_GEN_1802 & _GEN_113303 : ~(_GEN_113401 & _GEN_1802) & _GEN_113303) : _GEN_113303;
  wire        _GEN_113538 = _GEN_1168 ? (_GEN_113470 ? ~(&lcam_ldq_idx_1) & _GEN_113304 : _GEN_1170 ? ~(&lcam_ldq_idx_1) & _GEN_113304 : ~(_GEN_113401 & (&lcam_ldq_idx_1)) & _GEN_113304) : _GEN_113304;
  wire        _GEN_113741 = _GEN_1171 ? (_GEN_113704 ? (|lcam_ldq_idx_0) & _GEN_113507 : _GEN_1173 ? (|lcam_ldq_idx_0) & _GEN_113507 : ~(_GEN_113869 & ~(|lcam_ldq_idx_0)) & _GEN_113507) : _GEN_113507;
  wire        _GEN_113742 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1743 & _GEN_113508 : _GEN_1173 ? ~_GEN_1743 & _GEN_113508 : ~(_GEN_113869 & _GEN_1743) & _GEN_113508) : _GEN_113508;
  wire        _GEN_113743 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1744 & _GEN_113509 : _GEN_1173 ? ~_GEN_1744 & _GEN_113509 : ~(_GEN_113869 & _GEN_1744) & _GEN_113509) : _GEN_113509;
  wire        _GEN_113744 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1745 & _GEN_113510 : _GEN_1173 ? ~_GEN_1745 & _GEN_113510 : ~(_GEN_113869 & _GEN_1745) & _GEN_113510) : _GEN_113510;
  wire        _GEN_113745 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1746 & _GEN_113511 : _GEN_1173 ? ~_GEN_1746 & _GEN_113511 : ~(_GEN_113869 & _GEN_1746) & _GEN_113511) : _GEN_113511;
  wire        _GEN_113746 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1747 & _GEN_113512 : _GEN_1173 ? ~_GEN_1747 & _GEN_113512 : ~(_GEN_113869 & _GEN_1747) & _GEN_113512) : _GEN_113512;
  wire        _GEN_113747 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1748 & _GEN_113513 : _GEN_1173 ? ~_GEN_1748 & _GEN_113513 : ~(_GEN_113869 & _GEN_1748) & _GEN_113513) : _GEN_113513;
  wire        _GEN_113748 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1749 & _GEN_113514 : _GEN_1173 ? ~_GEN_1749 & _GEN_113514 : ~(_GEN_113869 & _GEN_1749) & _GEN_113514) : _GEN_113514;
  wire        _GEN_113749 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1750 & _GEN_113515 : _GEN_1173 ? ~_GEN_1750 & _GEN_113515 : ~(_GEN_113869 & _GEN_1750) & _GEN_113515) : _GEN_113515;
  wire        _GEN_113750 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1751 & _GEN_113516 : _GEN_1173 ? ~_GEN_1751 & _GEN_113516 : ~(_GEN_113869 & _GEN_1751) & _GEN_113516) : _GEN_113516;
  wire        _GEN_113751 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1752 & _GEN_113517 : _GEN_1173 ? ~_GEN_1752 & _GEN_113517 : ~(_GEN_113869 & _GEN_1752) & _GEN_113517) : _GEN_113517;
  wire        _GEN_113752 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1753 & _GEN_113518 : _GEN_1173 ? ~_GEN_1753 & _GEN_113518 : ~(_GEN_113869 & _GEN_1753) & _GEN_113518) : _GEN_113518;
  wire        _GEN_113753 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1754 & _GEN_113519 : _GEN_1173 ? ~_GEN_1754 & _GEN_113519 : ~(_GEN_113869 & _GEN_1754) & _GEN_113519) : _GEN_113519;
  wire        _GEN_113754 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1755 & _GEN_113520 : _GEN_1173 ? ~_GEN_1755 & _GEN_113520 : ~(_GEN_113869 & _GEN_1755) & _GEN_113520) : _GEN_113520;
  wire        _GEN_113755 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1756 & _GEN_113521 : _GEN_1173 ? ~_GEN_1756 & _GEN_113521 : ~(_GEN_113869 & _GEN_1756) & _GEN_113521) : _GEN_113521;
  wire        _GEN_113756 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1757 & _GEN_113522 : _GEN_1173 ? ~_GEN_1757 & _GEN_113522 : ~(_GEN_113869 & _GEN_1757) & _GEN_113522) : _GEN_113522;
  wire        _GEN_113757 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1758 & _GEN_113523 : _GEN_1173 ? ~_GEN_1758 & _GEN_113523 : ~(_GEN_113869 & _GEN_1758) & _GEN_113523) : _GEN_113523;
  wire        _GEN_113758 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1759 & _GEN_113524 : _GEN_1173 ? ~_GEN_1759 & _GEN_113524 : ~(_GEN_113869 & _GEN_1759) & _GEN_113524) : _GEN_113524;
  wire        _GEN_113759 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1760 & _GEN_113525 : _GEN_1173 ? ~_GEN_1760 & _GEN_113525 : ~(_GEN_113869 & _GEN_1760) & _GEN_113525) : _GEN_113525;
  wire        _GEN_113760 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1761 & _GEN_113526 : _GEN_1173 ? ~_GEN_1761 & _GEN_113526 : ~(_GEN_113869 & _GEN_1761) & _GEN_113526) : _GEN_113526;
  wire        _GEN_113761 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1762 & _GEN_113527 : _GEN_1173 ? ~_GEN_1762 & _GEN_113527 : ~(_GEN_113869 & _GEN_1762) & _GEN_113527) : _GEN_113527;
  wire        _GEN_113762 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1763 & _GEN_113528 : _GEN_1173 ? ~_GEN_1763 & _GEN_113528 : ~(_GEN_113869 & _GEN_1763) & _GEN_113528) : _GEN_113528;
  wire        _GEN_113763 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1764 & _GEN_113529 : _GEN_1173 ? ~_GEN_1764 & _GEN_113529 : ~(_GEN_113869 & _GEN_1764) & _GEN_113529) : _GEN_113529;
  wire        _GEN_113764 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1765 & _GEN_113530 : _GEN_1173 ? ~_GEN_1765 & _GEN_113530 : ~(_GEN_113869 & _GEN_1765) & _GEN_113530) : _GEN_113530;
  wire        _GEN_113765 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1766 & _GEN_113531 : _GEN_1173 ? ~_GEN_1766 & _GEN_113531 : ~(_GEN_113869 & _GEN_1766) & _GEN_113531) : _GEN_113531;
  wire        _GEN_113766 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1767 & _GEN_113532 : _GEN_1173 ? ~_GEN_1767 & _GEN_113532 : ~(_GEN_113869 & _GEN_1767) & _GEN_113532) : _GEN_113532;
  wire        _GEN_113767 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1768 & _GEN_113533 : _GEN_1173 ? ~_GEN_1768 & _GEN_113533 : ~(_GEN_113869 & _GEN_1768) & _GEN_113533) : _GEN_113533;
  wire        _GEN_113768 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1769 & _GEN_113534 : _GEN_1173 ? ~_GEN_1769 & _GEN_113534 : ~(_GEN_113869 & _GEN_1769) & _GEN_113534) : _GEN_113534;
  wire        _GEN_113769 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1770 & _GEN_113535 : _GEN_1173 ? ~_GEN_1770 & _GEN_113535 : ~(_GEN_113869 & _GEN_1770) & _GEN_113535) : _GEN_113535;
  wire        _GEN_113770 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1771 & _GEN_113536 : _GEN_1173 ? ~_GEN_1771 & _GEN_113536 : ~(_GEN_113869 & _GEN_1771) & _GEN_113536) : _GEN_113536;
  wire        _GEN_113771 = _GEN_1171 ? (_GEN_113704 ? ~_GEN_1772 & _GEN_113537 : _GEN_1173 ? ~_GEN_1772 & _GEN_113537 : ~(_GEN_113869 & _GEN_1772) & _GEN_113537) : _GEN_113537;
  wire        _GEN_113772 = _GEN_1171 ? (_GEN_113704 ? ~(&lcam_ldq_idx_0) & _GEN_113538 : _GEN_1173 ? ~(&lcam_ldq_idx_0) & _GEN_113538 : ~(_GEN_113869 & (&lcam_ldq_idx_0)) & _GEN_113538) : _GEN_113538;
  wire        ld_xcpt_valid = failed_loads_0 | failed_loads_1 | failed_loads_2 | failed_loads_3 | failed_loads_4 | failed_loads_5 | failed_loads_6 | failed_loads_7 | failed_loads_8 | failed_loads_9 | failed_loads_10 | failed_loads_11 | failed_loads_12 | failed_loads_13 | failed_loads_14 | failed_loads_15 | failed_loads_16 | failed_loads_17 | failed_loads_18 | failed_loads_19 | failed_loads_20 | failed_loads_21 | failed_loads_22 | failed_loads_23 | failed_loads_24 | failed_loads_25 | failed_loads_26 | failed_loads_27 | failed_loads_28 | failed_loads_29 | failed_loads_30 | failed_loads_31;
  wire        use_mem_xcpt = mem_xcpt_valid & (mem_xcpt_uop_rob_idx < casez_tmp_178 ^ mem_xcpt_uop_rob_idx < io_core_rob_head_idx ^ casez_tmp_178 < io_core_rob_head_idx) | ~ld_xcpt_valid;
  wire [19:0] xcpt_uop_br_mask = use_mem_xcpt ? (is_older ? mem_xcpt_uops_1_br_mask : mem_xcpt_uops_0_br_mask) : casez_tmp_179;
  wire        _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded = _io_core_exe_0_iresp_valid_output | _io_core_exe_0_fresp_valid_output;
  wire        _GEN_1867 = casez_tmp_203 & live;
  wire        _GEN_1868 = _GEN_1180 & _GEN_1867 & ~(|wb_forward_ldq_idx_0);
  wire        _GEN_1869 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h1;
  wire        _GEN_1870 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h2;
  wire        _GEN_1871 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h3;
  wire        _GEN_1872 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h4;
  wire        _GEN_1873 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h5;
  wire        _GEN_1874 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h6;
  wire        _GEN_1875 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h7;
  wire        _GEN_1876 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h8;
  wire        _GEN_1877 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h9;
  wire        _GEN_1878 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'hA;
  wire        _GEN_1879 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'hB;
  wire        _GEN_1880 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'hC;
  wire        _GEN_1881 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'hD;
  wire        _GEN_1882 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'hE;
  wire        _GEN_1883 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'hF;
  wire        _GEN_1884 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h10;
  wire        _GEN_1885 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h11;
  wire        _GEN_1886 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h12;
  wire        _GEN_1887 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h13;
  wire        _GEN_1888 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h14;
  wire        _GEN_1889 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h15;
  wire        _GEN_1890 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h16;
  wire        _GEN_1891 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h17;
  wire        _GEN_1892 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h18;
  wire        _GEN_1893 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h19;
  wire        _GEN_1894 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h1A;
  wire        _GEN_1895 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h1B;
  wire        _GEN_1896 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h1C;
  wire        _GEN_1897 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h1D;
  wire        _GEN_1898 = _GEN_1180 & _GEN_1867 & wb_forward_ldq_idx_0 == 5'h1E;
  wire        _GEN_1899 = _GEN_1180 & _GEN_1867 & (&wb_forward_ldq_idx_0);
  wire        _GEN_1900 = _GEN_1179 | ~_GEN_1868;
  wire        _GEN_1901 = _GEN_1179 | ~_GEN_1869;
  wire        _GEN_1902 = _GEN_1179 | ~_GEN_1870;
  wire        _GEN_1903 = _GEN_1179 | ~_GEN_1871;
  wire        _GEN_1904 = _GEN_1179 | ~_GEN_1872;
  wire        _GEN_1905 = _GEN_1179 | ~_GEN_1873;
  wire        _GEN_1906 = _GEN_1179 | ~_GEN_1874;
  wire        _GEN_1907 = _GEN_1179 | ~_GEN_1875;
  wire        _GEN_1908 = _GEN_1179 | ~_GEN_1876;
  wire        _GEN_1909 = _GEN_1179 | ~_GEN_1877;
  wire        _GEN_1910 = _GEN_1179 | ~_GEN_1878;
  wire        _GEN_1911 = _GEN_1179 | ~_GEN_1879;
  wire        _GEN_1912 = _GEN_1179 | ~_GEN_1880;
  wire        _GEN_1913 = _GEN_1179 | ~_GEN_1881;
  wire        _GEN_1914 = _GEN_1179 | ~_GEN_1882;
  wire        _GEN_1915 = _GEN_1179 | ~_GEN_1883;
  wire        _GEN_1916 = _GEN_1179 | ~_GEN_1884;
  wire        _GEN_1917 = _GEN_1179 | ~_GEN_1885;
  wire        _GEN_1918 = _GEN_1179 | ~_GEN_1886;
  wire        _GEN_1919 = _GEN_1179 | ~_GEN_1887;
  wire        _GEN_1920 = _GEN_1179 | ~_GEN_1888;
  wire        _GEN_1921 = _GEN_1179 | ~_GEN_1889;
  wire        _GEN_1922 = _GEN_1179 | ~_GEN_1890;
  wire        _GEN_1923 = _GEN_1179 | ~_GEN_1891;
  wire        _GEN_1924 = _GEN_1179 | ~_GEN_1892;
  wire        _GEN_1925 = _GEN_1179 | ~_GEN_1893;
  wire        _GEN_1926 = _GEN_1179 | ~_GEN_1894;
  wire        _GEN_1927 = _GEN_1179 | ~_GEN_1895;
  wire        _GEN_1928 = _GEN_1179 | ~_GEN_1896;
  wire        _GEN_1929 = _GEN_1179 | ~_GEN_1897;
  wire        _GEN_1930 = _GEN_1179 | ~_GEN_1898;
  wire        _GEN_1931 = _GEN_1179 | ~_GEN_1899;
  wire        _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded = _io_core_exe_1_iresp_valid_output | _io_core_exe_1_fresp_valid_output;
  wire        _GEN_1932 = casez_tmp_236 & live_1;
  wire        _GEN_1933 = _GEN_1184 & _GEN_1932 & ~(|wb_forward_ldq_idx_1);
  wire        _GEN_1934 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h1;
  wire        _GEN_1935 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h2;
  wire        _GEN_1936 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h3;
  wire        _GEN_1937 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h4;
  wire        _GEN_1938 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h5;
  wire        _GEN_1939 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h6;
  wire        _GEN_1940 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h7;
  wire        _GEN_1941 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h8;
  wire        _GEN_1942 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h9;
  wire        _GEN_1943 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'hA;
  wire        _GEN_1944 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'hB;
  wire        _GEN_1945 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'hC;
  wire        _GEN_1946 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'hD;
  wire        _GEN_1947 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'hE;
  wire        _GEN_1948 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'hF;
  wire        _GEN_1949 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h10;
  wire        _GEN_1950 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h11;
  wire        _GEN_1951 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h12;
  wire        _GEN_1952 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h13;
  wire        _GEN_1953 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h14;
  wire        _GEN_1954 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h15;
  wire        _GEN_1955 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h16;
  wire        _GEN_1956 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h17;
  wire        _GEN_1957 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h18;
  wire        _GEN_1958 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h19;
  wire        _GEN_1959 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h1A;
  wire        _GEN_1960 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h1B;
  wire        _GEN_1961 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h1C;
  wire        _GEN_1962 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h1D;
  wire        _GEN_1963 = _GEN_1184 & _GEN_1932 & wb_forward_ldq_idx_1 == 5'h1E;
  wire        _GEN_1964 = _GEN_1184 & _GEN_1932 & (&wb_forward_ldq_idx_1);
  wire        _GEN_1965 = _GEN_1183 | ~_GEN_1933;
  wire        _GEN_1966 = _GEN_1183 | ~_GEN_1934;
  wire        _GEN_1967 = _GEN_1183 | ~_GEN_1935;
  wire        _GEN_1968 = _GEN_1183 | ~_GEN_1936;
  wire        _GEN_1969 = _GEN_1183 | ~_GEN_1937;
  wire        _GEN_1970 = _GEN_1183 | ~_GEN_1938;
  wire        _GEN_1971 = _GEN_1183 | ~_GEN_1939;
  wire        _GEN_1972 = _GEN_1183 | ~_GEN_1940;
  wire        _GEN_1973 = _GEN_1183 | ~_GEN_1941;
  wire        _GEN_1974 = _GEN_1183 | ~_GEN_1942;
  wire        _GEN_1975 = _GEN_1183 | ~_GEN_1943;
  wire        _GEN_1976 = _GEN_1183 | ~_GEN_1944;
  wire        _GEN_1977 = _GEN_1183 | ~_GEN_1945;
  wire        _GEN_1978 = _GEN_1183 | ~_GEN_1946;
  wire        _GEN_1979 = _GEN_1183 | ~_GEN_1947;
  wire        _GEN_1980 = _GEN_1183 | ~_GEN_1948;
  wire        _GEN_1981 = _GEN_1183 | ~_GEN_1949;
  wire        _GEN_1982 = _GEN_1183 | ~_GEN_1950;
  wire        _GEN_1983 = _GEN_1183 | ~_GEN_1951;
  wire        _GEN_1984 = _GEN_1183 | ~_GEN_1952;
  wire        _GEN_1985 = _GEN_1183 | ~_GEN_1953;
  wire        _GEN_1986 = _GEN_1183 | ~_GEN_1954;
  wire        _GEN_1987 = _GEN_1183 | ~_GEN_1955;
  wire        _GEN_1988 = _GEN_1183 | ~_GEN_1956;
  wire        _GEN_1989 = _GEN_1183 | ~_GEN_1957;
  wire        _GEN_1990 = _GEN_1183 | ~_GEN_1958;
  wire        _GEN_1991 = _GEN_1183 | ~_GEN_1959;
  wire        _GEN_1992 = _GEN_1183 | ~_GEN_1960;
  wire        _GEN_1993 = _GEN_1183 | ~_GEN_1961;
  wire        _GEN_1994 = _GEN_1183 | ~_GEN_1962;
  wire        _GEN_1995 = _GEN_1183 | ~_GEN_1963;
  wire        _GEN_1996 = _GEN_1183 | ~_GEN_1964;
  wire        _GEN_1997 = stq_0_valid & (|_GEN_1186);
  wire        _GEN_1998 = stq_1_valid & (|_GEN_1187);
  wire        _GEN_1999 = stq_2_valid & (|_GEN_1188);
  wire        _GEN_2000 = stq_3_valid & (|_GEN_1189);
  wire        _GEN_2001 = stq_4_valid & (|_GEN_1190);
  wire        _GEN_2002 = stq_5_valid & (|_GEN_1191);
  wire        _GEN_2003 = stq_6_valid & (|_GEN_1192);
  wire        _GEN_2004 = stq_7_valid & (|_GEN_1193);
  wire        _GEN_2005 = stq_8_valid & (|_GEN_1194);
  wire        _GEN_2006 = stq_9_valid & (|_GEN_1195);
  wire        _GEN_2007 = stq_10_valid & (|_GEN_1196);
  wire        _GEN_2008 = stq_11_valid & (|_GEN_1197);
  wire        _GEN_2009 = stq_12_valid & (|_GEN_1198);
  wire        _GEN_2010 = stq_13_valid & (|_GEN_1199);
  wire        _GEN_2011 = stq_14_valid & (|_GEN_1200);
  wire        _GEN_2012 = stq_15_valid & (|_GEN_1201);
  wire        _GEN_2013 = stq_16_valid & (|_GEN_1202);
  wire        _GEN_2014 = stq_17_valid & (|_GEN_1203);
  wire        _GEN_2015 = stq_18_valid & (|_GEN_1204);
  wire        _GEN_2016 = stq_19_valid & (|_GEN_1205);
  wire        _GEN_2017 = stq_20_valid & (|_GEN_1206);
  wire        _GEN_2018 = stq_21_valid & (|_GEN_1207);
  wire        _GEN_2019 = stq_22_valid & (|_GEN_1208);
  wire        _GEN_2020 = stq_23_valid & (|_GEN_1209);
  wire        _GEN_2021 = stq_24_valid & (|_GEN_1210);
  wire        _GEN_2022 = stq_25_valid & (|_GEN_1211);
  wire        _GEN_2023 = stq_26_valid & (|_GEN_1212);
  wire        _GEN_2024 = stq_27_valid & (|_GEN_1213);
  wire        _GEN_2025 = stq_28_valid & (|_GEN_1214);
  wire        _GEN_2026 = stq_29_valid & (|_GEN_1215);
  wire        _GEN_2027 = stq_30_valid & (|_GEN_1216);
  wire        _GEN_2028 = stq_31_valid & (|_GEN_1217);
  wire        _GEN_2029 = ldq_0_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_0_bits_uop_br_mask));
  wire        _GEN_2030 = ldq_1_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_1_bits_uop_br_mask));
  wire        _GEN_2031 = ldq_2_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_2_bits_uop_br_mask));
  wire        _GEN_2032 = ldq_3_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_3_bits_uop_br_mask));
  wire        _GEN_2033 = ldq_4_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_4_bits_uop_br_mask));
  wire        _GEN_2034 = ldq_5_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_5_bits_uop_br_mask));
  wire        _GEN_2035 = ldq_6_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_6_bits_uop_br_mask));
  wire        _GEN_2036 = ldq_7_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_7_bits_uop_br_mask));
  wire        _GEN_2037 = ldq_8_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_8_bits_uop_br_mask));
  wire        _GEN_2038 = ldq_9_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_9_bits_uop_br_mask));
  wire        _GEN_2039 = ldq_10_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_10_bits_uop_br_mask));
  wire        _GEN_2040 = ldq_11_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_11_bits_uop_br_mask));
  wire        _GEN_2041 = ldq_12_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_12_bits_uop_br_mask));
  wire        _GEN_2042 = ldq_13_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_13_bits_uop_br_mask));
  wire        _GEN_2043 = ldq_14_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_14_bits_uop_br_mask));
  wire        _GEN_2044 = ldq_15_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_15_bits_uop_br_mask));
  wire        _GEN_2045 = ldq_16_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_16_bits_uop_br_mask));
  wire        _GEN_2046 = ldq_17_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_17_bits_uop_br_mask));
  wire        _GEN_2047 = ldq_18_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_18_bits_uop_br_mask));
  wire        _GEN_2048 = ldq_19_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_19_bits_uop_br_mask));
  wire        _GEN_2049 = ldq_20_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_20_bits_uop_br_mask));
  wire        _GEN_2050 = ldq_21_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_21_bits_uop_br_mask));
  wire        _GEN_2051 = ldq_22_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_22_bits_uop_br_mask));
  wire        _GEN_2052 = ldq_23_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_23_bits_uop_br_mask));
  wire        _GEN_2053 = ldq_24_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_24_bits_uop_br_mask));
  wire        _GEN_2054 = ldq_25_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_25_bits_uop_br_mask));
  wire        _GEN_2055 = ldq_26_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_26_bits_uop_br_mask));
  wire        _GEN_2056 = ldq_27_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_27_bits_uop_br_mask));
  wire        _GEN_2057 = ldq_28_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_28_bits_uop_br_mask));
  wire        _GEN_2058 = ldq_29_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_29_bits_uop_br_mask));
  wire        _GEN_2059 = ldq_30_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_30_bits_uop_br_mask));
  wire        _GEN_2060 = ldq_31_valid & (|(io_core_brupdate_b1_mispredict_mask & ldq_31_bits_uop_br_mask));
  wire        _GEN_2061 = idx == 5'h0;
  wire        _GEN_2062 = idx == 5'h1;
  wire        _GEN_2063 = idx == 5'h2;
  wire        _GEN_2064 = idx == 5'h3;
  wire        _GEN_2065 = idx == 5'h4;
  wire        _GEN_2066 = idx == 5'h5;
  wire        _GEN_2067 = idx == 5'h6;
  wire        _GEN_2068 = idx == 5'h7;
  wire        _GEN_2069 = idx == 5'h8;
  wire        _GEN_2070 = idx == 5'h9;
  wire        _GEN_2071 = idx == 5'hA;
  wire        _GEN_2072 = idx == 5'hB;
  wire        _GEN_2073 = idx == 5'hC;
  wire        _GEN_2074 = idx == 5'hD;
  wire        _GEN_2075 = idx == 5'hE;
  wire        _GEN_2076 = idx == 5'hF;
  wire        _GEN_2077 = idx == 5'h10;
  wire        _GEN_2078 = idx == 5'h11;
  wire        _GEN_2079 = idx == 5'h12;
  wire        _GEN_2080 = idx == 5'h13;
  wire        _GEN_2081 = idx == 5'h14;
  wire        _GEN_2082 = idx == 5'h15;
  wire        _GEN_2083 = idx == 5'h16;
  wire        _GEN_2084 = idx == 5'h17;
  wire        _GEN_2085 = idx == 5'h18;
  wire        _GEN_2086 = idx == 5'h19;
  wire        _GEN_2087 = idx == 5'h1A;
  wire        _GEN_2088 = idx == 5'h1B;
  wire        _GEN_2089 = idx == 5'h1C;
  wire        _GEN_2090 = idx == 5'h1D;
  wire        _GEN_2091 = idx == 5'h1E;
  wire        _GEN_2092 = _GEN_2061 | _GEN_2029;
  wire        _GEN_2093 = _GEN_2062 | _GEN_2030;
  wire        _GEN_2094 = _GEN_2063 | _GEN_2031;
  wire        _GEN_2095 = _GEN_2064 | _GEN_2032;
  wire        _GEN_2096 = _GEN_2065 | _GEN_2033;
  wire        _GEN_2097 = _GEN_2066 | _GEN_2034;
  wire        _GEN_2098 = _GEN_2067 | _GEN_2035;
  wire        _GEN_2099 = _GEN_2068 | _GEN_2036;
  wire        _GEN_2100 = _GEN_2069 | _GEN_2037;
  wire        _GEN_2101 = _GEN_2070 | _GEN_2038;
  wire        _GEN_2102 = _GEN_2071 | _GEN_2039;
  wire        _GEN_2103 = _GEN_2072 | _GEN_2040;
  wire        _GEN_2104 = _GEN_2073 | _GEN_2041;
  wire        _GEN_2105 = _GEN_2074 | _GEN_2042;
  wire        _GEN_2106 = _GEN_2075 | _GEN_2043;
  wire        _GEN_2107 = _GEN_2076 | _GEN_2044;
  wire        _GEN_2108 = _GEN_2077 | _GEN_2045;
  wire        _GEN_2109 = _GEN_2078 | _GEN_2046;
  wire        _GEN_2110 = _GEN_2079 | _GEN_2047;
  wire        _GEN_2111 = _GEN_2080 | _GEN_2048;
  wire        _GEN_2112 = _GEN_2081 | _GEN_2049;
  wire        _GEN_2113 = _GEN_2082 | _GEN_2050;
  wire        _GEN_2114 = _GEN_2083 | _GEN_2051;
  wire        _GEN_2115 = _GEN_2084 | _GEN_2052;
  wire        _GEN_2116 = _GEN_2085 | _GEN_2053;
  wire        _GEN_2117 = _GEN_2086 | _GEN_2054;
  wire        _GEN_2118 = _GEN_2087 | _GEN_2055;
  wire        _GEN_2119 = _GEN_2088 | _GEN_2056;
  wire        _GEN_2120 = _GEN_2089 | _GEN_2057;
  wire        _GEN_2121 = _GEN_2090 | _GEN_2058;
  wire        _GEN_2122 = _GEN_2091 | _GEN_2059;
  wire        _GEN_2123 = (&idx) | _GEN_2060;
  wire        _GEN_2124 = commit_store & _GEN_2061;
  wire        _GEN_2125 = commit_store & _GEN_2062;
  wire        _GEN_2126 = commit_store & _GEN_2063;
  wire        _GEN_2127 = commit_store & _GEN_2064;
  wire        _GEN_2128 = commit_store & _GEN_2065;
  wire        _GEN_2129 = commit_store & _GEN_2066;
  wire        _GEN_2130 = commit_store & _GEN_2067;
  wire        _GEN_2131 = commit_store & _GEN_2068;
  wire        _GEN_2132 = commit_store & _GEN_2069;
  wire        _GEN_2133 = commit_store & _GEN_2070;
  wire        _GEN_2134 = commit_store & _GEN_2071;
  wire        _GEN_2135 = commit_store & _GEN_2072;
  wire        _GEN_2136 = commit_store & _GEN_2073;
  wire        _GEN_2137 = commit_store & _GEN_2074;
  wire        _GEN_2138 = commit_store & _GEN_2075;
  wire        _GEN_2139 = commit_store & _GEN_2076;
  wire        _GEN_2140 = commit_store & _GEN_2077;
  wire        _GEN_2141 = commit_store & _GEN_2078;
  wire        _GEN_2142 = commit_store & _GEN_2079;
  wire        _GEN_2143 = commit_store & _GEN_2080;
  wire        _GEN_2144 = commit_store & _GEN_2081;
  wire        _GEN_2145 = commit_store & _GEN_2082;
  wire        _GEN_2146 = commit_store & _GEN_2083;
  wire        _GEN_2147 = commit_store & _GEN_2084;
  wire        _GEN_2148 = commit_store & _GEN_2085;
  wire        _GEN_2149 = commit_store & _GEN_2086;
  wire        _GEN_2150 = commit_store & _GEN_2087;
  wire        _GEN_2151 = commit_store & _GEN_2088;
  wire        _GEN_2152 = commit_store & _GEN_2089;
  wire        _GEN_2153 = commit_store & _GEN_2090;
  wire        _GEN_2154 = commit_store & _GEN_2091;
  wire        _GEN_2155 = commit_store & (&idx);
  wire        _GEN_2156 = commit_store | ~commit_load;
  wire        _GEN_2157 = commit_store | ~(commit_load & _GEN_2061);
  wire        _GEN_2158 = commit_store | ~(commit_load & _GEN_2062);
  wire        _GEN_2159 = commit_store | ~(commit_load & _GEN_2063);
  wire        _GEN_2160 = commit_store | ~(commit_load & _GEN_2064);
  wire        _GEN_2161 = commit_store | ~(commit_load & _GEN_2065);
  wire        _GEN_2162 = commit_store | ~(commit_load & _GEN_2066);
  wire        _GEN_2163 = commit_store | ~(commit_load & _GEN_2067);
  wire        _GEN_2164 = commit_store | ~(commit_load & _GEN_2068);
  wire        _GEN_2165 = commit_store | ~(commit_load & _GEN_2069);
  wire        _GEN_2166 = commit_store | ~(commit_load & _GEN_2070);
  wire        _GEN_2167 = commit_store | ~(commit_load & _GEN_2071);
  wire        _GEN_2168 = commit_store | ~(commit_load & _GEN_2072);
  wire        _GEN_2169 = commit_store | ~(commit_load & _GEN_2073);
  wire        _GEN_2170 = commit_store | ~(commit_load & _GEN_2074);
  wire        _GEN_2171 = commit_store | ~(commit_load & _GEN_2075);
  wire        _GEN_2172 = commit_store | ~(commit_load & _GEN_2076);
  wire        _GEN_2173 = commit_store | ~(commit_load & _GEN_2077);
  wire        _GEN_2174 = commit_store | ~(commit_load & _GEN_2078);
  wire        _GEN_2175 = commit_store | ~(commit_load & _GEN_2079);
  wire        _GEN_2176 = commit_store | ~(commit_load & _GEN_2080);
  wire        _GEN_2177 = commit_store | ~(commit_load & _GEN_2081);
  wire        _GEN_2178 = commit_store | ~(commit_load & _GEN_2082);
  wire        _GEN_2179 = commit_store | ~(commit_load & _GEN_2083);
  wire        _GEN_2180 = commit_store | ~(commit_load & _GEN_2084);
  wire        _GEN_2181 = commit_store | ~(commit_load & _GEN_2085);
  wire        _GEN_2182 = commit_store | ~(commit_load & _GEN_2086);
  wire        _GEN_2183 = commit_store | ~(commit_load & _GEN_2087);
  wire        _GEN_2184 = commit_store | ~(commit_load & _GEN_2088);
  wire        _GEN_2185 = commit_store | ~(commit_load & _GEN_2089);
  wire        _GEN_2186 = commit_store | ~(commit_load & _GEN_2090);
  wire        _GEN_2187 = commit_store | ~(commit_load & _GEN_2091);
  wire        _GEN_2188 = commit_store | ~(commit_load & (&idx));
  wire        _GEN_2189 = idx_1 == 5'h0;
  wire        _GEN_2190 = idx_1 == 5'h1;
  wire        _GEN_2191 = idx_1 == 5'h2;
  wire        _GEN_2192 = idx_1 == 5'h3;
  wire        _GEN_2193 = idx_1 == 5'h4;
  wire        _GEN_2194 = idx_1 == 5'h5;
  wire        _GEN_2195 = idx_1 == 5'h6;
  wire        _GEN_2196 = idx_1 == 5'h7;
  wire        _GEN_2197 = idx_1 == 5'h8;
  wire        _GEN_2198 = idx_1 == 5'h9;
  wire        _GEN_2199 = idx_1 == 5'hA;
  wire        _GEN_2200 = idx_1 == 5'hB;
  wire        _GEN_2201 = idx_1 == 5'hC;
  wire        _GEN_2202 = idx_1 == 5'hD;
  wire        _GEN_2203 = idx_1 == 5'hE;
  wire        _GEN_2204 = idx_1 == 5'hF;
  wire        _GEN_2205 = idx_1 == 5'h10;
  wire        _GEN_2206 = idx_1 == 5'h11;
  wire        _GEN_2207 = idx_1 == 5'h12;
  wire        _GEN_2208 = idx_1 == 5'h13;
  wire        _GEN_2209 = idx_1 == 5'h14;
  wire        _GEN_2210 = idx_1 == 5'h15;
  wire        _GEN_2211 = idx_1 == 5'h16;
  wire        _GEN_2212 = idx_1 == 5'h17;
  wire        _GEN_2213 = idx_1 == 5'h18;
  wire        _GEN_2214 = idx_1 == 5'h19;
  wire        _GEN_2215 = idx_1 == 5'h1A;
  wire        _GEN_2216 = idx_1 == 5'h1B;
  wire        _GEN_2217 = idx_1 == 5'h1C;
  wire        _GEN_2218 = idx_1 == 5'h1D;
  wire        _GEN_2219 = idx_1 == 5'h1E;
  wire        _GEN_137950 = commit_store_1 ? _GEN_2189 | _GEN_2124 | _GEN_55040 : _GEN_2124 | _GEN_55040;
  wire        _GEN_137951 = commit_store_1 ? _GEN_2190 | _GEN_2125 | _GEN_55041 : _GEN_2125 | _GEN_55041;
  wire        _GEN_137952 = commit_store_1 ? _GEN_2191 | _GEN_2126 | _GEN_55042 : _GEN_2126 | _GEN_55042;
  wire        _GEN_137953 = commit_store_1 ? _GEN_2192 | _GEN_2127 | _GEN_55043 : _GEN_2127 | _GEN_55043;
  wire        _GEN_137954 = commit_store_1 ? _GEN_2193 | _GEN_2128 | _GEN_55044 : _GEN_2128 | _GEN_55044;
  wire        _GEN_137955 = commit_store_1 ? _GEN_2194 | _GEN_2129 | _GEN_55045 : _GEN_2129 | _GEN_55045;
  wire        _GEN_137956 = commit_store_1 ? _GEN_2195 | _GEN_2130 | _GEN_55046 : _GEN_2130 | _GEN_55046;
  wire        _GEN_137957 = commit_store_1 ? _GEN_2196 | _GEN_2131 | _GEN_55047 : _GEN_2131 | _GEN_55047;
  wire        _GEN_137958 = commit_store_1 ? _GEN_2197 | _GEN_2132 | _GEN_55048 : _GEN_2132 | _GEN_55048;
  wire        _GEN_137959 = commit_store_1 ? _GEN_2198 | _GEN_2133 | _GEN_55049 : _GEN_2133 | _GEN_55049;
  wire        _GEN_137960 = commit_store_1 ? _GEN_2199 | _GEN_2134 | _GEN_55050 : _GEN_2134 | _GEN_55050;
  wire        _GEN_137961 = commit_store_1 ? _GEN_2200 | _GEN_2135 | _GEN_55051 : _GEN_2135 | _GEN_55051;
  wire        _GEN_137962 = commit_store_1 ? _GEN_2201 | _GEN_2136 | _GEN_55052 : _GEN_2136 | _GEN_55052;
  wire        _GEN_137963 = commit_store_1 ? _GEN_2202 | _GEN_2137 | _GEN_55053 : _GEN_2137 | _GEN_55053;
  wire        _GEN_137964 = commit_store_1 ? _GEN_2203 | _GEN_2138 | _GEN_55054 : _GEN_2138 | _GEN_55054;
  wire        _GEN_137965 = commit_store_1 ? _GEN_2204 | _GEN_2139 | _GEN_55055 : _GEN_2139 | _GEN_55055;
  wire        _GEN_137966 = commit_store_1 ? _GEN_2205 | _GEN_2140 | _GEN_55056 : _GEN_2140 | _GEN_55056;
  wire        _GEN_137967 = commit_store_1 ? _GEN_2206 | _GEN_2141 | _GEN_55057 : _GEN_2141 | _GEN_55057;
  wire        _GEN_137968 = commit_store_1 ? _GEN_2207 | _GEN_2142 | _GEN_55058 : _GEN_2142 | _GEN_55058;
  wire        _GEN_137969 = commit_store_1 ? _GEN_2208 | _GEN_2143 | _GEN_55059 : _GEN_2143 | _GEN_55059;
  wire        _GEN_137970 = commit_store_1 ? _GEN_2209 | _GEN_2144 | _GEN_55060 : _GEN_2144 | _GEN_55060;
  wire        _GEN_137971 = commit_store_1 ? _GEN_2210 | _GEN_2145 | _GEN_55061 : _GEN_2145 | _GEN_55061;
  wire        _GEN_137972 = commit_store_1 ? _GEN_2211 | _GEN_2146 | _GEN_55062 : _GEN_2146 | _GEN_55062;
  wire        _GEN_137973 = commit_store_1 ? _GEN_2212 | _GEN_2147 | _GEN_55063 : _GEN_2147 | _GEN_55063;
  wire        _GEN_137974 = commit_store_1 ? _GEN_2213 | _GEN_2148 | _GEN_55064 : _GEN_2148 | _GEN_55064;
  wire        _GEN_137975 = commit_store_1 ? _GEN_2214 | _GEN_2149 | _GEN_55065 : _GEN_2149 | _GEN_55065;
  wire        _GEN_137976 = commit_store_1 ? _GEN_2215 | _GEN_2150 | _GEN_55066 : _GEN_2150 | _GEN_55066;
  wire        _GEN_137977 = commit_store_1 ? _GEN_2216 | _GEN_2151 | _GEN_55067 : _GEN_2151 | _GEN_55067;
  wire        _GEN_137978 = commit_store_1 ? _GEN_2217 | _GEN_2152 | _GEN_55068 : _GEN_2152 | _GEN_55068;
  wire        _GEN_137979 = commit_store_1 ? _GEN_2218 | _GEN_2153 | _GEN_55069 : _GEN_2153 | _GEN_55069;
  wire        _GEN_137980 = commit_store_1 ? _GEN_2219 | _GEN_2154 | _GEN_55070 : _GEN_2154 | _GEN_55070;
  wire        _GEN_137981 = commit_store_1 ? (&idx_1) | _GEN_2155 | _GEN_55071 : _GEN_2155 | _GEN_55071;
  wire        _GEN_2220 = commit_store_1 | ~(commit_load_1 & _GEN_2189);
  wire        _GEN_2221 = commit_store_1 | ~(commit_load_1 & _GEN_2190);
  wire        _GEN_2222 = commit_store_1 | ~(commit_load_1 & _GEN_2191);
  wire        _GEN_2223 = commit_store_1 | ~(commit_load_1 & _GEN_2192);
  wire        _GEN_2224 = commit_store_1 | ~(commit_load_1 & _GEN_2193);
  wire        _GEN_2225 = commit_store_1 | ~(commit_load_1 & _GEN_2194);
  wire        _GEN_2226 = commit_store_1 | ~(commit_load_1 & _GEN_2195);
  wire        _GEN_2227 = commit_store_1 | ~(commit_load_1 & _GEN_2196);
  wire        _GEN_2228 = commit_store_1 | ~(commit_load_1 & _GEN_2197);
  wire        _GEN_2229 = commit_store_1 | ~(commit_load_1 & _GEN_2198);
  wire        _GEN_2230 = commit_store_1 | ~(commit_load_1 & _GEN_2199);
  wire        _GEN_2231 = commit_store_1 | ~(commit_load_1 & _GEN_2200);
  wire        _GEN_2232 = commit_store_1 | ~(commit_load_1 & _GEN_2201);
  wire        _GEN_2233 = commit_store_1 | ~(commit_load_1 & _GEN_2202);
  wire        _GEN_2234 = commit_store_1 | ~(commit_load_1 & _GEN_2203);
  wire        _GEN_2235 = commit_store_1 | ~(commit_load_1 & _GEN_2204);
  wire        _GEN_2236 = commit_store_1 | ~(commit_load_1 & _GEN_2205);
  wire        _GEN_2237 = commit_store_1 | ~(commit_load_1 & _GEN_2206);
  wire        _GEN_2238 = commit_store_1 | ~(commit_load_1 & _GEN_2207);
  wire        _GEN_2239 = commit_store_1 | ~(commit_load_1 & _GEN_2208);
  wire        _GEN_2240 = commit_store_1 | ~(commit_load_1 & _GEN_2209);
  wire        _GEN_2241 = commit_store_1 | ~(commit_load_1 & _GEN_2210);
  wire        _GEN_2242 = commit_store_1 | ~(commit_load_1 & _GEN_2211);
  wire        _GEN_2243 = commit_store_1 | ~(commit_load_1 & _GEN_2212);
  wire        _GEN_2244 = commit_store_1 | ~(commit_load_1 & _GEN_2213);
  wire        _GEN_2245 = commit_store_1 | ~(commit_load_1 & _GEN_2214);
  wire        _GEN_2246 = commit_store_1 | ~(commit_load_1 & _GEN_2215);
  wire        _GEN_2247 = commit_store_1 | ~(commit_load_1 & _GEN_2216);
  wire        _GEN_2248 = commit_store_1 | ~(commit_load_1 & _GEN_2217);
  wire        _GEN_2249 = commit_store_1 | ~(commit_load_1 & _GEN_2218);
  wire        _GEN_2250 = commit_store_1 | ~(commit_load_1 & _GEN_2219);
  wire        _GEN_2251 = commit_store_1 | ~(commit_load_1 & (&idx_1));
  wire        _GEN_2252 = idx_2 == 5'h0;
  wire        _GEN_2253 = idx_2 == 5'h1;
  wire        _GEN_2254 = idx_2 == 5'h2;
  wire        _GEN_2255 = idx_2 == 5'h3;
  wire        _GEN_2256 = idx_2 == 5'h4;
  wire        _GEN_2257 = idx_2 == 5'h5;
  wire        _GEN_2258 = idx_2 == 5'h6;
  wire        _GEN_2259 = idx_2 == 5'h7;
  wire        _GEN_2260 = idx_2 == 5'h8;
  wire        _GEN_2261 = idx_2 == 5'h9;
  wire        _GEN_2262 = idx_2 == 5'hA;
  wire        _GEN_2263 = idx_2 == 5'hB;
  wire        _GEN_2264 = idx_2 == 5'hC;
  wire        _GEN_2265 = idx_2 == 5'hD;
  wire        _GEN_2266 = idx_2 == 5'hE;
  wire        _GEN_2267 = idx_2 == 5'hF;
  wire        _GEN_2268 = idx_2 == 5'h10;
  wire        _GEN_2269 = idx_2 == 5'h11;
  wire        _GEN_2270 = idx_2 == 5'h12;
  wire        _GEN_2271 = idx_2 == 5'h13;
  wire        _GEN_2272 = idx_2 == 5'h14;
  wire        _GEN_2273 = idx_2 == 5'h15;
  wire        _GEN_2274 = idx_2 == 5'h16;
  wire        _GEN_2275 = idx_2 == 5'h17;
  wire        _GEN_2276 = idx_2 == 5'h18;
  wire        _GEN_2277 = idx_2 == 5'h19;
  wire        _GEN_2278 = idx_2 == 5'h1A;
  wire        _GEN_2279 = idx_2 == 5'h1B;
  wire        _GEN_2280 = idx_2 == 5'h1C;
  wire        _GEN_2281 = idx_2 == 5'h1D;
  wire        _GEN_2282 = idx_2 == 5'h1E;
  wire        _GEN_2283 = commit_store_2 & _GEN_2252;
  wire        _GEN_2284 = commit_store_2 & _GEN_2253;
  wire        _GEN_2285 = commit_store_2 & _GEN_2254;
  wire        _GEN_2286 = commit_store_2 & _GEN_2255;
  wire        _GEN_2287 = commit_store_2 & _GEN_2256;
  wire        _GEN_2288 = commit_store_2 & _GEN_2257;
  wire        _GEN_2289 = commit_store_2 & _GEN_2258;
  wire        _GEN_2290 = commit_store_2 & _GEN_2259;
  wire        _GEN_2291 = commit_store_2 & _GEN_2260;
  wire        _GEN_2292 = commit_store_2 & _GEN_2261;
  wire        _GEN_2293 = commit_store_2 & _GEN_2262;
  wire        _GEN_2294 = commit_store_2 & _GEN_2263;
  wire        _GEN_2295 = commit_store_2 & _GEN_2264;
  wire        _GEN_2296 = commit_store_2 & _GEN_2265;
  wire        _GEN_2297 = commit_store_2 & _GEN_2266;
  wire        _GEN_2298 = commit_store_2 & _GEN_2267;
  wire        _GEN_2299 = commit_store_2 & _GEN_2268;
  wire        _GEN_2300 = commit_store_2 & _GEN_2269;
  wire        _GEN_2301 = commit_store_2 & _GEN_2270;
  wire        _GEN_2302 = commit_store_2 & _GEN_2271;
  wire        _GEN_2303 = commit_store_2 & _GEN_2272;
  wire        _GEN_2304 = commit_store_2 & _GEN_2273;
  wire        _GEN_2305 = commit_store_2 & _GEN_2274;
  wire        _GEN_2306 = commit_store_2 & _GEN_2275;
  wire        _GEN_2307 = commit_store_2 & _GEN_2276;
  wire        _GEN_2308 = commit_store_2 & _GEN_2277;
  wire        _GEN_2309 = commit_store_2 & _GEN_2278;
  wire        _GEN_2310 = commit_store_2 & _GEN_2279;
  wire        _GEN_2311 = commit_store_2 & _GEN_2280;
  wire        _GEN_2312 = commit_store_2 & _GEN_2281;
  wire        _GEN_2313 = commit_store_2 & _GEN_2282;
  wire        _GEN_2314 = commit_store_2 & (&idx_2);
  wire        _GEN_2315 = commit_store_2 | ~(commit_load_2 & _GEN_2252);
  wire        _GEN_2316 = commit_store_2 | ~(commit_load_2 & _GEN_2253);
  wire        _GEN_2317 = commit_store_2 | ~(commit_load_2 & _GEN_2254);
  wire        _GEN_2318 = commit_store_2 | ~(commit_load_2 & _GEN_2255);
  wire        _GEN_2319 = commit_store_2 | ~(commit_load_2 & _GEN_2256);
  wire        _GEN_2320 = commit_store_2 | ~(commit_load_2 & _GEN_2257);
  wire        _GEN_2321 = commit_store_2 | ~(commit_load_2 & _GEN_2258);
  wire        _GEN_2322 = commit_store_2 | ~(commit_load_2 & _GEN_2259);
  wire        _GEN_2323 = commit_store_2 | ~(commit_load_2 & _GEN_2260);
  wire        _GEN_2324 = commit_store_2 | ~(commit_load_2 & _GEN_2261);
  wire        _GEN_2325 = commit_store_2 | ~(commit_load_2 & _GEN_2262);
  wire        _GEN_2326 = commit_store_2 | ~(commit_load_2 & _GEN_2263);
  wire        _GEN_2327 = commit_store_2 | ~(commit_load_2 & _GEN_2264);
  wire        _GEN_2328 = commit_store_2 | ~(commit_load_2 & _GEN_2265);
  wire        _GEN_2329 = commit_store_2 | ~(commit_load_2 & _GEN_2266);
  wire        _GEN_2330 = commit_store_2 | ~(commit_load_2 & _GEN_2267);
  wire        _GEN_2331 = commit_store_2 | ~(commit_load_2 & _GEN_2268);
  wire        _GEN_2332 = commit_store_2 | ~(commit_load_2 & _GEN_2269);
  wire        _GEN_2333 = commit_store_2 | ~(commit_load_2 & _GEN_2270);
  wire        _GEN_2334 = commit_store_2 | ~(commit_load_2 & _GEN_2271);
  wire        _GEN_2335 = commit_store_2 | ~(commit_load_2 & _GEN_2272);
  wire        _GEN_2336 = commit_store_2 | ~(commit_load_2 & _GEN_2273);
  wire        _GEN_2337 = commit_store_2 | ~(commit_load_2 & _GEN_2274);
  wire        _GEN_2338 = commit_store_2 | ~(commit_load_2 & _GEN_2275);
  wire        _GEN_2339 = commit_store_2 | ~(commit_load_2 & _GEN_2276);
  wire        _GEN_2340 = commit_store_2 | ~(commit_load_2 & _GEN_2277);
  wire        _GEN_2341 = commit_store_2 | ~(commit_load_2 & _GEN_2278);
  wire        _GEN_2342 = commit_store_2 | ~(commit_load_2 & _GEN_2279);
  wire        _GEN_2343 = commit_store_2 | ~(commit_load_2 & _GEN_2280);
  wire        _GEN_2344 = commit_store_2 | ~(commit_load_2 & _GEN_2281);
  wire        _GEN_2345 = commit_store_2 | ~(commit_load_2 & _GEN_2282);
  wire        _GEN_2346 = commit_store_2 | ~(commit_load_2 & (&idx_2));
  wire        _GEN_2347 = idx_3 == 5'h0;
  wire        _GEN_2348 = idx_3 == 5'h1;
  wire        _GEN_2349 = idx_3 == 5'h2;
  wire        _GEN_2350 = idx_3 == 5'h3;
  wire        _GEN_2351 = idx_3 == 5'h4;
  wire        _GEN_2352 = idx_3 == 5'h5;
  wire        _GEN_2353 = idx_3 == 5'h6;
  wire        _GEN_2354 = idx_3 == 5'h7;
  wire        _GEN_2355 = idx_3 == 5'h8;
  wire        _GEN_2356 = idx_3 == 5'h9;
  wire        _GEN_2357 = idx_3 == 5'hA;
  wire        _GEN_2358 = idx_3 == 5'hB;
  wire        _GEN_2359 = idx_3 == 5'hC;
  wire        _GEN_2360 = idx_3 == 5'hD;
  wire        _GEN_2361 = idx_3 == 5'hE;
  wire        _GEN_2362 = idx_3 == 5'hF;
  wire        _GEN_2363 = idx_3 == 5'h10;
  wire        _GEN_2364 = idx_3 == 5'h11;
  wire        _GEN_2365 = idx_3 == 5'h12;
  wire        _GEN_2366 = idx_3 == 5'h13;
  wire        _GEN_2367 = idx_3 == 5'h14;
  wire        _GEN_2368 = idx_3 == 5'h15;
  wire        _GEN_2369 = idx_3 == 5'h16;
  wire        _GEN_2370 = idx_3 == 5'h17;
  wire        _GEN_2371 = idx_3 == 5'h18;
  wire        _GEN_2372 = idx_3 == 5'h19;
  wire        _GEN_2373 = idx_3 == 5'h1A;
  wire        _GEN_2374 = idx_3 == 5'h1B;
  wire        _GEN_2375 = idx_3 == 5'h1C;
  wire        _GEN_2376 = idx_3 == 5'h1D;
  wire        _GEN_2377 = idx_3 == 5'h1E;
  wire        _GEN_2378 = commit_store_3 | ~(commit_load_3 & _GEN_2347);
  wire        _GEN_2379 = commit_store_3 | ~(commit_load_3 & _GEN_2348);
  wire        _GEN_2380 = commit_store_3 | ~(commit_load_3 & _GEN_2349);
  wire        _GEN_2381 = commit_store_3 | ~(commit_load_3 & _GEN_2350);
  wire        _GEN_2382 = commit_store_3 | ~(commit_load_3 & _GEN_2351);
  wire        _GEN_2383 = commit_store_3 | ~(commit_load_3 & _GEN_2352);
  wire        _GEN_2384 = commit_store_3 | ~(commit_load_3 & _GEN_2353);
  wire        _GEN_2385 = commit_store_3 | ~(commit_load_3 & _GEN_2354);
  wire        _GEN_2386 = commit_store_3 | ~(commit_load_3 & _GEN_2355);
  wire        _GEN_2387 = commit_store_3 | ~(commit_load_3 & _GEN_2356);
  wire        _GEN_2388 = commit_store_3 | ~(commit_load_3 & _GEN_2357);
  wire        _GEN_2389 = commit_store_3 | ~(commit_load_3 & _GEN_2358);
  wire        _GEN_2390 = commit_store_3 | ~(commit_load_3 & _GEN_2359);
  wire        _GEN_2391 = commit_store_3 | ~(commit_load_3 & _GEN_2360);
  wire        _GEN_2392 = commit_store_3 | ~(commit_load_3 & _GEN_2361);
  wire        _GEN_2393 = commit_store_3 | ~(commit_load_3 & _GEN_2362);
  wire        _GEN_2394 = commit_store_3 | ~(commit_load_3 & _GEN_2363);
  wire        _GEN_2395 = commit_store_3 | ~(commit_load_3 & _GEN_2364);
  wire        _GEN_2396 = commit_store_3 | ~(commit_load_3 & _GEN_2365);
  wire        _GEN_2397 = commit_store_3 | ~(commit_load_3 & _GEN_2366);
  wire        _GEN_2398 = commit_store_3 | ~(commit_load_3 & _GEN_2367);
  wire        _GEN_2399 = commit_store_3 | ~(commit_load_3 & _GEN_2368);
  wire        _GEN_2400 = commit_store_3 | ~(commit_load_3 & _GEN_2369);
  wire        _GEN_2401 = commit_store_3 | ~(commit_load_3 & _GEN_2370);
  wire        _GEN_2402 = commit_store_3 | ~(commit_load_3 & _GEN_2371);
  wire        _GEN_2403 = commit_store_3 | ~(commit_load_3 & _GEN_2372);
  wire        _GEN_2404 = commit_store_3 | ~(commit_load_3 & _GEN_2373);
  wire        _GEN_2405 = commit_store_3 | ~(commit_load_3 & _GEN_2374);
  wire        _GEN_2406 = commit_store_3 | ~(commit_load_3 & _GEN_2375);
  wire        _GEN_2407 = commit_store_3 | ~(commit_load_3 & _GEN_2376);
  wire        _GEN_2408 = commit_store_3 | ~(commit_load_3 & _GEN_2377);
  wire        _GEN_2409 = commit_store_3 | ~(commit_load_3 & (&idx_3));
  wire        _GEN_2410 = stq_head == 5'h0;
  wire        _GEN_2411 = _GEN_2410 | _GEN_1997;
  wire        _GEN_2412 = _GEN_1237 | _GEN_1998;
  wire        _GEN_2413 = _GEN_1238 | _GEN_1999;
  wire        _GEN_2414 = _GEN_1239 | _GEN_2000;
  wire        _GEN_2415 = _GEN_1240 | _GEN_2001;
  wire        _GEN_2416 = _GEN_1241 | _GEN_2002;
  wire        _GEN_2417 = _GEN_1242 | _GEN_2003;
  wire        _GEN_2418 = _GEN_1243 | _GEN_2004;
  wire        _GEN_2419 = _GEN_1244 | _GEN_2005;
  wire        _GEN_2420 = _GEN_1245 | _GEN_2006;
  wire        _GEN_2421 = _GEN_1246 | _GEN_2007;
  wire        _GEN_2422 = _GEN_1247 | _GEN_2008;
  wire        _GEN_2423 = _GEN_1248 | _GEN_2009;
  wire        _GEN_2424 = _GEN_1249 | _GEN_2010;
  wire        _GEN_2425 = _GEN_1250 | _GEN_2011;
  wire        _GEN_2426 = _GEN_1251 | _GEN_2012;
  wire        _GEN_2427 = _GEN_1252 | _GEN_2013;
  wire        _GEN_2428 = _GEN_1253 | _GEN_2014;
  wire        _GEN_2429 = _GEN_1254 | _GEN_2015;
  wire        _GEN_2430 = _GEN_1255 | _GEN_2016;
  wire        _GEN_2431 = _GEN_1256 | _GEN_2017;
  wire        _GEN_2432 = _GEN_1257 | _GEN_2018;
  wire        _GEN_2433 = _GEN_1258 | _GEN_2019;
  wire        _GEN_2434 = _GEN_1259 | _GEN_2020;
  wire        _GEN_2435 = _GEN_1260 | _GEN_2021;
  wire        _GEN_2436 = _GEN_1261 | _GEN_2022;
  wire        _GEN_2437 = _GEN_1262 | _GEN_2023;
  wire        _GEN_2438 = _GEN_1263 | _GEN_2024;
  wire        _GEN_2439 = _GEN_1264 | _GEN_2025;
  wire        _GEN_2440 = _GEN_1265 | _GEN_2026;
  wire        _GEN_2441 = _GEN_1266 | _GEN_2027;
  wire        _GEN_2442 = (&stq_head) | _GEN_2028;
  wire        _GEN_2443 = clear_store & _GEN_2410;
  wire        _GEN_2444 = clear_store & _GEN_1237;
  wire        _GEN_2445 = clear_store & _GEN_1238;
  wire        _GEN_2446 = clear_store & _GEN_1239;
  wire        _GEN_2447 = clear_store & _GEN_1240;
  wire        _GEN_2448 = clear_store & _GEN_1241;
  wire        _GEN_2449 = clear_store & _GEN_1242;
  wire        _GEN_2450 = clear_store & _GEN_1243;
  wire        _GEN_2451 = clear_store & _GEN_1244;
  wire        _GEN_2452 = clear_store & _GEN_1245;
  wire        _GEN_2453 = clear_store & _GEN_1246;
  wire        _GEN_2454 = clear_store & _GEN_1247;
  wire        _GEN_2455 = clear_store & _GEN_1248;
  wire        _GEN_2456 = clear_store & _GEN_1249;
  wire        _GEN_2457 = clear_store & _GEN_1250;
  wire        _GEN_2458 = clear_store & _GEN_1251;
  wire        _GEN_2459 = clear_store & _GEN_1252;
  wire        _GEN_2460 = clear_store & _GEN_1253;
  wire        _GEN_2461 = clear_store & _GEN_1254;
  wire        _GEN_2462 = clear_store & _GEN_1255;
  wire        _GEN_2463 = clear_store & _GEN_1256;
  wire        _GEN_2464 = clear_store & _GEN_1257;
  wire        _GEN_2465 = clear_store & _GEN_1258;
  wire        _GEN_2466 = clear_store & _GEN_1259;
  wire        _GEN_2467 = clear_store & _GEN_1260;
  wire        _GEN_2468 = clear_store & _GEN_1261;
  wire        _GEN_2469 = clear_store & _GEN_1262;
  wire        _GEN_2470 = clear_store & _GEN_1263;
  wire        _GEN_2471 = clear_store & _GEN_1264;
  wire        _GEN_2472 = clear_store & _GEN_1265;
  wire        _GEN_2473 = clear_store & _GEN_1266;
  wire        _GEN_2474 = clear_store & (&stq_head);
  wire        _GEN_2475 = ~(|hella_state) & io_hellacache_req_valid;
  wire        _GEN_2476 = ~(|hella_state) & _GEN_2475;
  wire        _GEN_2477 = (|hella_state) & _GEN_140251;
  wire        _GEN_2478 = ~(|hella_state) | ~_GEN_140251;
  wire        _GEN_140325 = ~stq_0_bits_committed & ~stq_0_bits_succeeded;
  wire        _GEN_140329 = ~stq_1_bits_committed & ~stq_1_bits_succeeded;
  wire        _GEN_140333 = ~stq_2_bits_committed & ~stq_2_bits_succeeded;
  wire        _GEN_140337 = ~stq_3_bits_committed & ~stq_3_bits_succeeded;
  wire        _GEN_140341 = ~stq_4_bits_committed & ~stq_4_bits_succeeded;
  wire        _GEN_140345 = ~stq_5_bits_committed & ~stq_5_bits_succeeded;
  wire        _GEN_140349 = ~stq_6_bits_committed & ~stq_6_bits_succeeded;
  wire        _GEN_140353 = ~stq_7_bits_committed & ~stq_7_bits_succeeded;
  wire        _GEN_140357 = ~stq_8_bits_committed & ~stq_8_bits_succeeded;
  wire        _GEN_140361 = ~stq_9_bits_committed & ~stq_9_bits_succeeded;
  wire        _GEN_140365 = ~stq_10_bits_committed & ~stq_10_bits_succeeded;
  wire        _GEN_140369 = ~stq_11_bits_committed & ~stq_11_bits_succeeded;
  wire        _GEN_140373 = ~stq_12_bits_committed & ~stq_12_bits_succeeded;
  wire        _GEN_140377 = ~stq_13_bits_committed & ~stq_13_bits_succeeded;
  wire        _GEN_140381 = ~stq_14_bits_committed & ~stq_14_bits_succeeded;
  wire        _GEN_140385 = ~stq_15_bits_committed & ~stq_15_bits_succeeded;
  wire        _GEN_140389 = ~stq_16_bits_committed & ~stq_16_bits_succeeded;
  wire        _GEN_140393 = ~stq_17_bits_committed & ~stq_17_bits_succeeded;
  wire        _GEN_140397 = ~stq_18_bits_committed & ~stq_18_bits_succeeded;
  wire        _GEN_140401 = ~stq_19_bits_committed & ~stq_19_bits_succeeded;
  wire        _GEN_140405 = ~stq_20_bits_committed & ~stq_20_bits_succeeded;
  wire        _GEN_140409 = ~stq_21_bits_committed & ~stq_21_bits_succeeded;
  wire        _GEN_140413 = ~stq_22_bits_committed & ~stq_22_bits_succeeded;
  wire        _GEN_140417 = ~stq_23_bits_committed & ~stq_23_bits_succeeded;
  wire        _GEN_140421 = ~stq_24_bits_committed & ~stq_24_bits_succeeded;
  wire        _GEN_140425 = ~stq_25_bits_committed & ~stq_25_bits_succeeded;
  wire        _GEN_140429 = ~stq_26_bits_committed & ~stq_26_bits_succeeded;
  wire        _GEN_140433 = ~stq_27_bits_committed & ~stq_27_bits_succeeded;
  wire        _GEN_140437 = ~stq_28_bits_committed & ~stq_28_bits_succeeded;
  wire        _GEN_140441 = ~stq_29_bits_committed & ~stq_29_bits_succeeded;
  wire        _GEN_140445 = ~stq_30_bits_committed & ~stq_30_bits_succeeded;
  wire        _GEN_140449 = ~stq_31_bits_committed & ~stq_31_bits_succeeded;
  wire        _GEN_2479 = _GEN_1234 & (reset | _GEN_140325);
  wire        _GEN_2480 = _GEN_1234 & (reset | _GEN_140329);
  wire        _GEN_2481 = _GEN_1234 & (reset | _GEN_140333);
  wire        _GEN_2482 = _GEN_1234 & (reset | _GEN_140337);
  wire        _GEN_2483 = _GEN_1234 & (reset | _GEN_140341);
  wire        _GEN_2484 = _GEN_1234 & (reset | _GEN_140345);
  wire        _GEN_2485 = _GEN_1234 & (reset | _GEN_140349);
  wire        _GEN_2486 = _GEN_1234 & (reset | _GEN_140353);
  wire        _GEN_2487 = _GEN_1234 & (reset | _GEN_140357);
  wire        _GEN_2488 = _GEN_1234 & (reset | _GEN_140361);
  wire        _GEN_2489 = _GEN_1234 & (reset | _GEN_140365);
  wire        _GEN_2490 = _GEN_1234 & (reset | _GEN_140369);
  wire        _GEN_2491 = _GEN_1234 & (reset | _GEN_140373);
  wire        _GEN_2492 = _GEN_1234 & (reset | _GEN_140377);
  wire        _GEN_2493 = _GEN_1234 & (reset | _GEN_140381);
  wire        _GEN_2494 = _GEN_1234 & (reset | _GEN_140385);
  wire        _GEN_2495 = _GEN_1234 & (reset | _GEN_140389);
  wire        _GEN_2496 = _GEN_1234 & (reset | _GEN_140393);
  wire        _GEN_2497 = _GEN_1234 & (reset | _GEN_140397);
  wire        _GEN_2498 = _GEN_1234 & (reset | _GEN_140401);
  wire        _GEN_2499 = _GEN_1234 & (reset | _GEN_140405);
  wire        _GEN_2500 = _GEN_1234 & (reset | _GEN_140409);
  wire        _GEN_2501 = _GEN_1234 & (reset | _GEN_140413);
  wire        _GEN_2502 = _GEN_1234 & (reset | _GEN_140417);
  wire        _GEN_2503 = _GEN_1234 & (reset | _GEN_140421);
  wire        _GEN_2504 = _GEN_1234 & (reset | _GEN_140425);
  wire        _GEN_2505 = _GEN_1234 & (reset | _GEN_140429);
  wire        _GEN_2506 = _GEN_1234 & (reset | _GEN_140433);
  wire        _GEN_2507 = _GEN_1234 & (reset | _GEN_140437);
  wire        _GEN_2508 = _GEN_1234 & (reset | _GEN_140441);
  wire        _GEN_2509 = _GEN_1234 & (reset | _GEN_140445);
  wire        _GEN_2510 = _GEN_1234 & (reset | _GEN_140449);
  wire [5:0]  _ldq_wakeup_idx_idx_T_42 = _ldq_wakeup_idx_T_167 & _temp_bits_T_40 ? 6'h14 : _ldq_wakeup_idx_T_175 & _temp_bits_T_42 ? 6'h15 : _ldq_wakeup_idx_T_183 & _temp_bits_T_44 ? 6'h16 : _ldq_wakeup_idx_T_191 & _temp_bits_T_46 ? 6'h17 : _ldq_wakeup_idx_T_199 & _temp_bits_T_48 ? 6'h18 : _ldq_wakeup_idx_T_207 & _temp_bits_T_50 ? 6'h19 : _ldq_wakeup_idx_T_215 & _temp_bits_T_52 ? 6'h1A : _ldq_wakeup_idx_T_223 & _temp_bits_T_54 ? 6'h1B : _ldq_wakeup_idx_T_231 & _temp_bits_T_56 ? 6'h1C : _ldq_wakeup_idx_T_239 & _temp_bits_T_58 ? 6'h1D : _ldq_wakeup_idx_T_247 & _temp_bits_T_60 ? 6'h1E : ldq_31_bits_addr_valid & ~ldq_31_bits_executed & ~ldq_31_bits_succeeded & ~ldq_31_bits_addr_is_virtual & ~ldq_retry_idx_block_31 ? 6'h1F : _ldq_wakeup_idx_T_7 ? 6'h20 : _ldq_wakeup_idx_T_15 ? 6'h21 : _ldq_wakeup_idx_T_23 ? 6'h22 : _ldq_wakeup_idx_T_31 ? 6'h23 : _ldq_wakeup_idx_T_39 ? 6'h24 : _ldq_wakeup_idx_T_47 ? 6'h25 : _ldq_wakeup_idx_T_55 ? 6'h26 : _ldq_wakeup_idx_T_63 ? 6'h27 : _ldq_wakeup_idx_T_71 ? 6'h28 : _ldq_wakeup_idx_T_79 ? 6'h29 : _ldq_wakeup_idx_T_87 ? 6'h2A : _ldq_wakeup_idx_T_95 ? 6'h2B : _ldq_wakeup_idx_T_103 ? 6'h2C : _ldq_wakeup_idx_T_111 ? 6'h2D : _ldq_wakeup_idx_T_119 ? 6'h2E : _ldq_wakeup_idx_T_127 ? 6'h2F : _ldq_wakeup_idx_T_135 ? 6'h30 : _ldq_wakeup_idx_T_143 ? 6'h31 : _ldq_wakeup_idx_T_151 ? 6'h32 : _ldq_wakeup_idx_T_159 ? 6'h33 : _ldq_wakeup_idx_T_167 ? 6'h34 : _ldq_wakeup_idx_T_175 ? 6'h35 : _ldq_wakeup_idx_T_183 ? 6'h36 : _ldq_wakeup_idx_T_191 ? 6'h37 : _ldq_wakeup_idx_T_199 ? 6'h38 : _ldq_wakeup_idx_T_207 ? 6'h39 : _ldq_wakeup_idx_T_215 ? 6'h3A : _ldq_wakeup_idx_T_223 ? 6'h3B : _ldq_wakeup_idx_T_231 ? 6'h3C : _ldq_wakeup_idx_T_239 ? 6'h3D : {5'h1F, ~_ldq_wakeup_idx_T_247};
  wire [5:0]  _ldq_retry_idx_idx_T_42 = _ldq_retry_idx_T_62 & _temp_bits_T_40 ? 6'h14 : _ldq_retry_idx_T_65 & _temp_bits_T_42 ? 6'h15 : _ldq_retry_idx_T_68 & _temp_bits_T_44 ? 6'h16 : _ldq_retry_idx_T_71 & _temp_bits_T_46 ? 6'h17 : _ldq_retry_idx_T_74 & _temp_bits_T_48 ? 6'h18 : _ldq_retry_idx_T_77 & _temp_bits_T_50 ? 6'h19 : _ldq_retry_idx_T_80 & _temp_bits_T_52 ? 6'h1A : _ldq_retry_idx_T_83 & _temp_bits_T_54 ? 6'h1B : _ldq_retry_idx_T_86 & _temp_bits_T_56 ? 6'h1C : _ldq_retry_idx_T_89 & _temp_bits_T_58 ? 6'h1D : _ldq_retry_idx_T_92 & _temp_bits_T_60 ? 6'h1E : ldq_31_bits_addr_valid & ldq_31_bits_addr_is_virtual & ~ldq_retry_idx_block_31 ? 6'h1F : _ldq_retry_idx_T_2 ? 6'h20 : _ldq_retry_idx_T_5 ? 6'h21 : _ldq_retry_idx_T_8 ? 6'h22 : _ldq_retry_idx_T_11 ? 6'h23 : _ldq_retry_idx_T_14 ? 6'h24 : _ldq_retry_idx_T_17 ? 6'h25 : _ldq_retry_idx_T_20 ? 6'h26 : _ldq_retry_idx_T_23 ? 6'h27 : _ldq_retry_idx_T_26 ? 6'h28 : _ldq_retry_idx_T_29 ? 6'h29 : _ldq_retry_idx_T_32 ? 6'h2A : _ldq_retry_idx_T_35 ? 6'h2B : _ldq_retry_idx_T_38 ? 6'h2C : _ldq_retry_idx_T_41 ? 6'h2D : _ldq_retry_idx_T_44 ? 6'h2E : _ldq_retry_idx_T_47 ? 6'h2F : _ldq_retry_idx_T_50 ? 6'h30 : _ldq_retry_idx_T_53 ? 6'h31 : _ldq_retry_idx_T_56 ? 6'h32 : _ldq_retry_idx_T_59 ? 6'h33 : _ldq_retry_idx_T_62 ? 6'h34 : _ldq_retry_idx_T_65 ? 6'h35 : _ldq_retry_idx_T_68 ? 6'h36 : _ldq_retry_idx_T_71 ? 6'h37 : _ldq_retry_idx_T_74 ? 6'h38 : _ldq_retry_idx_T_77 ? 6'h39 : _ldq_retry_idx_T_80 ? 6'h3A : _ldq_retry_idx_T_83 ? 6'h3B : _ldq_retry_idx_T_86 ? 6'h3C : _ldq_retry_idx_T_89 ? 6'h3D : {5'h1F, ~_ldq_retry_idx_T_92};
  wire [5:0]  _stq_retry_idx_idx_T_42 = _stq_retry_idx_T_20 & stq_commit_head < 5'h15 ? 6'h14 : _stq_retry_idx_T_21 & stq_commit_head < 5'h16 ? 6'h15 : _stq_retry_idx_T_22 & stq_commit_head < 5'h17 ? 6'h16 : _stq_retry_idx_T_23 & stq_commit_head[4:3] != 2'h3 ? 6'h17 : _stq_retry_idx_T_24 & stq_commit_head < 5'h19 ? 6'h18 : _stq_retry_idx_T_25 & stq_commit_head < 5'h1A ? 6'h19 : _stq_retry_idx_T_26 & stq_commit_head < 5'h1B ? 6'h1A : _stq_retry_idx_T_27 & stq_commit_head[4:2] != 3'h7 ? 6'h1B : _stq_retry_idx_T_28 & stq_commit_head < 5'h1D ? 6'h1C : _stq_retry_idx_T_29 & stq_commit_head[4:1] != 4'hF ? 6'h1D : _stq_retry_idx_T_30 & stq_commit_head != 5'h1F ? 6'h1E : stq_31_bits_addr_valid & stq_31_bits_addr_is_virtual ? 6'h1F : _stq_retry_idx_T ? 6'h20 : _stq_retry_idx_T_1 ? 6'h21 : _stq_retry_idx_T_2 ? 6'h22 : _stq_retry_idx_T_3 ? 6'h23 : _stq_retry_idx_T_4 ? 6'h24 : _stq_retry_idx_T_5 ? 6'h25 : _stq_retry_idx_T_6 ? 6'h26 : _stq_retry_idx_T_7 ? 6'h27 : _stq_retry_idx_T_8 ? 6'h28 : _stq_retry_idx_T_9 ? 6'h29 : _stq_retry_idx_T_10 ? 6'h2A : _stq_retry_idx_T_11 ? 6'h2B : _stq_retry_idx_T_12 ? 6'h2C : _stq_retry_idx_T_13 ? 6'h2D : _stq_retry_idx_T_14 ? 6'h2E : _stq_retry_idx_T_15 ? 6'h2F : _stq_retry_idx_T_16 ? 6'h30 : _stq_retry_idx_T_17 ? 6'h31 : _stq_retry_idx_T_18 ? 6'h32 : _stq_retry_idx_T_19 ? 6'h33 : _stq_retry_idx_T_20 ? 6'h34 : _stq_retry_idx_T_21 ? 6'h35 : _stq_retry_idx_T_22 ? 6'h36 : _stq_retry_idx_T_23 ? 6'h37 : _stq_retry_idx_T_24 ? 6'h38 : _stq_retry_idx_T_25 ? 6'h39 : _stq_retry_idx_T_26 ? 6'h3A : _stq_retry_idx_T_27 ? 6'h3B : _stq_retry_idx_T_28 ? 6'h3C : _stq_retry_idx_T_29 ? 6'h3D : {5'h1F, ~_stq_retry_idx_T_30};
  always @(posedge clock) begin
    ldq_0_valid <= ~_GEN_1234 & _GEN_2378 & _GEN_2315 & _GEN_2220 & (_GEN_2156 ? ~_GEN_2029 & _GEN_49600 : ~_GEN_2092 & _GEN_49600);
    if (_GEN_297) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_0_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_0_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_0_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_0_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_0_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_199) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_0_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_0_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_0_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_0_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_132) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_0_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_0_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_0_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_34) begin
      ldq_0_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_0_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_0_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_0_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_0_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_0_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_0_bits_st_dep_mask <= next_live_store_mask;
      ldq_0_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_0_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_0_bits_st_dep_mask;
    if (ldq_0_valid)
      ldq_0_bits_uop_br_mask <= ldq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_297)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_199)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_132)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_34)
      ldq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1649) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_0_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_0_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_0_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_0_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_0_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_0_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_0_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_0_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_0_bits_addr_bits <= hella_req_addr;
        else
          ldq_0_bits_addr_bits <= 40'h0;
      end
      else
        ldq_0_bits_addr_bits <= _GEN_338;
      ldq_0_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_0_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1553) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_0_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_0_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_0_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_0_bits_addr_bits <= _GEN_332;
        else
          ldq_0_bits_addr_bits <= 40'h0;
      end
      else
        ldq_0_bits_addr_bits <= _GEN_334;
      ldq_0_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_0_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_297)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_199)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_132)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_34)
      ldq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_0_bits_addr_valid <= ~_GEN_1234 & _GEN_2378 & _GEN_2315 & _GEN_2220 & (_GEN_2156 ? ~_GEN_2029 & _GEN_81718 : ~_GEN_2092 & _GEN_81718);
    ldq_0_bits_executed <= ~_GEN_1234 & _GEN_2378 & _GEN_2315 & _GEN_2220 & _GEN_2157 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_354) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116695)) & ((_GEN_1174 ? (_GEN_113938 ? (|lcam_ldq_idx_1) & _GEN_113741 : _GEN_1176 ? (|lcam_ldq_idx_1) & _GEN_113741 : ~(_GEN_113869 & ~(|lcam_ldq_idx_1)) & _GEN_113741) : _GEN_113741) | (dis_ld_val_3 ? ~_GEN_1396 & _GEN_24736 : ~_GEN_199 & _GEN_24736));
    ldq_0_bits_succeeded <= _GEN_2378 & _GEN_2315 & _GEN_2220 & _GEN_2157 & (_GEN_1965 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h0 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1900 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h0 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1396 & _GEN_24768 : ~_GEN_199 & _GEN_24768) : casez_tmp_203) : casez_tmp_236);
    ldq_0_bits_order_fail <= _GEN_2378 & _GEN_2315 & _GEN_2220 & _GEN_2157 & (_GEN_357 ? _GEN_83271 : _GEN_360 ? _GEN_361 | _GEN_83271 : _GEN_365 | _GEN_83271);
    ldq_0_bits_observed <= _GEN_357 | (dis_ld_val_3 ? ~_GEN_1396 & _GEN_24832 : ~_GEN_199 & _GEN_24832);
    ldq_0_bits_forward_std_val <= _GEN_2378 & _GEN_2315 & _GEN_2220 & _GEN_2157 & (~_GEN_1183 & _GEN_1933 | ~_GEN_1179 & _GEN_1868 | (dis_ld_val_3 ? ~_GEN_1396 & _GEN_24864 : ~_GEN_199 & _GEN_24864));
    if (_GEN_1965) begin
      if (_GEN_1900) begin
      end
      else
        ldq_0_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_0_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_1_valid <= ~_GEN_1234 & _GEN_2379 & _GEN_2316 & _GEN_2221 & (_GEN_2156 ? ~_GEN_2030 & _GEN_49601 : ~_GEN_2093 & _GEN_49601);
    if (_GEN_298) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_1_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_1_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_1_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_1_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_1_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_200) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_1_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_1_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_1_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_1_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_133) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_1_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_1_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_1_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_35) begin
      ldq_1_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_1_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_1_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_1_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_1_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_1_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_1_bits_st_dep_mask <= next_live_store_mask;
      ldq_1_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_1_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_1_bits_st_dep_mask;
    if (ldq_1_valid)
      ldq_1_bits_uop_br_mask <= ldq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_298)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_200)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_133)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_35)
      ldq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1650) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_1_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_1_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_1_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_1_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_1_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_1_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_1_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_1_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_1_bits_addr_bits <= hella_req_addr;
        else
          ldq_1_bits_addr_bits <= 40'h0;
      end
      else
        ldq_1_bits_addr_bits <= _GEN_338;
      ldq_1_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_1_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1554) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_1_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_1_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_1_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_1_bits_addr_bits <= _GEN_332;
        else
          ldq_1_bits_addr_bits <= 40'h0;
      end
      else
        ldq_1_bits_addr_bits <= _GEN_334;
      ldq_1_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_1_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_298)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_200)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_133)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_35)
      ldq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_1_bits_addr_valid <= ~_GEN_1234 & _GEN_2379 & _GEN_2316 & _GEN_2221 & (_GEN_2156 ? ~_GEN_2030 & _GEN_81719 : ~_GEN_2093 & _GEN_81719);
    ldq_1_bits_executed <= ~_GEN_1234 & _GEN_2379 & _GEN_2316 & _GEN_2221 & _GEN_2158 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_374) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116696)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1773 & _GEN_113742 : _GEN_1176 ? ~_GEN_1773 & _GEN_113742 : ~(_GEN_113869 & _GEN_1773) & _GEN_113742) : _GEN_113742) | (dis_ld_val_3 ? ~_GEN_1397 & _GEN_24737 : ~_GEN_200 & _GEN_24737));
    ldq_1_bits_succeeded <= _GEN_2379 & _GEN_2316 & _GEN_2221 & _GEN_2158 & (_GEN_1966 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1901 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1397 & _GEN_24769 : ~_GEN_200 & _GEN_24769) : casez_tmp_203) : casez_tmp_236);
    ldq_1_bits_order_fail <= _GEN_2379 & _GEN_2316 & _GEN_2221 & _GEN_2158 & (_GEN_377 ? _GEN_83769 : _GEN_379 ? _GEN_380 | _GEN_83769 : _GEN_384 | _GEN_83769);
    ldq_1_bits_observed <= _GEN_377 | (dis_ld_val_3 ? ~_GEN_1397 & _GEN_24833 : ~_GEN_200 & _GEN_24833);
    ldq_1_bits_forward_std_val <= _GEN_2379 & _GEN_2316 & _GEN_2221 & _GEN_2158 & (~_GEN_1183 & _GEN_1934 | ~_GEN_1179 & _GEN_1869 | (dis_ld_val_3 ? ~_GEN_1397 & _GEN_24865 : ~_GEN_200 & _GEN_24865));
    if (_GEN_1966) begin
      if (_GEN_1901) begin
      end
      else
        ldq_1_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_1_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_2_valid <= ~_GEN_1234 & _GEN_2380 & _GEN_2317 & _GEN_2222 & (_GEN_2156 ? ~_GEN_2031 & _GEN_49602 : ~_GEN_2094 & _GEN_49602);
    if (_GEN_299) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_2_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_2_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_2_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_2_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_2_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_201) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_2_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_2_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_2_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_2_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_134) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_2_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_2_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_2_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_36) begin
      ldq_2_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_2_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_2_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_2_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_2_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_2_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_2_bits_st_dep_mask <= next_live_store_mask;
      ldq_2_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_2_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_2_bits_st_dep_mask;
    if (ldq_2_valid)
      ldq_2_bits_uop_br_mask <= ldq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_299)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_201)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_134)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_36)
      ldq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1651) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_2_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_2_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_2_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_2_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_2_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_2_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_2_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_2_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_2_bits_addr_bits <= hella_req_addr;
        else
          ldq_2_bits_addr_bits <= 40'h0;
      end
      else
        ldq_2_bits_addr_bits <= _GEN_338;
      ldq_2_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_2_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1555) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_2_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_2_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_2_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_2_bits_addr_bits <= _GEN_332;
        else
          ldq_2_bits_addr_bits <= 40'h0;
      end
      else
        ldq_2_bits_addr_bits <= _GEN_334;
      ldq_2_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_2_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_299)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_201)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_134)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_36)
      ldq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_2_bits_addr_valid <= ~_GEN_1234 & _GEN_2380 & _GEN_2317 & _GEN_2222 & (_GEN_2156 ? ~_GEN_2031 & _GEN_81720 : ~_GEN_2094 & _GEN_81720);
    ldq_2_bits_executed <= ~_GEN_1234 & _GEN_2380 & _GEN_2317 & _GEN_2222 & _GEN_2159 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_394) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116697)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1774 & _GEN_113743 : _GEN_1176 ? ~_GEN_1774 & _GEN_113743 : ~(_GEN_113869 & _GEN_1774) & _GEN_113743) : _GEN_113743) | (dis_ld_val_3 ? ~_GEN_1398 & _GEN_24738 : ~_GEN_201 & _GEN_24738));
    ldq_2_bits_succeeded <= _GEN_2380 & _GEN_2317 & _GEN_2222 & _GEN_2159 & (_GEN_1967 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h2 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1902 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h2 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1398 & _GEN_24770 : ~_GEN_201 & _GEN_24770) : casez_tmp_203) : casez_tmp_236);
    ldq_2_bits_order_fail <= _GEN_2380 & _GEN_2317 & _GEN_2222 & _GEN_2159 & (_GEN_397 ? _GEN_84267 : _GEN_399 ? _GEN_400 | _GEN_84267 : _GEN_404 | _GEN_84267);
    ldq_2_bits_observed <= _GEN_397 | (dis_ld_val_3 ? ~_GEN_1398 & _GEN_24834 : ~_GEN_201 & _GEN_24834);
    ldq_2_bits_forward_std_val <= _GEN_2380 & _GEN_2317 & _GEN_2222 & _GEN_2159 & (~_GEN_1183 & _GEN_1935 | ~_GEN_1179 & _GEN_1870 | (dis_ld_val_3 ? ~_GEN_1398 & _GEN_24866 : ~_GEN_201 & _GEN_24866));
    if (_GEN_1967) begin
      if (_GEN_1902) begin
      end
      else
        ldq_2_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_2_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_3_valid <= ~_GEN_1234 & _GEN_2381 & _GEN_2318 & _GEN_2223 & (_GEN_2156 ? ~_GEN_2032 & _GEN_49603 : ~_GEN_2095 & _GEN_49603);
    if (_GEN_300) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_3_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_3_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_3_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_3_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_3_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_202) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_3_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_3_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_3_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_3_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_135) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_3_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_3_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_3_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_37) begin
      ldq_3_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_3_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_3_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_3_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_3_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_3_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_3_bits_st_dep_mask <= next_live_store_mask;
      ldq_3_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_3_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_3_bits_st_dep_mask;
    if (ldq_3_valid)
      ldq_3_bits_uop_br_mask <= ldq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_300)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_202)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_135)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_37)
      ldq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1652) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_3_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_3_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_3_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_3_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_3_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_3_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_3_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_3_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_3_bits_addr_bits <= hella_req_addr;
        else
          ldq_3_bits_addr_bits <= 40'h0;
      end
      else
        ldq_3_bits_addr_bits <= _GEN_338;
      ldq_3_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_3_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1556) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_3_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_3_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_3_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_3_bits_addr_bits <= _GEN_332;
        else
          ldq_3_bits_addr_bits <= 40'h0;
      end
      else
        ldq_3_bits_addr_bits <= _GEN_334;
      ldq_3_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_3_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_300)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_202)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_135)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_37)
      ldq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_3_bits_addr_valid <= ~_GEN_1234 & _GEN_2381 & _GEN_2318 & _GEN_2223 & (_GEN_2156 ? ~_GEN_2032 & _GEN_81721 : ~_GEN_2095 & _GEN_81721);
    ldq_3_bits_executed <= ~_GEN_1234 & _GEN_2381 & _GEN_2318 & _GEN_2223 & _GEN_2160 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_414) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116698)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1775 & _GEN_113744 : _GEN_1176 ? ~_GEN_1775 & _GEN_113744 : ~(_GEN_113869 & _GEN_1775) & _GEN_113744) : _GEN_113744) | (dis_ld_val_3 ? ~_GEN_1399 & _GEN_24739 : ~_GEN_202 & _GEN_24739));
    ldq_3_bits_succeeded <= _GEN_2381 & _GEN_2318 & _GEN_2223 & _GEN_2160 & (_GEN_1968 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h3 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1903 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h3 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1399 & _GEN_24771 : ~_GEN_202 & _GEN_24771) : casez_tmp_203) : casez_tmp_236);
    ldq_3_bits_order_fail <= _GEN_2381 & _GEN_2318 & _GEN_2223 & _GEN_2160 & (_GEN_417 ? _GEN_84765 : _GEN_419 ? _GEN_420 | _GEN_84765 : _GEN_424 | _GEN_84765);
    ldq_3_bits_observed <= _GEN_417 | (dis_ld_val_3 ? ~_GEN_1399 & _GEN_24835 : ~_GEN_202 & _GEN_24835);
    ldq_3_bits_forward_std_val <= _GEN_2381 & _GEN_2318 & _GEN_2223 & _GEN_2160 & (~_GEN_1183 & _GEN_1936 | ~_GEN_1179 & _GEN_1871 | (dis_ld_val_3 ? ~_GEN_1399 & _GEN_24867 : ~_GEN_202 & _GEN_24867));
    if (_GEN_1968) begin
      if (_GEN_1903) begin
      end
      else
        ldq_3_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_3_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_4_valid <= ~_GEN_1234 & _GEN_2382 & _GEN_2319 & _GEN_2224 & (_GEN_2156 ? ~_GEN_2033 & _GEN_49604 : ~_GEN_2096 & _GEN_49604);
    if (_GEN_301) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_4_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_4_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_4_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_4_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_4_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_203) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_4_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_4_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_4_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_4_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_136) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_4_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_4_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_4_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_38) begin
      ldq_4_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_4_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_4_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_4_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_4_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_4_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_4_bits_st_dep_mask <= next_live_store_mask;
      ldq_4_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_4_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_4_bits_st_dep_mask;
    if (ldq_4_valid)
      ldq_4_bits_uop_br_mask <= ldq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_301)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_203)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_136)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_38)
      ldq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1653) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_4_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_4_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_4_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_4_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_4_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_4_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_4_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_4_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_4_bits_addr_bits <= hella_req_addr;
        else
          ldq_4_bits_addr_bits <= 40'h0;
      end
      else
        ldq_4_bits_addr_bits <= _GEN_338;
      ldq_4_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_4_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1557) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_4_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_4_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_4_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_4_bits_addr_bits <= _GEN_332;
        else
          ldq_4_bits_addr_bits <= 40'h0;
      end
      else
        ldq_4_bits_addr_bits <= _GEN_334;
      ldq_4_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_4_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_301)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_203)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_136)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_38)
      ldq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_4_bits_addr_valid <= ~_GEN_1234 & _GEN_2382 & _GEN_2319 & _GEN_2224 & (_GEN_2156 ? ~_GEN_2033 & _GEN_81722 : ~_GEN_2096 & _GEN_81722);
    ldq_4_bits_executed <= ~_GEN_1234 & _GEN_2382 & _GEN_2319 & _GEN_2224 & _GEN_2161 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_434) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116699)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1776 & _GEN_113745 : _GEN_1176 ? ~_GEN_1776 & _GEN_113745 : ~(_GEN_113869 & _GEN_1776) & _GEN_113745) : _GEN_113745) | (dis_ld_val_3 ? ~_GEN_1400 & _GEN_24740 : ~_GEN_203 & _GEN_24740));
    ldq_4_bits_succeeded <= _GEN_2382 & _GEN_2319 & _GEN_2224 & _GEN_2161 & (_GEN_1969 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h4 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1904 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h4 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1400 & _GEN_24772 : ~_GEN_203 & _GEN_24772) : casez_tmp_203) : casez_tmp_236);
    ldq_4_bits_order_fail <= _GEN_2382 & _GEN_2319 & _GEN_2224 & _GEN_2161 & (_GEN_437 ? _GEN_85263 : _GEN_439 ? _GEN_440 | _GEN_85263 : _GEN_444 | _GEN_85263);
    ldq_4_bits_observed <= _GEN_437 | (dis_ld_val_3 ? ~_GEN_1400 & _GEN_24836 : ~_GEN_203 & _GEN_24836);
    ldq_4_bits_forward_std_val <= _GEN_2382 & _GEN_2319 & _GEN_2224 & _GEN_2161 & (~_GEN_1183 & _GEN_1937 | ~_GEN_1179 & _GEN_1872 | (dis_ld_val_3 ? ~_GEN_1400 & _GEN_24868 : ~_GEN_203 & _GEN_24868));
    if (_GEN_1969) begin
      if (_GEN_1904) begin
      end
      else
        ldq_4_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_4_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_5_valid <= ~_GEN_1234 & _GEN_2383 & _GEN_2320 & _GEN_2225 & (_GEN_2156 ? ~_GEN_2034 & _GEN_49605 : ~_GEN_2097 & _GEN_49605);
    if (_GEN_302) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_5_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_5_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_5_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_5_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_5_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_204) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_5_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_5_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_5_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_5_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_137) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_5_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_5_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_5_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_39) begin
      ldq_5_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_5_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_5_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_5_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_5_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_5_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_5_bits_st_dep_mask <= next_live_store_mask;
      ldq_5_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_5_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_5_bits_st_dep_mask;
    if (ldq_5_valid)
      ldq_5_bits_uop_br_mask <= ldq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_302)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_204)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_137)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_39)
      ldq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1654) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_5_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_5_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_5_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_5_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_5_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_5_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_5_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_5_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_5_bits_addr_bits <= hella_req_addr;
        else
          ldq_5_bits_addr_bits <= 40'h0;
      end
      else
        ldq_5_bits_addr_bits <= _GEN_338;
      ldq_5_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_5_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1558) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_5_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_5_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_5_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_5_bits_addr_bits <= _GEN_332;
        else
          ldq_5_bits_addr_bits <= 40'h0;
      end
      else
        ldq_5_bits_addr_bits <= _GEN_334;
      ldq_5_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_5_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_302)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_204)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_137)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_39)
      ldq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_5_bits_addr_valid <= ~_GEN_1234 & _GEN_2383 & _GEN_2320 & _GEN_2225 & (_GEN_2156 ? ~_GEN_2034 & _GEN_81723 : ~_GEN_2097 & _GEN_81723);
    ldq_5_bits_executed <= ~_GEN_1234 & _GEN_2383 & _GEN_2320 & _GEN_2225 & _GEN_2162 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_454) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116700)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1777 & _GEN_113746 : _GEN_1176 ? ~_GEN_1777 & _GEN_113746 : ~(_GEN_113869 & _GEN_1777) & _GEN_113746) : _GEN_113746) | (dis_ld_val_3 ? ~_GEN_1401 & _GEN_24741 : ~_GEN_204 & _GEN_24741));
    ldq_5_bits_succeeded <= _GEN_2383 & _GEN_2320 & _GEN_2225 & _GEN_2162 & (_GEN_1970 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h5 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1905 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h5 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1401 & _GEN_24773 : ~_GEN_204 & _GEN_24773) : casez_tmp_203) : casez_tmp_236);
    ldq_5_bits_order_fail <= _GEN_2383 & _GEN_2320 & _GEN_2225 & _GEN_2162 & (_GEN_457 ? _GEN_85761 : _GEN_459 ? _GEN_460 | _GEN_85761 : _GEN_464 | _GEN_85761);
    ldq_5_bits_observed <= _GEN_457 | (dis_ld_val_3 ? ~_GEN_1401 & _GEN_24837 : ~_GEN_204 & _GEN_24837);
    ldq_5_bits_forward_std_val <= _GEN_2383 & _GEN_2320 & _GEN_2225 & _GEN_2162 & (~_GEN_1183 & _GEN_1938 | ~_GEN_1179 & _GEN_1873 | (dis_ld_val_3 ? ~_GEN_1401 & _GEN_24869 : ~_GEN_204 & _GEN_24869));
    if (_GEN_1970) begin
      if (_GEN_1905) begin
      end
      else
        ldq_5_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_5_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_6_valid <= ~_GEN_1234 & _GEN_2384 & _GEN_2321 & _GEN_2226 & (_GEN_2156 ? ~_GEN_2035 & _GEN_49606 : ~_GEN_2098 & _GEN_49606);
    if (_GEN_303) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_6_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_6_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_6_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_6_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_6_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_205) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_6_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_6_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_6_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_6_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_138) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_6_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_6_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_6_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_40) begin
      ldq_6_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_6_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_6_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_6_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_6_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_6_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_6_bits_st_dep_mask <= next_live_store_mask;
      ldq_6_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_6_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_6_bits_st_dep_mask;
    if (ldq_6_valid)
      ldq_6_bits_uop_br_mask <= ldq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_303)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_205)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_138)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_40)
      ldq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1655) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_6_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_6_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_6_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_6_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_6_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_6_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_6_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_6_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_6_bits_addr_bits <= hella_req_addr;
        else
          ldq_6_bits_addr_bits <= 40'h0;
      end
      else
        ldq_6_bits_addr_bits <= _GEN_338;
      ldq_6_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_6_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1559) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_6_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_6_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_6_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_6_bits_addr_bits <= _GEN_332;
        else
          ldq_6_bits_addr_bits <= 40'h0;
      end
      else
        ldq_6_bits_addr_bits <= _GEN_334;
      ldq_6_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_6_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_303)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_205)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_138)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_40)
      ldq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_6_bits_addr_valid <= ~_GEN_1234 & _GEN_2384 & _GEN_2321 & _GEN_2226 & (_GEN_2156 ? ~_GEN_2035 & _GEN_81724 : ~_GEN_2098 & _GEN_81724);
    ldq_6_bits_executed <= ~_GEN_1234 & _GEN_2384 & _GEN_2321 & _GEN_2226 & _GEN_2163 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_474) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116701)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1778 & _GEN_113747 : _GEN_1176 ? ~_GEN_1778 & _GEN_113747 : ~(_GEN_113869 & _GEN_1778) & _GEN_113747) : _GEN_113747) | (dis_ld_val_3 ? ~_GEN_1402 & _GEN_24742 : ~_GEN_205 & _GEN_24742));
    ldq_6_bits_succeeded <= _GEN_2384 & _GEN_2321 & _GEN_2226 & _GEN_2163 & (_GEN_1971 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h6 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1906 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h6 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1402 & _GEN_24774 : ~_GEN_205 & _GEN_24774) : casez_tmp_203) : casez_tmp_236);
    ldq_6_bits_order_fail <= _GEN_2384 & _GEN_2321 & _GEN_2226 & _GEN_2163 & (_GEN_477 ? _GEN_86259 : _GEN_479 ? _GEN_480 | _GEN_86259 : _GEN_484 | _GEN_86259);
    ldq_6_bits_observed <= _GEN_477 | (dis_ld_val_3 ? ~_GEN_1402 & _GEN_24838 : ~_GEN_205 & _GEN_24838);
    ldq_6_bits_forward_std_val <= _GEN_2384 & _GEN_2321 & _GEN_2226 & _GEN_2163 & (~_GEN_1183 & _GEN_1939 | ~_GEN_1179 & _GEN_1874 | (dis_ld_val_3 ? ~_GEN_1402 & _GEN_24870 : ~_GEN_205 & _GEN_24870));
    if (_GEN_1971) begin
      if (_GEN_1906) begin
      end
      else
        ldq_6_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_6_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_7_valid <= ~_GEN_1234 & _GEN_2385 & _GEN_2322 & _GEN_2227 & (_GEN_2156 ? ~_GEN_2036 & _GEN_49607 : ~_GEN_2099 & _GEN_49607);
    if (_GEN_304) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_7_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_7_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_7_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_7_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_7_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_206) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_7_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_7_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_7_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_7_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_139) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_7_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_7_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_7_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_41) begin
      ldq_7_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_7_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_7_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_7_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_7_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_7_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_7_bits_st_dep_mask <= next_live_store_mask;
      ldq_7_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_7_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_7_bits_st_dep_mask;
    if (ldq_7_valid)
      ldq_7_bits_uop_br_mask <= ldq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_304)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_206)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_139)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_41)
      ldq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1656) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_7_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_7_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_7_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_7_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_7_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_7_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_7_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_7_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_7_bits_addr_bits <= hella_req_addr;
        else
          ldq_7_bits_addr_bits <= 40'h0;
      end
      else
        ldq_7_bits_addr_bits <= _GEN_338;
      ldq_7_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_7_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1560) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_7_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_7_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_7_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_7_bits_addr_bits <= _GEN_332;
        else
          ldq_7_bits_addr_bits <= 40'h0;
      end
      else
        ldq_7_bits_addr_bits <= _GEN_334;
      ldq_7_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_7_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_304)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_206)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_139)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_41)
      ldq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_7_bits_addr_valid <= ~_GEN_1234 & _GEN_2385 & _GEN_2322 & _GEN_2227 & (_GEN_2156 ? ~_GEN_2036 & _GEN_81725 : ~_GEN_2099 & _GEN_81725);
    ldq_7_bits_executed <= ~_GEN_1234 & _GEN_2385 & _GEN_2322 & _GEN_2227 & _GEN_2164 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_494) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116702)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1779 & _GEN_113748 : _GEN_1176 ? ~_GEN_1779 & _GEN_113748 : ~(_GEN_113869 & _GEN_1779) & _GEN_113748) : _GEN_113748) | (dis_ld_val_3 ? ~_GEN_1403 & _GEN_24743 : ~_GEN_206 & _GEN_24743));
    ldq_7_bits_succeeded <= _GEN_2385 & _GEN_2322 & _GEN_2227 & _GEN_2164 & (_GEN_1972 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h7 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1907 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h7 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1403 & _GEN_24775 : ~_GEN_206 & _GEN_24775) : casez_tmp_203) : casez_tmp_236);
    ldq_7_bits_order_fail <= _GEN_2385 & _GEN_2322 & _GEN_2227 & _GEN_2164 & (_GEN_497 ? _GEN_86757 : _GEN_499 ? _GEN_500 | _GEN_86757 : _GEN_504 | _GEN_86757);
    ldq_7_bits_observed <= _GEN_497 | (dis_ld_val_3 ? ~_GEN_1403 & _GEN_24839 : ~_GEN_206 & _GEN_24839);
    ldq_7_bits_forward_std_val <= _GEN_2385 & _GEN_2322 & _GEN_2227 & _GEN_2164 & (~_GEN_1183 & _GEN_1940 | ~_GEN_1179 & _GEN_1875 | (dis_ld_val_3 ? ~_GEN_1403 & _GEN_24871 : ~_GEN_206 & _GEN_24871));
    if (_GEN_1972) begin
      if (_GEN_1907) begin
      end
      else
        ldq_7_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_7_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_8_valid <= ~_GEN_1234 & _GEN_2386 & _GEN_2323 & _GEN_2228 & (_GEN_2156 ? ~_GEN_2037 & _GEN_49608 : ~_GEN_2100 & _GEN_49608);
    if (_GEN_305) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_8_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_8_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_8_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_8_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_8_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_207) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_8_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_8_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_8_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_8_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_140) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_8_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_8_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_8_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_42) begin
      ldq_8_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_8_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_8_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_8_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_8_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_8_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_8_bits_st_dep_mask <= next_live_store_mask;
      ldq_8_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_8_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_8_bits_st_dep_mask;
    if (ldq_8_valid)
      ldq_8_bits_uop_br_mask <= ldq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_305)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_207)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_140)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_42)
      ldq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1657) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_8_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_8_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_8_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_8_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_8_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_8_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_8_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_8_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_8_bits_addr_bits <= hella_req_addr;
        else
          ldq_8_bits_addr_bits <= 40'h0;
      end
      else
        ldq_8_bits_addr_bits <= _GEN_338;
      ldq_8_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_8_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1561) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_8_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_8_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_8_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_8_bits_addr_bits <= _GEN_332;
        else
          ldq_8_bits_addr_bits <= 40'h0;
      end
      else
        ldq_8_bits_addr_bits <= _GEN_334;
      ldq_8_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_8_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_305)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_207)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_140)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_42)
      ldq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_8_bits_addr_valid <= ~_GEN_1234 & _GEN_2386 & _GEN_2323 & _GEN_2228 & (_GEN_2156 ? ~_GEN_2037 & _GEN_81726 : ~_GEN_2100 & _GEN_81726);
    ldq_8_bits_executed <= ~_GEN_1234 & _GEN_2386 & _GEN_2323 & _GEN_2228 & _GEN_2165 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_514) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116703)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1780 & _GEN_113749 : _GEN_1176 ? ~_GEN_1780 & _GEN_113749 : ~(_GEN_113869 & _GEN_1780) & _GEN_113749) : _GEN_113749) | (dis_ld_val_3 ? ~_GEN_1404 & _GEN_24744 : ~_GEN_207 & _GEN_24744));
    ldq_8_bits_succeeded <= _GEN_2386 & _GEN_2323 & _GEN_2228 & _GEN_2165 & (_GEN_1973 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h8 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1908 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h8 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1404 & _GEN_24776 : ~_GEN_207 & _GEN_24776) : casez_tmp_203) : casez_tmp_236);
    ldq_8_bits_order_fail <= _GEN_2386 & _GEN_2323 & _GEN_2228 & _GEN_2165 & (_GEN_517 ? _GEN_87255 : _GEN_519 ? _GEN_520 | _GEN_87255 : _GEN_524 | _GEN_87255);
    ldq_8_bits_observed <= _GEN_517 | (dis_ld_val_3 ? ~_GEN_1404 & _GEN_24840 : ~_GEN_207 & _GEN_24840);
    ldq_8_bits_forward_std_val <= _GEN_2386 & _GEN_2323 & _GEN_2228 & _GEN_2165 & (~_GEN_1183 & _GEN_1941 | ~_GEN_1179 & _GEN_1876 | (dis_ld_val_3 ? ~_GEN_1404 & _GEN_24872 : ~_GEN_207 & _GEN_24872));
    if (_GEN_1973) begin
      if (_GEN_1908) begin
      end
      else
        ldq_8_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_8_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_9_valid <= ~_GEN_1234 & _GEN_2387 & _GEN_2324 & _GEN_2229 & (_GEN_2156 ? ~_GEN_2038 & _GEN_49609 : ~_GEN_2101 & _GEN_49609);
    if (_GEN_306) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_9_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_9_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_9_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_9_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_9_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_208) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_9_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_9_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_9_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_9_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_141) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_9_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_9_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_9_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_43) begin
      ldq_9_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_9_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_9_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_9_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_9_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_9_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_9_bits_st_dep_mask <= next_live_store_mask;
      ldq_9_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_9_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_9_bits_st_dep_mask;
    if (ldq_9_valid)
      ldq_9_bits_uop_br_mask <= ldq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_306)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_208)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_141)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_43)
      ldq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1658) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_9_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_9_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_9_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_9_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_9_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_9_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_9_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_9_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_9_bits_addr_bits <= hella_req_addr;
        else
          ldq_9_bits_addr_bits <= 40'h0;
      end
      else
        ldq_9_bits_addr_bits <= _GEN_338;
      ldq_9_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_9_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1562) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_9_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_9_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_9_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_9_bits_addr_bits <= _GEN_332;
        else
          ldq_9_bits_addr_bits <= 40'h0;
      end
      else
        ldq_9_bits_addr_bits <= _GEN_334;
      ldq_9_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_9_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_306)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_208)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_141)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_43)
      ldq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_9_bits_addr_valid <= ~_GEN_1234 & _GEN_2387 & _GEN_2324 & _GEN_2229 & (_GEN_2156 ? ~_GEN_2038 & _GEN_81727 : ~_GEN_2101 & _GEN_81727);
    ldq_9_bits_executed <= ~_GEN_1234 & _GEN_2387 & _GEN_2324 & _GEN_2229 & _GEN_2166 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_534) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116704)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1781 & _GEN_113750 : _GEN_1176 ? ~_GEN_1781 & _GEN_113750 : ~(_GEN_113869 & _GEN_1781) & _GEN_113750) : _GEN_113750) | (dis_ld_val_3 ? ~_GEN_1405 & _GEN_24745 : ~_GEN_208 & _GEN_24745));
    ldq_9_bits_succeeded <= _GEN_2387 & _GEN_2324 & _GEN_2229 & _GEN_2166 & (_GEN_1974 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h9 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1909 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h9 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1405 & _GEN_24777 : ~_GEN_208 & _GEN_24777) : casez_tmp_203) : casez_tmp_236);
    ldq_9_bits_order_fail <= _GEN_2387 & _GEN_2324 & _GEN_2229 & _GEN_2166 & (_GEN_537 ? _GEN_87753 : _GEN_539 ? _GEN_540 | _GEN_87753 : _GEN_544 | _GEN_87753);
    ldq_9_bits_observed <= _GEN_537 | (dis_ld_val_3 ? ~_GEN_1405 & _GEN_24841 : ~_GEN_208 & _GEN_24841);
    ldq_9_bits_forward_std_val <= _GEN_2387 & _GEN_2324 & _GEN_2229 & _GEN_2166 & (~_GEN_1183 & _GEN_1942 | ~_GEN_1179 & _GEN_1877 | (dis_ld_val_3 ? ~_GEN_1405 & _GEN_24873 : ~_GEN_208 & _GEN_24873));
    if (_GEN_1974) begin
      if (_GEN_1909) begin
      end
      else
        ldq_9_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_9_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_10_valid <= ~_GEN_1234 & _GEN_2388 & _GEN_2325 & _GEN_2230 & (_GEN_2156 ? ~_GEN_2039 & _GEN_49610 : ~_GEN_2102 & _GEN_49610);
    if (_GEN_307) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_10_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_10_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_10_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_10_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_10_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_209) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_10_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_10_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_10_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_10_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_142) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_10_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_10_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_10_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_44) begin
      ldq_10_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_10_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_10_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_10_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_10_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_10_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_10_bits_st_dep_mask <= next_live_store_mask;
      ldq_10_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_10_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_10_bits_st_dep_mask;
    if (ldq_10_valid)
      ldq_10_bits_uop_br_mask <= ldq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_307)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_209)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_142)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_44)
      ldq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1659) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_10_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_10_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_10_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_10_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_10_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_10_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_10_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_10_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_10_bits_addr_bits <= hella_req_addr;
        else
          ldq_10_bits_addr_bits <= 40'h0;
      end
      else
        ldq_10_bits_addr_bits <= _GEN_338;
      ldq_10_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_10_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1563) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_10_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_10_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_10_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_10_bits_addr_bits <= _GEN_332;
        else
          ldq_10_bits_addr_bits <= 40'h0;
      end
      else
        ldq_10_bits_addr_bits <= _GEN_334;
      ldq_10_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_10_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_307)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_209)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_142)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_44)
      ldq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_10_bits_addr_valid <= ~_GEN_1234 & _GEN_2388 & _GEN_2325 & _GEN_2230 & (_GEN_2156 ? ~_GEN_2039 & _GEN_81728 : ~_GEN_2102 & _GEN_81728);
    ldq_10_bits_executed <= ~_GEN_1234 & _GEN_2388 & _GEN_2325 & _GEN_2230 & _GEN_2167 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_554) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116705)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1782 & _GEN_113751 : _GEN_1176 ? ~_GEN_1782 & _GEN_113751 : ~(_GEN_113869 & _GEN_1782) & _GEN_113751) : _GEN_113751) | (dis_ld_val_3 ? ~_GEN_1406 & _GEN_24746 : ~_GEN_209 & _GEN_24746));
    ldq_10_bits_succeeded <= _GEN_2388 & _GEN_2325 & _GEN_2230 & _GEN_2167 & (_GEN_1975 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hA ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1910 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hA ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1406 & _GEN_24778 : ~_GEN_209 & _GEN_24778) : casez_tmp_203) : casez_tmp_236);
    ldq_10_bits_order_fail <= _GEN_2388 & _GEN_2325 & _GEN_2230 & _GEN_2167 & (_GEN_557 ? _GEN_88251 : _GEN_559 ? _GEN_560 | _GEN_88251 : _GEN_564 | _GEN_88251);
    ldq_10_bits_observed <= _GEN_557 | (dis_ld_val_3 ? ~_GEN_1406 & _GEN_24842 : ~_GEN_209 & _GEN_24842);
    ldq_10_bits_forward_std_val <= _GEN_2388 & _GEN_2325 & _GEN_2230 & _GEN_2167 & (~_GEN_1183 & _GEN_1943 | ~_GEN_1179 & _GEN_1878 | (dis_ld_val_3 ? ~_GEN_1406 & _GEN_24874 : ~_GEN_209 & _GEN_24874));
    if (_GEN_1975) begin
      if (_GEN_1910) begin
      end
      else
        ldq_10_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_10_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_11_valid <= ~_GEN_1234 & _GEN_2389 & _GEN_2326 & _GEN_2231 & (_GEN_2156 ? ~_GEN_2040 & _GEN_49611 : ~_GEN_2103 & _GEN_49611);
    if (_GEN_308) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_11_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_11_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_11_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_11_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_11_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_210) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_11_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_11_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_11_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_11_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_143) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_11_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_11_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_11_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_45) begin
      ldq_11_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_11_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_11_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_11_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_11_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_11_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_11_bits_st_dep_mask <= next_live_store_mask;
      ldq_11_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_11_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_11_bits_st_dep_mask;
    if (ldq_11_valid)
      ldq_11_bits_uop_br_mask <= ldq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_308)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_210)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_143)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_45)
      ldq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1660) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_11_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_11_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_11_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_11_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_11_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_11_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_11_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_11_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_11_bits_addr_bits <= hella_req_addr;
        else
          ldq_11_bits_addr_bits <= 40'h0;
      end
      else
        ldq_11_bits_addr_bits <= _GEN_338;
      ldq_11_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_11_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1564) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_11_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_11_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_11_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_11_bits_addr_bits <= _GEN_332;
        else
          ldq_11_bits_addr_bits <= 40'h0;
      end
      else
        ldq_11_bits_addr_bits <= _GEN_334;
      ldq_11_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_11_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_308)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_210)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_143)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_45)
      ldq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_11_bits_addr_valid <= ~_GEN_1234 & _GEN_2389 & _GEN_2326 & _GEN_2231 & (_GEN_2156 ? ~_GEN_2040 & _GEN_81729 : ~_GEN_2103 & _GEN_81729);
    ldq_11_bits_executed <= ~_GEN_1234 & _GEN_2389 & _GEN_2326 & _GEN_2231 & _GEN_2168 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_574) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116706)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1783 & _GEN_113752 : _GEN_1176 ? ~_GEN_1783 & _GEN_113752 : ~(_GEN_113869 & _GEN_1783) & _GEN_113752) : _GEN_113752) | (dis_ld_val_3 ? ~_GEN_1407 & _GEN_24747 : ~_GEN_210 & _GEN_24747));
    ldq_11_bits_succeeded <= _GEN_2389 & _GEN_2326 & _GEN_2231 & _GEN_2168 & (_GEN_1976 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hB ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1911 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hB ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1407 & _GEN_24779 : ~_GEN_210 & _GEN_24779) : casez_tmp_203) : casez_tmp_236);
    ldq_11_bits_order_fail <= _GEN_2389 & _GEN_2326 & _GEN_2231 & _GEN_2168 & (_GEN_577 ? _GEN_88749 : _GEN_579 ? _GEN_580 | _GEN_88749 : _GEN_584 | _GEN_88749);
    ldq_11_bits_observed <= _GEN_577 | (dis_ld_val_3 ? ~_GEN_1407 & _GEN_24843 : ~_GEN_210 & _GEN_24843);
    ldq_11_bits_forward_std_val <= _GEN_2389 & _GEN_2326 & _GEN_2231 & _GEN_2168 & (~_GEN_1183 & _GEN_1944 | ~_GEN_1179 & _GEN_1879 | (dis_ld_val_3 ? ~_GEN_1407 & _GEN_24875 : ~_GEN_210 & _GEN_24875));
    if (_GEN_1976) begin
      if (_GEN_1911) begin
      end
      else
        ldq_11_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_11_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_12_valid <= ~_GEN_1234 & _GEN_2390 & _GEN_2327 & _GEN_2232 & (_GEN_2156 ? ~_GEN_2041 & _GEN_49612 : ~_GEN_2104 & _GEN_49612);
    if (_GEN_309) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_12_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_12_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_12_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_12_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_12_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_211) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_12_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_12_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_12_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_12_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_144) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_12_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_12_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_12_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_46) begin
      ldq_12_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_12_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_12_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_12_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_12_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_12_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_12_bits_st_dep_mask <= next_live_store_mask;
      ldq_12_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_12_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_12_bits_st_dep_mask;
    if (ldq_12_valid)
      ldq_12_bits_uop_br_mask <= ldq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_309)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_211)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_144)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_46)
      ldq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1661) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_12_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_12_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_12_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_12_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_12_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_12_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_12_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_12_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_12_bits_addr_bits <= hella_req_addr;
        else
          ldq_12_bits_addr_bits <= 40'h0;
      end
      else
        ldq_12_bits_addr_bits <= _GEN_338;
      ldq_12_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_12_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1565) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_12_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_12_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_12_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_12_bits_addr_bits <= _GEN_332;
        else
          ldq_12_bits_addr_bits <= 40'h0;
      end
      else
        ldq_12_bits_addr_bits <= _GEN_334;
      ldq_12_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_12_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_309)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_211)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_144)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_46)
      ldq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_12_bits_addr_valid <= ~_GEN_1234 & _GEN_2390 & _GEN_2327 & _GEN_2232 & (_GEN_2156 ? ~_GEN_2041 & _GEN_81730 : ~_GEN_2104 & _GEN_81730);
    ldq_12_bits_executed <= ~_GEN_1234 & _GEN_2390 & _GEN_2327 & _GEN_2232 & _GEN_2169 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_594) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116707)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1784 & _GEN_113753 : _GEN_1176 ? ~_GEN_1784 & _GEN_113753 : ~(_GEN_113869 & _GEN_1784) & _GEN_113753) : _GEN_113753) | (dis_ld_val_3 ? ~_GEN_1408 & _GEN_24748 : ~_GEN_211 & _GEN_24748));
    ldq_12_bits_succeeded <= _GEN_2390 & _GEN_2327 & _GEN_2232 & _GEN_2169 & (_GEN_1977 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hC ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1912 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hC ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1408 & _GEN_24780 : ~_GEN_211 & _GEN_24780) : casez_tmp_203) : casez_tmp_236);
    ldq_12_bits_order_fail <= _GEN_2390 & _GEN_2327 & _GEN_2232 & _GEN_2169 & (_GEN_597 ? _GEN_89247 : _GEN_599 ? _GEN_600 | _GEN_89247 : _GEN_604 | _GEN_89247);
    ldq_12_bits_observed <= _GEN_597 | (dis_ld_val_3 ? ~_GEN_1408 & _GEN_24844 : ~_GEN_211 & _GEN_24844);
    ldq_12_bits_forward_std_val <= _GEN_2390 & _GEN_2327 & _GEN_2232 & _GEN_2169 & (~_GEN_1183 & _GEN_1945 | ~_GEN_1179 & _GEN_1880 | (dis_ld_val_3 ? ~_GEN_1408 & _GEN_24876 : ~_GEN_211 & _GEN_24876));
    if (_GEN_1977) begin
      if (_GEN_1912) begin
      end
      else
        ldq_12_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_12_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_13_valid <= ~_GEN_1234 & _GEN_2391 & _GEN_2328 & _GEN_2233 & (_GEN_2156 ? ~_GEN_2042 & _GEN_49613 : ~_GEN_2105 & _GEN_49613);
    if (_GEN_310) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_13_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_13_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_13_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_13_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_13_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_212) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_13_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_13_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_13_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_13_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_145) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_13_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_13_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_13_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_47) begin
      ldq_13_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_13_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_13_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_13_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_13_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_13_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_13_bits_st_dep_mask <= next_live_store_mask;
      ldq_13_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_13_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_13_bits_st_dep_mask;
    if (ldq_13_valid)
      ldq_13_bits_uop_br_mask <= ldq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_310)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_212)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_145)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_47)
      ldq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1662) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_13_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_13_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_13_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_13_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_13_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_13_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_13_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_13_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_13_bits_addr_bits <= hella_req_addr;
        else
          ldq_13_bits_addr_bits <= 40'h0;
      end
      else
        ldq_13_bits_addr_bits <= _GEN_338;
      ldq_13_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_13_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1566) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_13_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_13_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_13_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_13_bits_addr_bits <= _GEN_332;
        else
          ldq_13_bits_addr_bits <= 40'h0;
      end
      else
        ldq_13_bits_addr_bits <= _GEN_334;
      ldq_13_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_13_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_310)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_212)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_145)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_47)
      ldq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_13_bits_addr_valid <= ~_GEN_1234 & _GEN_2391 & _GEN_2328 & _GEN_2233 & (_GEN_2156 ? ~_GEN_2042 & _GEN_81731 : ~_GEN_2105 & _GEN_81731);
    ldq_13_bits_executed <= ~_GEN_1234 & _GEN_2391 & _GEN_2328 & _GEN_2233 & _GEN_2170 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_614) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116708)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1785 & _GEN_113754 : _GEN_1176 ? ~_GEN_1785 & _GEN_113754 : ~(_GEN_113869 & _GEN_1785) & _GEN_113754) : _GEN_113754) | (dis_ld_val_3 ? ~_GEN_1409 & _GEN_24749 : ~_GEN_212 & _GEN_24749));
    ldq_13_bits_succeeded <= _GEN_2391 & _GEN_2328 & _GEN_2233 & _GEN_2170 & (_GEN_1978 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hD ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1913 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hD ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1409 & _GEN_24781 : ~_GEN_212 & _GEN_24781) : casez_tmp_203) : casez_tmp_236);
    ldq_13_bits_order_fail <= _GEN_2391 & _GEN_2328 & _GEN_2233 & _GEN_2170 & (_GEN_617 ? _GEN_89745 : _GEN_619 ? _GEN_620 | _GEN_89745 : _GEN_624 | _GEN_89745);
    ldq_13_bits_observed <= _GEN_617 | (dis_ld_val_3 ? ~_GEN_1409 & _GEN_24845 : ~_GEN_212 & _GEN_24845);
    ldq_13_bits_forward_std_val <= _GEN_2391 & _GEN_2328 & _GEN_2233 & _GEN_2170 & (~_GEN_1183 & _GEN_1946 | ~_GEN_1179 & _GEN_1881 | (dis_ld_val_3 ? ~_GEN_1409 & _GEN_24877 : ~_GEN_212 & _GEN_24877));
    if (_GEN_1978) begin
      if (_GEN_1913) begin
      end
      else
        ldq_13_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_13_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_14_valid <= ~_GEN_1234 & _GEN_2392 & _GEN_2329 & _GEN_2234 & (_GEN_2156 ? ~_GEN_2043 & _GEN_49614 : ~_GEN_2106 & _GEN_49614);
    if (_GEN_311) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_14_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_14_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_14_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_14_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_14_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_213) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_14_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_14_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_14_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_14_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_146) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_14_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_14_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_14_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_48) begin
      ldq_14_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_14_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_14_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_14_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_14_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_14_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_14_bits_st_dep_mask <= next_live_store_mask;
      ldq_14_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_14_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_14_bits_st_dep_mask;
    if (ldq_14_valid)
      ldq_14_bits_uop_br_mask <= ldq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_311)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_213)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_146)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_48)
      ldq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1663) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_14_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_14_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_14_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_14_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_14_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_14_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_14_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_14_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_14_bits_addr_bits <= hella_req_addr;
        else
          ldq_14_bits_addr_bits <= 40'h0;
      end
      else
        ldq_14_bits_addr_bits <= _GEN_338;
      ldq_14_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_14_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1567) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_14_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_14_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_14_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_14_bits_addr_bits <= _GEN_332;
        else
          ldq_14_bits_addr_bits <= 40'h0;
      end
      else
        ldq_14_bits_addr_bits <= _GEN_334;
      ldq_14_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_14_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_311)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_213)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_146)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_48)
      ldq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_14_bits_addr_valid <= ~_GEN_1234 & _GEN_2392 & _GEN_2329 & _GEN_2234 & (_GEN_2156 ? ~_GEN_2043 & _GEN_81732 : ~_GEN_2106 & _GEN_81732);
    ldq_14_bits_executed <= ~_GEN_1234 & _GEN_2392 & _GEN_2329 & _GEN_2234 & _GEN_2171 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_634) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116709)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1786 & _GEN_113755 : _GEN_1176 ? ~_GEN_1786 & _GEN_113755 : ~(_GEN_113869 & _GEN_1786) & _GEN_113755) : _GEN_113755) | (dis_ld_val_3 ? ~_GEN_1410 & _GEN_24750 : ~_GEN_213 & _GEN_24750));
    ldq_14_bits_succeeded <= _GEN_2392 & _GEN_2329 & _GEN_2234 & _GEN_2171 & (_GEN_1979 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hE ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1914 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hE ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1410 & _GEN_24782 : ~_GEN_213 & _GEN_24782) : casez_tmp_203) : casez_tmp_236);
    ldq_14_bits_order_fail <= _GEN_2392 & _GEN_2329 & _GEN_2234 & _GEN_2171 & (_GEN_637 ? _GEN_90243 : _GEN_639 ? _GEN_640 | _GEN_90243 : _GEN_644 | _GEN_90243);
    ldq_14_bits_observed <= _GEN_637 | (dis_ld_val_3 ? ~_GEN_1410 & _GEN_24846 : ~_GEN_213 & _GEN_24846);
    ldq_14_bits_forward_std_val <= _GEN_2392 & _GEN_2329 & _GEN_2234 & _GEN_2171 & (~_GEN_1183 & _GEN_1947 | ~_GEN_1179 & _GEN_1882 | (dis_ld_val_3 ? ~_GEN_1410 & _GEN_24878 : ~_GEN_213 & _GEN_24878));
    if (_GEN_1979) begin
      if (_GEN_1914) begin
      end
      else
        ldq_14_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_14_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_15_valid <= ~_GEN_1234 & _GEN_2393 & _GEN_2330 & _GEN_2235 & (_GEN_2156 ? ~_GEN_2044 & _GEN_49615 : ~_GEN_2107 & _GEN_49615);
    if (_GEN_312) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_15_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_15_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_15_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_15_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_15_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_214) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_15_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_15_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_15_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_15_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_147) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_15_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_15_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_15_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_49) begin
      ldq_15_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_15_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_15_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_15_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_15_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_15_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_15_bits_st_dep_mask <= next_live_store_mask;
      ldq_15_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_15_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_15_bits_st_dep_mask;
    if (ldq_15_valid)
      ldq_15_bits_uop_br_mask <= ldq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_312)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_214)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_147)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_49)
      ldq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1664) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_15_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_15_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_15_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_15_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_15_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_15_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_15_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_15_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_15_bits_addr_bits <= hella_req_addr;
        else
          ldq_15_bits_addr_bits <= 40'h0;
      end
      else
        ldq_15_bits_addr_bits <= _GEN_338;
      ldq_15_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_15_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1568) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_15_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_15_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_15_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_15_bits_addr_bits <= _GEN_332;
        else
          ldq_15_bits_addr_bits <= 40'h0;
      end
      else
        ldq_15_bits_addr_bits <= _GEN_334;
      ldq_15_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_15_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_312)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_214)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_147)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_49)
      ldq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_15_bits_addr_valid <= ~_GEN_1234 & _GEN_2393 & _GEN_2330 & _GEN_2235 & (_GEN_2156 ? ~_GEN_2044 & _GEN_81733 : ~_GEN_2107 & _GEN_81733);
    ldq_15_bits_executed <= ~_GEN_1234 & _GEN_2393 & _GEN_2330 & _GEN_2235 & _GEN_2172 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_654) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116710)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1787 & _GEN_113756 : _GEN_1176 ? ~_GEN_1787 & _GEN_113756 : ~(_GEN_113869 & _GEN_1787) & _GEN_113756) : _GEN_113756) | (dis_ld_val_3 ? ~_GEN_1411 & _GEN_24751 : ~_GEN_214 & _GEN_24751));
    ldq_15_bits_succeeded <= _GEN_2393 & _GEN_2330 & _GEN_2235 & _GEN_2172 & (_GEN_1980 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'hF ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1915 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'hF ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1411 & _GEN_24783 : ~_GEN_214 & _GEN_24783) : casez_tmp_203) : casez_tmp_236);
    ldq_15_bits_order_fail <= _GEN_2393 & _GEN_2330 & _GEN_2235 & _GEN_2172 & (_GEN_657 ? _GEN_90741 : _GEN_659 ? _GEN_660 | _GEN_90741 : _GEN_664 | _GEN_90741);
    ldq_15_bits_observed <= _GEN_657 | (dis_ld_val_3 ? ~_GEN_1411 & _GEN_24847 : ~_GEN_214 & _GEN_24847);
    ldq_15_bits_forward_std_val <= _GEN_2393 & _GEN_2330 & _GEN_2235 & _GEN_2172 & (~_GEN_1183 & _GEN_1948 | ~_GEN_1179 & _GEN_1883 | (dis_ld_val_3 ? ~_GEN_1411 & _GEN_24879 : ~_GEN_214 & _GEN_24879));
    if (_GEN_1980) begin
      if (_GEN_1915) begin
      end
      else
        ldq_15_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_15_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_16_valid <= ~_GEN_1234 & _GEN_2394 & _GEN_2331 & _GEN_2236 & (_GEN_2156 ? ~_GEN_2045 & _GEN_49616 : ~_GEN_2108 & _GEN_49616);
    if (_GEN_313) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_16_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_16_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_16_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_16_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_16_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_215) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_16_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_16_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_16_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_16_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_148) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_16_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_16_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_16_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_50) begin
      ldq_16_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_16_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_16_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_16_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_16_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_16_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_16_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_16_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_16_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_16_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_16_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_16_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_16_bits_st_dep_mask <= next_live_store_mask;
      ldq_16_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_16_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_16_bits_st_dep_mask;
    if (ldq_16_valid)
      ldq_16_bits_uop_br_mask <= ldq_16_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_313)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_215)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_148)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_50)
      ldq_16_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1665) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_16_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_16_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_16_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_16_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_16_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_16_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_16_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_16_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_16_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_16_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_16_bits_addr_bits <= hella_req_addr;
        else
          ldq_16_bits_addr_bits <= 40'h0;
      end
      else
        ldq_16_bits_addr_bits <= _GEN_338;
      ldq_16_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_16_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1569) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_16_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_16_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_16_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_16_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_16_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_16_bits_addr_bits <= _GEN_332;
        else
          ldq_16_bits_addr_bits <= 40'h0;
      end
      else
        ldq_16_bits_addr_bits <= _GEN_334;
      ldq_16_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_16_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_313)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_215)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_148)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_50)
      ldq_16_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_16_bits_addr_valid <= ~_GEN_1234 & _GEN_2394 & _GEN_2331 & _GEN_2236 & (_GEN_2156 ? ~_GEN_2045 & _GEN_81734 : ~_GEN_2108 & _GEN_81734);
    ldq_16_bits_executed <= ~_GEN_1234 & _GEN_2394 & _GEN_2331 & _GEN_2236 & _GEN_2173 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_674) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116711)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1788 & _GEN_113757 : _GEN_1176 ? ~_GEN_1788 & _GEN_113757 : ~(_GEN_113869 & _GEN_1788) & _GEN_113757) : _GEN_113757) | (dis_ld_val_3 ? ~_GEN_1412 & _GEN_24752 : ~_GEN_215 & _GEN_24752));
    ldq_16_bits_succeeded <= _GEN_2394 & _GEN_2331 & _GEN_2236 & _GEN_2173 & (_GEN_1981 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h10 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1916 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h10 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1412 & _GEN_24784 : ~_GEN_215 & _GEN_24784) : casez_tmp_203) : casez_tmp_236);
    ldq_16_bits_order_fail <= _GEN_2394 & _GEN_2331 & _GEN_2236 & _GEN_2173 & (_GEN_677 ? _GEN_91239 : _GEN_679 ? _GEN_680 | _GEN_91239 : _GEN_684 | _GEN_91239);
    ldq_16_bits_observed <= _GEN_677 | (dis_ld_val_3 ? ~_GEN_1412 & _GEN_24848 : ~_GEN_215 & _GEN_24848);
    ldq_16_bits_forward_std_val <= _GEN_2394 & _GEN_2331 & _GEN_2236 & _GEN_2173 & (~_GEN_1183 & _GEN_1949 | ~_GEN_1179 & _GEN_1884 | (dis_ld_val_3 ? ~_GEN_1412 & _GEN_24880 : ~_GEN_215 & _GEN_24880));
    if (_GEN_1981) begin
      if (_GEN_1916) begin
      end
      else
        ldq_16_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_16_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_17_valid <= ~_GEN_1234 & _GEN_2395 & _GEN_2332 & _GEN_2237 & (_GEN_2156 ? ~_GEN_2046 & _GEN_49617 : ~_GEN_2109 & _GEN_49617);
    if (_GEN_314) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_17_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_17_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_17_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_17_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_17_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_216) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_17_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_17_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_17_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_17_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_149) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_17_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_17_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_17_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_51) begin
      ldq_17_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_17_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_17_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_17_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_17_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_17_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_17_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_17_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_17_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_17_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_17_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_17_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_17_bits_st_dep_mask <= next_live_store_mask;
      ldq_17_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_17_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_17_bits_st_dep_mask;
    if (ldq_17_valid)
      ldq_17_bits_uop_br_mask <= ldq_17_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_314)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_216)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_149)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_51)
      ldq_17_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1666) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_17_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_17_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_17_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_17_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_17_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_17_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_17_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_17_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_17_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_17_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_17_bits_addr_bits <= hella_req_addr;
        else
          ldq_17_bits_addr_bits <= 40'h0;
      end
      else
        ldq_17_bits_addr_bits <= _GEN_338;
      ldq_17_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_17_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1570) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_17_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_17_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_17_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_17_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_17_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_17_bits_addr_bits <= _GEN_332;
        else
          ldq_17_bits_addr_bits <= 40'h0;
      end
      else
        ldq_17_bits_addr_bits <= _GEN_334;
      ldq_17_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_17_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_314)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_216)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_149)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_51)
      ldq_17_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_17_bits_addr_valid <= ~_GEN_1234 & _GEN_2395 & _GEN_2332 & _GEN_2237 & (_GEN_2156 ? ~_GEN_2046 & _GEN_81735 : ~_GEN_2109 & _GEN_81735);
    ldq_17_bits_executed <= ~_GEN_1234 & _GEN_2395 & _GEN_2332 & _GEN_2237 & _GEN_2174 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_694) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116712)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1789 & _GEN_113758 : _GEN_1176 ? ~_GEN_1789 & _GEN_113758 : ~(_GEN_113869 & _GEN_1789) & _GEN_113758) : _GEN_113758) | (dis_ld_val_3 ? ~_GEN_1413 & _GEN_24753 : ~_GEN_216 & _GEN_24753));
    ldq_17_bits_succeeded <= _GEN_2395 & _GEN_2332 & _GEN_2237 & _GEN_2174 & (_GEN_1982 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h11 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1917 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h11 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1413 & _GEN_24785 : ~_GEN_216 & _GEN_24785) : casez_tmp_203) : casez_tmp_236);
    ldq_17_bits_order_fail <= _GEN_2395 & _GEN_2332 & _GEN_2237 & _GEN_2174 & (_GEN_697 ? _GEN_91737 : _GEN_699 ? _GEN_700 | _GEN_91737 : _GEN_704 | _GEN_91737);
    ldq_17_bits_observed <= _GEN_697 | (dis_ld_val_3 ? ~_GEN_1413 & _GEN_24849 : ~_GEN_216 & _GEN_24849);
    ldq_17_bits_forward_std_val <= _GEN_2395 & _GEN_2332 & _GEN_2237 & _GEN_2174 & (~_GEN_1183 & _GEN_1950 | ~_GEN_1179 & _GEN_1885 | (dis_ld_val_3 ? ~_GEN_1413 & _GEN_24881 : ~_GEN_216 & _GEN_24881));
    if (_GEN_1982) begin
      if (_GEN_1917) begin
      end
      else
        ldq_17_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_17_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_18_valid <= ~_GEN_1234 & _GEN_2396 & _GEN_2333 & _GEN_2238 & (_GEN_2156 ? ~_GEN_2047 & _GEN_49618 : ~_GEN_2110 & _GEN_49618);
    if (_GEN_315) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_18_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_18_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_18_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_18_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_18_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_217) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_18_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_18_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_18_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_18_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_150) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_18_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_18_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_18_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_52) begin
      ldq_18_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_18_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_18_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_18_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_18_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_18_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_18_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_18_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_18_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_18_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_18_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_18_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_18_bits_st_dep_mask <= next_live_store_mask;
      ldq_18_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_18_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_18_bits_st_dep_mask;
    if (ldq_18_valid)
      ldq_18_bits_uop_br_mask <= ldq_18_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_315)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_217)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_150)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_52)
      ldq_18_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1667) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_18_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_18_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_18_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_18_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_18_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_18_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_18_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_18_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_18_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_18_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_18_bits_addr_bits <= hella_req_addr;
        else
          ldq_18_bits_addr_bits <= 40'h0;
      end
      else
        ldq_18_bits_addr_bits <= _GEN_338;
      ldq_18_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_18_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1571) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_18_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_18_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_18_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_18_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_18_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_18_bits_addr_bits <= _GEN_332;
        else
          ldq_18_bits_addr_bits <= 40'h0;
      end
      else
        ldq_18_bits_addr_bits <= _GEN_334;
      ldq_18_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_18_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_315)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_217)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_150)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_52)
      ldq_18_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_18_bits_addr_valid <= ~_GEN_1234 & _GEN_2396 & _GEN_2333 & _GEN_2238 & (_GEN_2156 ? ~_GEN_2047 & _GEN_81736 : ~_GEN_2110 & _GEN_81736);
    ldq_18_bits_executed <= ~_GEN_1234 & _GEN_2396 & _GEN_2333 & _GEN_2238 & _GEN_2175 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_714) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116713)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1790 & _GEN_113759 : _GEN_1176 ? ~_GEN_1790 & _GEN_113759 : ~(_GEN_113869 & _GEN_1790) & _GEN_113759) : _GEN_113759) | (dis_ld_val_3 ? ~_GEN_1414 & _GEN_24754 : ~_GEN_217 & _GEN_24754));
    ldq_18_bits_succeeded <= _GEN_2396 & _GEN_2333 & _GEN_2238 & _GEN_2175 & (_GEN_1983 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h12 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1918 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h12 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1414 & _GEN_24786 : ~_GEN_217 & _GEN_24786) : casez_tmp_203) : casez_tmp_236);
    ldq_18_bits_order_fail <= _GEN_2396 & _GEN_2333 & _GEN_2238 & _GEN_2175 & (_GEN_717 ? _GEN_92235 : _GEN_719 ? _GEN_720 | _GEN_92235 : _GEN_724 | _GEN_92235);
    ldq_18_bits_observed <= _GEN_717 | (dis_ld_val_3 ? ~_GEN_1414 & _GEN_24850 : ~_GEN_217 & _GEN_24850);
    ldq_18_bits_forward_std_val <= _GEN_2396 & _GEN_2333 & _GEN_2238 & _GEN_2175 & (~_GEN_1183 & _GEN_1951 | ~_GEN_1179 & _GEN_1886 | (dis_ld_val_3 ? ~_GEN_1414 & _GEN_24882 : ~_GEN_217 & _GEN_24882));
    if (_GEN_1983) begin
      if (_GEN_1918) begin
      end
      else
        ldq_18_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_18_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_19_valid <= ~_GEN_1234 & _GEN_2397 & _GEN_2334 & _GEN_2239 & (_GEN_2156 ? ~_GEN_2048 & _GEN_49619 : ~_GEN_2111 & _GEN_49619);
    if (_GEN_316) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_19_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_19_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_19_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_19_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_19_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_218) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_19_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_19_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_19_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_19_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_151) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_19_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_19_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_19_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_53) begin
      ldq_19_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_19_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_19_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_19_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_19_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_19_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_19_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_19_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_19_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_19_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_19_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_19_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_19_bits_st_dep_mask <= next_live_store_mask;
      ldq_19_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_19_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_19_bits_st_dep_mask;
    if (ldq_19_valid)
      ldq_19_bits_uop_br_mask <= ldq_19_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_316)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_218)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_151)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_53)
      ldq_19_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1668) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_19_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_19_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_19_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_19_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_19_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_19_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_19_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_19_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_19_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_19_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_19_bits_addr_bits <= hella_req_addr;
        else
          ldq_19_bits_addr_bits <= 40'h0;
      end
      else
        ldq_19_bits_addr_bits <= _GEN_338;
      ldq_19_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_19_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1572) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_19_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_19_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_19_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_19_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_19_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_19_bits_addr_bits <= _GEN_332;
        else
          ldq_19_bits_addr_bits <= 40'h0;
      end
      else
        ldq_19_bits_addr_bits <= _GEN_334;
      ldq_19_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_19_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_316)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_218)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_151)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_53)
      ldq_19_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_19_bits_addr_valid <= ~_GEN_1234 & _GEN_2397 & _GEN_2334 & _GEN_2239 & (_GEN_2156 ? ~_GEN_2048 & _GEN_81737 : ~_GEN_2111 & _GEN_81737);
    ldq_19_bits_executed <= ~_GEN_1234 & _GEN_2397 & _GEN_2334 & _GEN_2239 & _GEN_2176 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_734) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116714)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1791 & _GEN_113760 : _GEN_1176 ? ~_GEN_1791 & _GEN_113760 : ~(_GEN_113869 & _GEN_1791) & _GEN_113760) : _GEN_113760) | (dis_ld_val_3 ? ~_GEN_1415 & _GEN_24755 : ~_GEN_218 & _GEN_24755));
    ldq_19_bits_succeeded <= _GEN_2397 & _GEN_2334 & _GEN_2239 & _GEN_2176 & (_GEN_1984 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h13 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1919 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h13 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1415 & _GEN_24787 : ~_GEN_218 & _GEN_24787) : casez_tmp_203) : casez_tmp_236);
    ldq_19_bits_order_fail <= _GEN_2397 & _GEN_2334 & _GEN_2239 & _GEN_2176 & (_GEN_737 ? _GEN_92733 : _GEN_739 ? _GEN_740 | _GEN_92733 : _GEN_744 | _GEN_92733);
    ldq_19_bits_observed <= _GEN_737 | (dis_ld_val_3 ? ~_GEN_1415 & _GEN_24851 : ~_GEN_218 & _GEN_24851);
    ldq_19_bits_forward_std_val <= _GEN_2397 & _GEN_2334 & _GEN_2239 & _GEN_2176 & (~_GEN_1183 & _GEN_1952 | ~_GEN_1179 & _GEN_1887 | (dis_ld_val_3 ? ~_GEN_1415 & _GEN_24883 : ~_GEN_218 & _GEN_24883));
    if (_GEN_1984) begin
      if (_GEN_1919) begin
      end
      else
        ldq_19_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_19_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_20_valid <= ~_GEN_1234 & _GEN_2398 & _GEN_2335 & _GEN_2240 & (_GEN_2156 ? ~_GEN_2049 & _GEN_49620 : ~_GEN_2112 & _GEN_49620);
    if (_GEN_317) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_20_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_20_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_20_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_20_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_20_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_219) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_20_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_20_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_20_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_20_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_152) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_20_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_20_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_20_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_54) begin
      ldq_20_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_20_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_20_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_20_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_20_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_20_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_20_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_20_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_20_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_20_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_20_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_20_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_20_bits_st_dep_mask <= next_live_store_mask;
      ldq_20_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_20_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_20_bits_st_dep_mask;
    if (ldq_20_valid)
      ldq_20_bits_uop_br_mask <= ldq_20_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_317)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_219)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_152)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_54)
      ldq_20_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1669) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_20_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_20_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_20_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_20_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_20_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_20_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_20_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_20_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_20_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_20_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_20_bits_addr_bits <= hella_req_addr;
        else
          ldq_20_bits_addr_bits <= 40'h0;
      end
      else
        ldq_20_bits_addr_bits <= _GEN_338;
      ldq_20_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_20_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1573) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_20_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_20_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_20_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_20_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_20_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_20_bits_addr_bits <= _GEN_332;
        else
          ldq_20_bits_addr_bits <= 40'h0;
      end
      else
        ldq_20_bits_addr_bits <= _GEN_334;
      ldq_20_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_20_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_317)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_219)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_152)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_54)
      ldq_20_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_20_bits_addr_valid <= ~_GEN_1234 & _GEN_2398 & _GEN_2335 & _GEN_2240 & (_GEN_2156 ? ~_GEN_2049 & _GEN_81738 : ~_GEN_2112 & _GEN_81738);
    ldq_20_bits_executed <= ~_GEN_1234 & _GEN_2398 & _GEN_2335 & _GEN_2240 & _GEN_2177 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_754) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116715)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1792 & _GEN_113761 : _GEN_1176 ? ~_GEN_1792 & _GEN_113761 : ~(_GEN_113869 & _GEN_1792) & _GEN_113761) : _GEN_113761) | (dis_ld_val_3 ? ~_GEN_1416 & _GEN_24756 : ~_GEN_219 & _GEN_24756));
    ldq_20_bits_succeeded <= _GEN_2398 & _GEN_2335 & _GEN_2240 & _GEN_2177 & (_GEN_1985 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h14 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1920 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h14 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1416 & _GEN_24788 : ~_GEN_219 & _GEN_24788) : casez_tmp_203) : casez_tmp_236);
    ldq_20_bits_order_fail <= _GEN_2398 & _GEN_2335 & _GEN_2240 & _GEN_2177 & (_GEN_757 ? _GEN_93231 : _GEN_759 ? _GEN_760 | _GEN_93231 : _GEN_764 | _GEN_93231);
    ldq_20_bits_observed <= _GEN_757 | (dis_ld_val_3 ? ~_GEN_1416 & _GEN_24852 : ~_GEN_219 & _GEN_24852);
    ldq_20_bits_forward_std_val <= _GEN_2398 & _GEN_2335 & _GEN_2240 & _GEN_2177 & (~_GEN_1183 & _GEN_1953 | ~_GEN_1179 & _GEN_1888 | (dis_ld_val_3 ? ~_GEN_1416 & _GEN_24884 : ~_GEN_219 & _GEN_24884));
    if (_GEN_1985) begin
      if (_GEN_1920) begin
      end
      else
        ldq_20_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_20_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_21_valid <= ~_GEN_1234 & _GEN_2399 & _GEN_2336 & _GEN_2241 & (_GEN_2156 ? ~_GEN_2050 & _GEN_49621 : ~_GEN_2113 & _GEN_49621);
    if (_GEN_318) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_21_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_21_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_21_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_21_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_21_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_220) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_21_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_21_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_21_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_21_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_153) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_21_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_21_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_21_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_55) begin
      ldq_21_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_21_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_21_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_21_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_21_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_21_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_21_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_21_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_21_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_21_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_21_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_21_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_21_bits_st_dep_mask <= next_live_store_mask;
      ldq_21_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_21_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_21_bits_st_dep_mask;
    if (ldq_21_valid)
      ldq_21_bits_uop_br_mask <= ldq_21_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_318)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_220)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_153)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_55)
      ldq_21_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1670) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_21_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_21_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_21_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_21_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_21_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_21_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_21_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_21_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_21_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_21_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_21_bits_addr_bits <= hella_req_addr;
        else
          ldq_21_bits_addr_bits <= 40'h0;
      end
      else
        ldq_21_bits_addr_bits <= _GEN_338;
      ldq_21_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_21_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1574) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_21_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_21_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_21_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_21_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_21_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_21_bits_addr_bits <= _GEN_332;
        else
          ldq_21_bits_addr_bits <= 40'h0;
      end
      else
        ldq_21_bits_addr_bits <= _GEN_334;
      ldq_21_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_21_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_318)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_220)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_153)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_55)
      ldq_21_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_21_bits_addr_valid <= ~_GEN_1234 & _GEN_2399 & _GEN_2336 & _GEN_2241 & (_GEN_2156 ? ~_GEN_2050 & _GEN_81739 : ~_GEN_2113 & _GEN_81739);
    ldq_21_bits_executed <= ~_GEN_1234 & _GEN_2399 & _GEN_2336 & _GEN_2241 & _GEN_2178 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_774) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116716)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1793 & _GEN_113762 : _GEN_1176 ? ~_GEN_1793 & _GEN_113762 : ~(_GEN_113869 & _GEN_1793) & _GEN_113762) : _GEN_113762) | (dis_ld_val_3 ? ~_GEN_1417 & _GEN_24757 : ~_GEN_220 & _GEN_24757));
    ldq_21_bits_succeeded <= _GEN_2399 & _GEN_2336 & _GEN_2241 & _GEN_2178 & (_GEN_1986 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h15 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1921 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h15 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1417 & _GEN_24789 : ~_GEN_220 & _GEN_24789) : casez_tmp_203) : casez_tmp_236);
    ldq_21_bits_order_fail <= _GEN_2399 & _GEN_2336 & _GEN_2241 & _GEN_2178 & (_GEN_777 ? _GEN_93729 : _GEN_779 ? _GEN_780 | _GEN_93729 : _GEN_784 | _GEN_93729);
    ldq_21_bits_observed <= _GEN_777 | (dis_ld_val_3 ? ~_GEN_1417 & _GEN_24853 : ~_GEN_220 & _GEN_24853);
    ldq_21_bits_forward_std_val <= _GEN_2399 & _GEN_2336 & _GEN_2241 & _GEN_2178 & (~_GEN_1183 & _GEN_1954 | ~_GEN_1179 & _GEN_1889 | (dis_ld_val_3 ? ~_GEN_1417 & _GEN_24885 : ~_GEN_220 & _GEN_24885));
    if (_GEN_1986) begin
      if (_GEN_1921) begin
      end
      else
        ldq_21_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_21_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_22_valid <= ~_GEN_1234 & _GEN_2400 & _GEN_2337 & _GEN_2242 & (_GEN_2156 ? ~_GEN_2051 & _GEN_49622 : ~_GEN_2114 & _GEN_49622);
    if (_GEN_319) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_22_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_22_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_22_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_22_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_22_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_221) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_22_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_22_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_22_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_22_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_154) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_22_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_22_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_22_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_56) begin
      ldq_22_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_22_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_22_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_22_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_22_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_22_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_22_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_22_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_22_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_22_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_22_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_22_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_22_bits_st_dep_mask <= next_live_store_mask;
      ldq_22_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_22_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_22_bits_st_dep_mask;
    if (ldq_22_valid)
      ldq_22_bits_uop_br_mask <= ldq_22_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_319)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_221)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_154)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_56)
      ldq_22_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1671) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_22_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_22_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_22_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_22_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_22_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_22_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_22_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_22_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_22_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_22_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_22_bits_addr_bits <= hella_req_addr;
        else
          ldq_22_bits_addr_bits <= 40'h0;
      end
      else
        ldq_22_bits_addr_bits <= _GEN_338;
      ldq_22_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_22_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1575) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_22_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_22_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_22_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_22_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_22_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_22_bits_addr_bits <= _GEN_332;
        else
          ldq_22_bits_addr_bits <= 40'h0;
      end
      else
        ldq_22_bits_addr_bits <= _GEN_334;
      ldq_22_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_22_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_319)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_221)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_154)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_56)
      ldq_22_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_22_bits_addr_valid <= ~_GEN_1234 & _GEN_2400 & _GEN_2337 & _GEN_2242 & (_GEN_2156 ? ~_GEN_2051 & _GEN_81740 : ~_GEN_2114 & _GEN_81740);
    ldq_22_bits_executed <= ~_GEN_1234 & _GEN_2400 & _GEN_2337 & _GEN_2242 & _GEN_2179 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_794) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116717)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1794 & _GEN_113763 : _GEN_1176 ? ~_GEN_1794 & _GEN_113763 : ~(_GEN_113869 & _GEN_1794) & _GEN_113763) : _GEN_113763) | (dis_ld_val_3 ? ~_GEN_1418 & _GEN_24758 : ~_GEN_221 & _GEN_24758));
    ldq_22_bits_succeeded <= _GEN_2400 & _GEN_2337 & _GEN_2242 & _GEN_2179 & (_GEN_1987 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h16 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1922 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h16 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1418 & _GEN_24790 : ~_GEN_221 & _GEN_24790) : casez_tmp_203) : casez_tmp_236);
    ldq_22_bits_order_fail <= _GEN_2400 & _GEN_2337 & _GEN_2242 & _GEN_2179 & (_GEN_797 ? _GEN_94227 : _GEN_799 ? _GEN_800 | _GEN_94227 : _GEN_804 | _GEN_94227);
    ldq_22_bits_observed <= _GEN_797 | (dis_ld_val_3 ? ~_GEN_1418 & _GEN_24854 : ~_GEN_221 & _GEN_24854);
    ldq_22_bits_forward_std_val <= _GEN_2400 & _GEN_2337 & _GEN_2242 & _GEN_2179 & (~_GEN_1183 & _GEN_1955 | ~_GEN_1179 & _GEN_1890 | (dis_ld_val_3 ? ~_GEN_1418 & _GEN_24886 : ~_GEN_221 & _GEN_24886));
    if (_GEN_1987) begin
      if (_GEN_1922) begin
      end
      else
        ldq_22_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_22_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_23_valid <= ~_GEN_1234 & _GEN_2401 & _GEN_2338 & _GEN_2243 & (_GEN_2156 ? ~_GEN_2052 & _GEN_49623 : ~_GEN_2115 & _GEN_49623);
    if (_GEN_320) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_23_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_23_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_23_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_23_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_23_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_222) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_23_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_23_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_23_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_23_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_155) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_23_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_23_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_23_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_57) begin
      ldq_23_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_23_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_23_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_23_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_23_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_23_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_23_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_23_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_23_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_23_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_23_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_23_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_23_bits_st_dep_mask <= next_live_store_mask;
      ldq_23_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_23_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_23_bits_st_dep_mask;
    if (ldq_23_valid)
      ldq_23_bits_uop_br_mask <= ldq_23_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_320)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_222)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_155)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_57)
      ldq_23_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1672) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_23_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_23_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_23_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_23_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_23_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_23_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_23_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_23_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_23_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_23_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_23_bits_addr_bits <= hella_req_addr;
        else
          ldq_23_bits_addr_bits <= 40'h0;
      end
      else
        ldq_23_bits_addr_bits <= _GEN_338;
      ldq_23_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_23_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1576) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_23_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_23_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_23_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_23_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_23_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_23_bits_addr_bits <= _GEN_332;
        else
          ldq_23_bits_addr_bits <= 40'h0;
      end
      else
        ldq_23_bits_addr_bits <= _GEN_334;
      ldq_23_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_23_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_320)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_222)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_155)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_57)
      ldq_23_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_23_bits_addr_valid <= ~_GEN_1234 & _GEN_2401 & _GEN_2338 & _GEN_2243 & (_GEN_2156 ? ~_GEN_2052 & _GEN_81741 : ~_GEN_2115 & _GEN_81741);
    ldq_23_bits_executed <= ~_GEN_1234 & _GEN_2401 & _GEN_2338 & _GEN_2243 & _GEN_2180 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_814) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116718)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1795 & _GEN_113764 : _GEN_1176 ? ~_GEN_1795 & _GEN_113764 : ~(_GEN_113869 & _GEN_1795) & _GEN_113764) : _GEN_113764) | (dis_ld_val_3 ? ~_GEN_1419 & _GEN_24759 : ~_GEN_222 & _GEN_24759));
    ldq_23_bits_succeeded <= _GEN_2401 & _GEN_2338 & _GEN_2243 & _GEN_2180 & (_GEN_1988 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h17 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1923 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h17 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1419 & _GEN_24791 : ~_GEN_222 & _GEN_24791) : casez_tmp_203) : casez_tmp_236);
    ldq_23_bits_order_fail <= _GEN_2401 & _GEN_2338 & _GEN_2243 & _GEN_2180 & (_GEN_817 ? _GEN_94725 : _GEN_819 ? _GEN_820 | _GEN_94725 : _GEN_824 | _GEN_94725);
    ldq_23_bits_observed <= _GEN_817 | (dis_ld_val_3 ? ~_GEN_1419 & _GEN_24855 : ~_GEN_222 & _GEN_24855);
    ldq_23_bits_forward_std_val <= _GEN_2401 & _GEN_2338 & _GEN_2243 & _GEN_2180 & (~_GEN_1183 & _GEN_1956 | ~_GEN_1179 & _GEN_1891 | (dis_ld_val_3 ? ~_GEN_1419 & _GEN_24887 : ~_GEN_222 & _GEN_24887));
    if (_GEN_1988) begin
      if (_GEN_1923) begin
      end
      else
        ldq_23_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_23_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_24_valid <= ~_GEN_1234 & _GEN_2402 & _GEN_2339 & _GEN_2244 & (_GEN_2156 ? ~_GEN_2053 & _GEN_49624 : ~_GEN_2116 & _GEN_49624);
    if (_GEN_321) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_24_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_24_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_24_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_24_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_24_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_223) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_24_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_24_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_24_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_24_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_156) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_24_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_24_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_24_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_58) begin
      ldq_24_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_24_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_24_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_24_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_24_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_24_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_24_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_24_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_24_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_24_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_24_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_24_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_24_bits_st_dep_mask <= next_live_store_mask;
      ldq_24_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_24_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_24_bits_st_dep_mask;
    if (ldq_24_valid)
      ldq_24_bits_uop_br_mask <= ldq_24_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_321)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_223)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_156)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_58)
      ldq_24_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1673) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_24_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_24_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_24_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_24_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_24_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_24_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_24_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_24_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_24_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_24_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_24_bits_addr_bits <= hella_req_addr;
        else
          ldq_24_bits_addr_bits <= 40'h0;
      end
      else
        ldq_24_bits_addr_bits <= _GEN_338;
      ldq_24_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_24_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1577) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_24_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_24_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_24_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_24_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_24_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_24_bits_addr_bits <= _GEN_332;
        else
          ldq_24_bits_addr_bits <= 40'h0;
      end
      else
        ldq_24_bits_addr_bits <= _GEN_334;
      ldq_24_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_24_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_321)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_223)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_156)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_58)
      ldq_24_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_24_bits_addr_valid <= ~_GEN_1234 & _GEN_2402 & _GEN_2339 & _GEN_2244 & (_GEN_2156 ? ~_GEN_2053 & _GEN_81742 : ~_GEN_2116 & _GEN_81742);
    ldq_24_bits_executed <= ~_GEN_1234 & _GEN_2402 & _GEN_2339 & _GEN_2244 & _GEN_2181 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_834) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116719)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1796 & _GEN_113765 : _GEN_1176 ? ~_GEN_1796 & _GEN_113765 : ~(_GEN_113869 & _GEN_1796) & _GEN_113765) : _GEN_113765) | (dis_ld_val_3 ? ~_GEN_1420 & _GEN_24760 : ~_GEN_223 & _GEN_24760));
    ldq_24_bits_succeeded <= _GEN_2402 & _GEN_2339 & _GEN_2244 & _GEN_2181 & (_GEN_1989 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h18 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1924 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h18 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1420 & _GEN_24792 : ~_GEN_223 & _GEN_24792) : casez_tmp_203) : casez_tmp_236);
    ldq_24_bits_order_fail <= _GEN_2402 & _GEN_2339 & _GEN_2244 & _GEN_2181 & (_GEN_837 ? _GEN_95223 : _GEN_839 ? _GEN_840 | _GEN_95223 : _GEN_844 | _GEN_95223);
    ldq_24_bits_observed <= _GEN_837 | (dis_ld_val_3 ? ~_GEN_1420 & _GEN_24856 : ~_GEN_223 & _GEN_24856);
    ldq_24_bits_forward_std_val <= _GEN_2402 & _GEN_2339 & _GEN_2244 & _GEN_2181 & (~_GEN_1183 & _GEN_1957 | ~_GEN_1179 & _GEN_1892 | (dis_ld_val_3 ? ~_GEN_1420 & _GEN_24888 : ~_GEN_223 & _GEN_24888));
    if (_GEN_1989) begin
      if (_GEN_1924) begin
      end
      else
        ldq_24_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_24_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_25_valid <= ~_GEN_1234 & _GEN_2403 & _GEN_2340 & _GEN_2245 & (_GEN_2156 ? ~_GEN_2054 & _GEN_49625 : ~_GEN_2117 & _GEN_49625);
    if (_GEN_322) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_25_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_25_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_25_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_25_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_25_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_224) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_25_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_25_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_25_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_25_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_157) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_25_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_25_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_25_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_59) begin
      ldq_25_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_25_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_25_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_25_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_25_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_25_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_25_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_25_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_25_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_25_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_25_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_25_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_25_bits_st_dep_mask <= next_live_store_mask;
      ldq_25_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_25_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_25_bits_st_dep_mask;
    if (ldq_25_valid)
      ldq_25_bits_uop_br_mask <= ldq_25_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_322)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_224)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_157)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_59)
      ldq_25_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1674) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_25_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_25_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_25_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_25_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_25_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_25_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_25_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_25_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_25_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_25_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_25_bits_addr_bits <= hella_req_addr;
        else
          ldq_25_bits_addr_bits <= 40'h0;
      end
      else
        ldq_25_bits_addr_bits <= _GEN_338;
      ldq_25_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_25_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1578) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_25_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_25_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_25_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_25_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_25_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_25_bits_addr_bits <= _GEN_332;
        else
          ldq_25_bits_addr_bits <= 40'h0;
      end
      else
        ldq_25_bits_addr_bits <= _GEN_334;
      ldq_25_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_25_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_322)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_224)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_157)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_59)
      ldq_25_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_25_bits_addr_valid <= ~_GEN_1234 & _GEN_2403 & _GEN_2340 & _GEN_2245 & (_GEN_2156 ? ~_GEN_2054 & _GEN_81743 : ~_GEN_2117 & _GEN_81743);
    ldq_25_bits_executed <= ~_GEN_1234 & _GEN_2403 & _GEN_2340 & _GEN_2245 & _GEN_2182 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_854) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116720)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1797 & _GEN_113766 : _GEN_1176 ? ~_GEN_1797 & _GEN_113766 : ~(_GEN_113869 & _GEN_1797) & _GEN_113766) : _GEN_113766) | (dis_ld_val_3 ? ~_GEN_1421 & _GEN_24761 : ~_GEN_224 & _GEN_24761));
    ldq_25_bits_succeeded <= _GEN_2403 & _GEN_2340 & _GEN_2245 & _GEN_2182 & (_GEN_1990 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h19 ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1925 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h19 ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1421 & _GEN_24793 : ~_GEN_224 & _GEN_24793) : casez_tmp_203) : casez_tmp_236);
    ldq_25_bits_order_fail <= _GEN_2403 & _GEN_2340 & _GEN_2245 & _GEN_2182 & (_GEN_857 ? _GEN_95721 : _GEN_859 ? _GEN_860 | _GEN_95721 : _GEN_864 | _GEN_95721);
    ldq_25_bits_observed <= _GEN_857 | (dis_ld_val_3 ? ~_GEN_1421 & _GEN_24857 : ~_GEN_224 & _GEN_24857);
    ldq_25_bits_forward_std_val <= _GEN_2403 & _GEN_2340 & _GEN_2245 & _GEN_2182 & (~_GEN_1183 & _GEN_1958 | ~_GEN_1179 & _GEN_1893 | (dis_ld_val_3 ? ~_GEN_1421 & _GEN_24889 : ~_GEN_224 & _GEN_24889));
    if (_GEN_1990) begin
      if (_GEN_1925) begin
      end
      else
        ldq_25_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_25_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_26_valid <= ~_GEN_1234 & _GEN_2404 & _GEN_2341 & _GEN_2246 & (_GEN_2156 ? ~_GEN_2055 & _GEN_49626 : ~_GEN_2118 & _GEN_49626);
    if (_GEN_323) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_26_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_26_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_26_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_26_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_26_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_225) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_26_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_26_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_26_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_26_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_158) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_26_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_26_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_26_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_60) begin
      ldq_26_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_26_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_26_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_26_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_26_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_26_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_26_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_26_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_26_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_26_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_26_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_26_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_26_bits_st_dep_mask <= next_live_store_mask;
      ldq_26_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_26_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_26_bits_st_dep_mask;
    if (ldq_26_valid)
      ldq_26_bits_uop_br_mask <= ldq_26_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_323)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_225)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_158)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_60)
      ldq_26_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1675) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_26_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_26_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_26_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_26_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_26_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_26_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_26_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_26_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_26_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_26_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_26_bits_addr_bits <= hella_req_addr;
        else
          ldq_26_bits_addr_bits <= 40'h0;
      end
      else
        ldq_26_bits_addr_bits <= _GEN_338;
      ldq_26_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_26_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1579) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_26_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_26_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_26_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_26_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_26_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_26_bits_addr_bits <= _GEN_332;
        else
          ldq_26_bits_addr_bits <= 40'h0;
      end
      else
        ldq_26_bits_addr_bits <= _GEN_334;
      ldq_26_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_26_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_323)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_225)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_158)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_60)
      ldq_26_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_26_bits_addr_valid <= ~_GEN_1234 & _GEN_2404 & _GEN_2341 & _GEN_2246 & (_GEN_2156 ? ~_GEN_2055 & _GEN_81744 : ~_GEN_2118 & _GEN_81744);
    ldq_26_bits_executed <= ~_GEN_1234 & _GEN_2404 & _GEN_2341 & _GEN_2246 & _GEN_2183 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_874) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116721)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1798 & _GEN_113767 : _GEN_1176 ? ~_GEN_1798 & _GEN_113767 : ~(_GEN_113869 & _GEN_1798) & _GEN_113767) : _GEN_113767) | (dis_ld_val_3 ? ~_GEN_1422 & _GEN_24762 : ~_GEN_225 & _GEN_24762));
    ldq_26_bits_succeeded <= _GEN_2404 & _GEN_2341 & _GEN_2246 & _GEN_2183 & (_GEN_1991 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1A ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1926 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1A ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1422 & _GEN_24794 : ~_GEN_225 & _GEN_24794) : casez_tmp_203) : casez_tmp_236);
    ldq_26_bits_order_fail <= _GEN_2404 & _GEN_2341 & _GEN_2246 & _GEN_2183 & (_GEN_877 ? _GEN_96219 : _GEN_879 ? _GEN_880 | _GEN_96219 : _GEN_884 | _GEN_96219);
    ldq_26_bits_observed <= _GEN_877 | (dis_ld_val_3 ? ~_GEN_1422 & _GEN_24858 : ~_GEN_225 & _GEN_24858);
    ldq_26_bits_forward_std_val <= _GEN_2404 & _GEN_2341 & _GEN_2246 & _GEN_2183 & (~_GEN_1183 & _GEN_1959 | ~_GEN_1179 & _GEN_1894 | (dis_ld_val_3 ? ~_GEN_1422 & _GEN_24890 : ~_GEN_225 & _GEN_24890));
    if (_GEN_1991) begin
      if (_GEN_1926) begin
      end
      else
        ldq_26_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_26_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_27_valid <= ~_GEN_1234 & _GEN_2405 & _GEN_2342 & _GEN_2247 & (_GEN_2156 ? ~_GEN_2056 & _GEN_49627 : ~_GEN_2119 & _GEN_49627);
    if (_GEN_324) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_27_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_27_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_27_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_27_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_27_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_226) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_27_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_27_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_27_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_27_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_159) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_27_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_27_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_27_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_61) begin
      ldq_27_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_27_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_27_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_27_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_27_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_27_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_27_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_27_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_27_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_27_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_27_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_27_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_27_bits_st_dep_mask <= next_live_store_mask;
      ldq_27_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_27_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_27_bits_st_dep_mask;
    if (ldq_27_valid)
      ldq_27_bits_uop_br_mask <= ldq_27_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_324)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_226)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_159)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_61)
      ldq_27_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1676) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_27_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_27_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_27_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_27_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_27_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_27_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_27_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_27_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_27_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_27_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_27_bits_addr_bits <= hella_req_addr;
        else
          ldq_27_bits_addr_bits <= 40'h0;
      end
      else
        ldq_27_bits_addr_bits <= _GEN_338;
      ldq_27_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_27_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1580) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_27_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_27_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_27_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_27_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_27_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_27_bits_addr_bits <= _GEN_332;
        else
          ldq_27_bits_addr_bits <= 40'h0;
      end
      else
        ldq_27_bits_addr_bits <= _GEN_334;
      ldq_27_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_27_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_324)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_226)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_159)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_61)
      ldq_27_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_27_bits_addr_valid <= ~_GEN_1234 & _GEN_2405 & _GEN_2342 & _GEN_2247 & (_GEN_2156 ? ~_GEN_2056 & _GEN_81745 : ~_GEN_2119 & _GEN_81745);
    ldq_27_bits_executed <= ~_GEN_1234 & _GEN_2405 & _GEN_2342 & _GEN_2247 & _GEN_2184 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_894) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116722)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1799 & _GEN_113768 : _GEN_1176 ? ~_GEN_1799 & _GEN_113768 : ~(_GEN_113869 & _GEN_1799) & _GEN_113768) : _GEN_113768) | (dis_ld_val_3 ? ~_GEN_1423 & _GEN_24763 : ~_GEN_226 & _GEN_24763));
    ldq_27_bits_succeeded <= _GEN_2405 & _GEN_2342 & _GEN_2247 & _GEN_2184 & (_GEN_1992 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1B ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1927 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1B ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1423 & _GEN_24795 : ~_GEN_226 & _GEN_24795) : casez_tmp_203) : casez_tmp_236);
    ldq_27_bits_order_fail <= _GEN_2405 & _GEN_2342 & _GEN_2247 & _GEN_2184 & (_GEN_897 ? _GEN_96717 : _GEN_899 ? _GEN_900 | _GEN_96717 : _GEN_904 | _GEN_96717);
    ldq_27_bits_observed <= _GEN_897 | (dis_ld_val_3 ? ~_GEN_1423 & _GEN_24859 : ~_GEN_226 & _GEN_24859);
    ldq_27_bits_forward_std_val <= _GEN_2405 & _GEN_2342 & _GEN_2247 & _GEN_2184 & (~_GEN_1183 & _GEN_1960 | ~_GEN_1179 & _GEN_1895 | (dis_ld_val_3 ? ~_GEN_1423 & _GEN_24891 : ~_GEN_226 & _GEN_24891));
    if (_GEN_1992) begin
      if (_GEN_1927) begin
      end
      else
        ldq_27_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_27_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_28_valid <= ~_GEN_1234 & _GEN_2406 & _GEN_2343 & _GEN_2248 & (_GEN_2156 ? ~_GEN_2057 & _GEN_49628 : ~_GEN_2120 & _GEN_49628);
    if (_GEN_325) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_28_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_28_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_28_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_28_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_28_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_227) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_28_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_28_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_28_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_28_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_160) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_28_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_28_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_28_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_62) begin
      ldq_28_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_28_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_28_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_28_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_28_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_28_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_28_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_28_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_28_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_28_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_28_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_28_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_28_bits_st_dep_mask <= next_live_store_mask;
      ldq_28_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_28_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_28_bits_st_dep_mask;
    if (ldq_28_valid)
      ldq_28_bits_uop_br_mask <= ldq_28_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_325)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_227)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_160)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_62)
      ldq_28_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1677) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_28_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_28_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_28_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_28_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_28_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_28_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_28_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_28_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_28_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_28_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_28_bits_addr_bits <= hella_req_addr;
        else
          ldq_28_bits_addr_bits <= 40'h0;
      end
      else
        ldq_28_bits_addr_bits <= _GEN_338;
      ldq_28_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_28_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1581) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_28_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_28_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_28_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_28_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_28_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_28_bits_addr_bits <= _GEN_332;
        else
          ldq_28_bits_addr_bits <= 40'h0;
      end
      else
        ldq_28_bits_addr_bits <= _GEN_334;
      ldq_28_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_28_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_325)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_227)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_160)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_62)
      ldq_28_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_28_bits_addr_valid <= ~_GEN_1234 & _GEN_2406 & _GEN_2343 & _GEN_2248 & (_GEN_2156 ? ~_GEN_2057 & _GEN_81746 : ~_GEN_2120 & _GEN_81746);
    ldq_28_bits_executed <= ~_GEN_1234 & _GEN_2406 & _GEN_2343 & _GEN_2248 & _GEN_2185 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_914) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116723)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1800 & _GEN_113769 : _GEN_1176 ? ~_GEN_1800 & _GEN_113769 : ~(_GEN_113869 & _GEN_1800) & _GEN_113769) : _GEN_113769) | (dis_ld_val_3 ? ~_GEN_1424 & _GEN_24764 : ~_GEN_227 & _GEN_24764));
    ldq_28_bits_succeeded <= _GEN_2406 & _GEN_2343 & _GEN_2248 & _GEN_2185 & (_GEN_1993 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1C ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1928 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1C ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1424 & _GEN_24796 : ~_GEN_227 & _GEN_24796) : casez_tmp_203) : casez_tmp_236);
    ldq_28_bits_order_fail <= _GEN_2406 & _GEN_2343 & _GEN_2248 & _GEN_2185 & (_GEN_917 ? _GEN_97215 : _GEN_919 ? _GEN_920 | _GEN_97215 : _GEN_924 | _GEN_97215);
    ldq_28_bits_observed <= _GEN_917 | (dis_ld_val_3 ? ~_GEN_1424 & _GEN_24860 : ~_GEN_227 & _GEN_24860);
    ldq_28_bits_forward_std_val <= _GEN_2406 & _GEN_2343 & _GEN_2248 & _GEN_2185 & (~_GEN_1183 & _GEN_1961 | ~_GEN_1179 & _GEN_1896 | (dis_ld_val_3 ? ~_GEN_1424 & _GEN_24892 : ~_GEN_227 & _GEN_24892));
    if (_GEN_1993) begin
      if (_GEN_1928) begin
      end
      else
        ldq_28_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_28_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_29_valid <= ~_GEN_1234 & _GEN_2407 & _GEN_2344 & _GEN_2249 & (_GEN_2156 ? ~_GEN_2058 & _GEN_49629 : ~_GEN_2121 & _GEN_49629);
    if (_GEN_326) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_29_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_29_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_29_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_29_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_29_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_228) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_29_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_29_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_29_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_29_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_161) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_29_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_29_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_29_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_63) begin
      ldq_29_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_29_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_29_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_29_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_29_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_29_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_29_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_29_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_29_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_29_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_29_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_29_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_29_bits_st_dep_mask <= next_live_store_mask;
      ldq_29_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_29_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_29_bits_st_dep_mask;
    if (ldq_29_valid)
      ldq_29_bits_uop_br_mask <= ldq_29_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_326)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_228)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_161)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_63)
      ldq_29_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1678) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_29_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_29_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_29_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_29_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_29_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_29_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_29_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_29_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_29_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_29_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_29_bits_addr_bits <= hella_req_addr;
        else
          ldq_29_bits_addr_bits <= 40'h0;
      end
      else
        ldq_29_bits_addr_bits <= _GEN_338;
      ldq_29_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_29_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1582) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_29_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_29_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_29_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_29_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_29_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_29_bits_addr_bits <= _GEN_332;
        else
          ldq_29_bits_addr_bits <= 40'h0;
      end
      else
        ldq_29_bits_addr_bits <= _GEN_334;
      ldq_29_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_29_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_326)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_228)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_161)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_63)
      ldq_29_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_29_bits_addr_valid <= ~_GEN_1234 & _GEN_2407 & _GEN_2344 & _GEN_2249 & (_GEN_2156 ? ~_GEN_2058 & _GEN_81747 : ~_GEN_2121 & _GEN_81747);
    ldq_29_bits_executed <= ~_GEN_1234 & _GEN_2407 & _GEN_2344 & _GEN_2249 & _GEN_2186 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_934) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116724)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1801 & _GEN_113770 : _GEN_1176 ? ~_GEN_1801 & _GEN_113770 : ~(_GEN_113869 & _GEN_1801) & _GEN_113770) : _GEN_113770) | (dis_ld_val_3 ? ~_GEN_1425 & _GEN_24765 : ~_GEN_228 & _GEN_24765));
    ldq_29_bits_succeeded <= _GEN_2407 & _GEN_2344 & _GEN_2249 & _GEN_2186 & (_GEN_1994 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1D ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1929 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1D ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1425 & _GEN_24797 : ~_GEN_228 & _GEN_24797) : casez_tmp_203) : casez_tmp_236);
    ldq_29_bits_order_fail <= _GEN_2407 & _GEN_2344 & _GEN_2249 & _GEN_2186 & (_GEN_937 ? _GEN_97713 : _GEN_939 ? _GEN_940 | _GEN_97713 : _GEN_944 | _GEN_97713);
    ldq_29_bits_observed <= _GEN_937 | (dis_ld_val_3 ? ~_GEN_1425 & _GEN_24861 : ~_GEN_228 & _GEN_24861);
    ldq_29_bits_forward_std_val <= _GEN_2407 & _GEN_2344 & _GEN_2249 & _GEN_2186 & (~_GEN_1183 & _GEN_1962 | ~_GEN_1179 & _GEN_1897 | (dis_ld_val_3 ? ~_GEN_1425 & _GEN_24893 : ~_GEN_228 & _GEN_24893));
    if (_GEN_1994) begin
      if (_GEN_1929) begin
      end
      else
        ldq_29_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_29_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_30_valid <= ~_GEN_1234 & _GEN_2408 & _GEN_2345 & _GEN_2250 & (_GEN_2156 ? ~_GEN_2059 & _GEN_49630 : ~_GEN_2122 & _GEN_49630);
    if (_GEN_327) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_30_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_30_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_30_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_30_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_30_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_229) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_30_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_30_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_30_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_30_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_162) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_30_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_30_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_30_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_64) begin
      ldq_30_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_30_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_30_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_30_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_30_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_30_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_30_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_30_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_30_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_30_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_30_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_30_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_30_bits_st_dep_mask <= next_live_store_mask;
      ldq_30_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_30_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_30_bits_st_dep_mask;
    if (ldq_30_valid)
      ldq_30_bits_uop_br_mask <= ldq_30_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_327)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_229)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_162)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_64)
      ldq_30_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & _GEN_1679) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_30_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_30_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_30_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_30_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_30_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_30_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_30_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_30_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_30_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_30_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_30_bits_addr_bits <= hella_req_addr;
        else
          ldq_30_bits_addr_bits <= 40'h0;
      end
      else
        ldq_30_bits_addr_bits <= _GEN_338;
      ldq_30_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_30_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1583) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_30_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_30_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_30_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_30_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_30_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_30_bits_addr_bits <= _GEN_332;
        else
          ldq_30_bits_addr_bits <= 40'h0;
      end
      else
        ldq_30_bits_addr_bits <= _GEN_334;
      ldq_30_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_30_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_327)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_229)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_162)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_64)
      ldq_30_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_30_bits_addr_valid <= ~_GEN_1234 & _GEN_2408 & _GEN_2345 & _GEN_2250 & (_GEN_2156 ? ~_GEN_2059 & _GEN_81748 : ~_GEN_2122 & _GEN_81748);
    ldq_30_bits_executed <= ~_GEN_1234 & _GEN_2408 & _GEN_2345 & _GEN_2250 & _GEN_2187 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_954) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & _GEN_116725)) & ((_GEN_1174 ? (_GEN_113938 ? ~_GEN_1802 & _GEN_113771 : _GEN_1176 ? ~_GEN_1802 & _GEN_113771 : ~(_GEN_113869 & _GEN_1802) & _GEN_113771) : _GEN_113771) | (dis_ld_val_3 ? ~_GEN_1426 & _GEN_24766 : ~_GEN_229 & _GEN_24766));
    ldq_30_bits_succeeded <= _GEN_2408 & _GEN_2345 & _GEN_2250 & _GEN_2187 & (_GEN_1995 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_ldq_idx == 5'h1E ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1930 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_ldq_idx == 5'h1E ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1426 & _GEN_24798 : ~_GEN_229 & _GEN_24798) : casez_tmp_203) : casez_tmp_236);
    ldq_30_bits_order_fail <= _GEN_2408 & _GEN_2345 & _GEN_2250 & _GEN_2187 & (_GEN_957 ? _GEN_98211 : _GEN_959 ? _GEN_960 | _GEN_98211 : _GEN_964 | _GEN_98211);
    ldq_30_bits_observed <= _GEN_957 | (dis_ld_val_3 ? ~_GEN_1426 & _GEN_24862 : ~_GEN_229 & _GEN_24862);
    ldq_30_bits_forward_std_val <= _GEN_2408 & _GEN_2345 & _GEN_2250 & _GEN_2187 & (~_GEN_1183 & _GEN_1963 | ~_GEN_1179 & _GEN_1898 | (dis_ld_val_3 ? ~_GEN_1426 & _GEN_24894 : ~_GEN_229 & _GEN_24894));
    if (_GEN_1995) begin
      if (_GEN_1930) begin
      end
      else
        ldq_30_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_30_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    ldq_31_valid <= ~_GEN_1234 & _GEN_2409 & _GEN_2346 & _GEN_2251 & (_GEN_2156 ? ~_GEN_2060 & _GEN_49631 : ~_GEN_2123 & _GEN_49631);
    if (_GEN_328) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_3_bits_uopc;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_3_bits_mem_signed;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_3_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_3_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_3_bits_uses_stq;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_3_bits_fp_val;
      ldq_31_bits_st_dep_mask <= _ldq_T_115_bits_st_dep_mask;
      if (dis_st_val_2)
        ldq_31_bits_youngest_stq_idx <= _GEN_166;
      else if (dis_st_val_1)
        ldq_31_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_31_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_31_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_230) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_2_bits_uopc;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_2_bits_mem_signed;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_2_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_2_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_2_bits_uses_stq;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_2_bits_fp_val;
      ldq_31_bits_st_dep_mask <= _ldq_T_75_bits_st_dep_mask;
      if (dis_st_val_1)
        ldq_31_bits_youngest_stq_idx <= _GEN_68;
      else if (dis_st_val)
        ldq_31_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_31_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_163) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_1_bits_uopc;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_1_bits_mem_signed;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_1_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_1_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_1_bits_uses_stq;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_1_bits_fp_val;
      ldq_31_bits_st_dep_mask <= _ldq_T_35_bits_st_dep_mask;
      if (dis_st_val)
        ldq_31_bits_youngest_stq_idx <= _GEN_1;
      else
        ldq_31_bits_youngest_stq_idx <= stq_tail;
    end
    else if (_GEN_65) begin
      ldq_31_bits_uop_uopc <= io_core_dis_uops_0_bits_uopc;
      ldq_31_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
      ldq_31_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
      ldq_31_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
      ldq_31_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
      ldq_31_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
      ldq_31_bits_uop_mem_signed <= io_core_dis_uops_0_bits_mem_signed;
      ldq_31_bits_uop_is_amo <= io_core_dis_uops_0_bits_is_amo;
      ldq_31_bits_uop_uses_ldq <= io_core_dis_uops_0_bits_uses_ldq;
      ldq_31_bits_uop_uses_stq <= io_core_dis_uops_0_bits_uses_stq;
      ldq_31_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
      ldq_31_bits_uop_fp_val <= io_core_dis_uops_0_bits_fp_val;
      ldq_31_bits_st_dep_mask <= next_live_store_mask;
      ldq_31_bits_youngest_stq_idx <= stq_tail;
    end
    else
      ldq_31_bits_st_dep_mask <= (_GEN_1267 | ~_ldq_31_bits_st_dep_mask_T) & ldq_31_bits_st_dep_mask;
    if (ldq_31_valid)
      ldq_31_bits_uop_br_mask <= ldq_31_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (_GEN_328)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
    else if (_GEN_230)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
    else if (_GEN_163)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
    else if (_GEN_65)
      ldq_31_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
    if (_GEN_341 & (&ldq_idx_1)) begin
      if (_exe_tlb_uop_T_9) begin
        if (_GEN_329)
          ldq_31_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_31_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else if (will_fire_load_retry_1)
        ldq_31_bits_uop_pdst <= casez_tmp_71;
      else if (will_fire_sta_retry_1)
        ldq_31_bits_uop_pdst <= casez_tmp_60;
      else
        ldq_31_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            ldq_31_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_31_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          ldq_31_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          ldq_31_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          ldq_31_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          ldq_31_bits_addr_bits <= hella_req_addr;
        else
          ldq_31_bits_addr_bits <= 40'h0;
      end
      else
        ldq_31_bits_addr_bits <= _GEN_338;
      ldq_31_bits_addr_is_virtual <= exe_tlb_miss_1;
      ldq_31_bits_addr_is_uncacheable <= _ldq_T_403_bits_addr_is_uncacheable;
    end
    else if (_GEN_1584) begin
      if (_exe_tlb_uop_T_2) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          ldq_31_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
        else
          ldq_31_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
      end
      else
        ldq_31_bits_uop_pdst <= 7'h0;
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            ldq_31_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            ldq_31_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          ldq_31_bits_addr_bits <= _GEN_332;
        else
          ldq_31_bits_addr_bits <= 40'h0;
      end
      else
        ldq_31_bits_addr_bits <= _GEN_334;
      ldq_31_bits_addr_is_virtual <= exe_tlb_miss_0;
      ldq_31_bits_addr_is_uncacheable <= _ldq_T_340_bits_addr_is_uncacheable;
    end
    else if (_GEN_328)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
    else if (_GEN_230)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
    else if (_GEN_163)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
    else if (_GEN_65)
      ldq_31_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
    ldq_31_bits_addr_valid <= ~_GEN_1234 & _GEN_2409 & _GEN_2346 & _GEN_2251 & (_GEN_2156 ? ~_GEN_2060 & _GEN_81749 : ~_GEN_2123 & _GEN_81749);
    ldq_31_bits_executed <= ~_GEN_1234 & _GEN_2409 & _GEN_2346 & _GEN_2251 & _GEN_2188 & (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | ~_GEN_973) & (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | ~(io_dmem_nack_0_bits_uop_uses_ldq & (&io_dmem_nack_0_bits_uop_ldq_idx))) & ((_GEN_1174 ? (_GEN_113938 ? ~(&lcam_ldq_idx_1) & _GEN_113772 : _GEN_1176 ? ~(&lcam_ldq_idx_1) & _GEN_113772 : ~(_GEN_113869 & (&lcam_ldq_idx_1)) & _GEN_113772) : _GEN_113772) | (dis_ld_val_3 ? ~_GEN_1427 & _GEN_24767 : ~_GEN_230 & _GEN_24767));
    ldq_31_bits_succeeded <= _GEN_2409 & _GEN_2346 & _GEN_2251 & _GEN_2188 & (_GEN_1996 ? (io_dmem_resp_1_valid & io_dmem_resp_1_bits_uop_uses_ldq & (&io_dmem_resp_1_bits_uop_ldq_idx) ? _ldq_io_dmem_resp_1_bits_uop_ldq_idx_bits_succeeded : _GEN_1931 ? (io_dmem_resp_0_valid & io_dmem_resp_0_bits_uop_uses_ldq & (&io_dmem_resp_0_bits_uop_ldq_idx) ? _ldq_io_dmem_resp_0_bits_uop_ldq_idx_bits_succeeded : dis_ld_val_3 ? ~_GEN_1427 & _GEN_24799 : ~_GEN_230 & _GEN_24799) : casez_tmp_203) : casez_tmp_236);
    ldq_31_bits_order_fail <= _GEN_2409 & _GEN_2346 & _GEN_2251 & _GEN_2188 & (_GEN_976 ? _GEN_98709 : _GEN_978 ? _GEN_979 | _GEN_98709 : _GEN_982 | _GEN_98709);
    ldq_31_bits_observed <= _GEN_976 | (dis_ld_val_3 ? ~_GEN_1427 & _GEN_24863 : ~_GEN_230 & _GEN_24863);
    ldq_31_bits_forward_std_val <= _GEN_2409 & _GEN_2346 & _GEN_2251 & _GEN_2188 & (~_GEN_1183 & _GEN_1964 | ~_GEN_1179 & _GEN_1899 | (dis_ld_val_3 ? ~_GEN_1427 & _GEN_24895 : ~_GEN_230 & _GEN_24895));
    if (_GEN_1996) begin
      if (_GEN_1931) begin
      end
      else
        ldq_31_bits_forward_stq_idx <= wb_forward_stq_idx_0;
    end
    else
      ldq_31_bits_forward_stq_idx <= wb_forward_stq_idx_1;
    stq_0_valid <= ~_GEN_2479 & (clear_store ? ~_GEN_2411 & _GEN_52416 : ~_GEN_1997 & _GEN_52416);
    if (_GEN_1235) begin
      stq_0_bits_uop_br_mask <= 20'h0;
      stq_0_bits_uop_rob_idx <= 7'h0;
      stq_0_bits_uop_ldq_idx <= 5'h0;
      stq_0_bits_uop_stq_idx <= 5'h0;
      stq_0_bits_uop_pdst <= 7'h0;
      stq_0_bits_uop_mem_cmd <= 5'h0;
      stq_0_bits_uop_mem_size <= 2'h0;
      stq_0_bits_uop_dst_rtype <= 2'h2;
      stq_1_bits_uop_br_mask <= 20'h0;
      stq_1_bits_uop_rob_idx <= 7'h0;
      stq_1_bits_uop_ldq_idx <= 5'h0;
      stq_1_bits_uop_stq_idx <= 5'h0;
      stq_1_bits_uop_pdst <= 7'h0;
      stq_1_bits_uop_mem_cmd <= 5'h0;
      stq_1_bits_uop_mem_size <= 2'h0;
      stq_1_bits_uop_dst_rtype <= 2'h2;
      stq_2_bits_uop_br_mask <= 20'h0;
      stq_2_bits_uop_rob_idx <= 7'h0;
      stq_2_bits_uop_ldq_idx <= 5'h0;
      stq_2_bits_uop_stq_idx <= 5'h0;
      stq_2_bits_uop_pdst <= 7'h0;
      stq_2_bits_uop_mem_cmd <= 5'h0;
      stq_2_bits_uop_mem_size <= 2'h0;
      stq_2_bits_uop_dst_rtype <= 2'h2;
      stq_3_bits_uop_br_mask <= 20'h0;
      stq_3_bits_uop_rob_idx <= 7'h0;
      stq_3_bits_uop_ldq_idx <= 5'h0;
      stq_3_bits_uop_stq_idx <= 5'h0;
      stq_3_bits_uop_pdst <= 7'h0;
      stq_3_bits_uop_mem_cmd <= 5'h0;
      stq_3_bits_uop_mem_size <= 2'h0;
      stq_3_bits_uop_dst_rtype <= 2'h2;
      stq_4_bits_uop_br_mask <= 20'h0;
      stq_4_bits_uop_rob_idx <= 7'h0;
      stq_4_bits_uop_ldq_idx <= 5'h0;
      stq_4_bits_uop_stq_idx <= 5'h0;
      stq_4_bits_uop_pdst <= 7'h0;
      stq_4_bits_uop_mem_cmd <= 5'h0;
      stq_4_bits_uop_mem_size <= 2'h0;
      stq_4_bits_uop_dst_rtype <= 2'h2;
      stq_5_bits_uop_br_mask <= 20'h0;
      stq_5_bits_uop_rob_idx <= 7'h0;
      stq_5_bits_uop_ldq_idx <= 5'h0;
      stq_5_bits_uop_stq_idx <= 5'h0;
      stq_5_bits_uop_pdst <= 7'h0;
      stq_5_bits_uop_mem_cmd <= 5'h0;
      stq_5_bits_uop_mem_size <= 2'h0;
      stq_5_bits_uop_dst_rtype <= 2'h2;
      stq_6_bits_uop_br_mask <= 20'h0;
      stq_6_bits_uop_rob_idx <= 7'h0;
      stq_6_bits_uop_ldq_idx <= 5'h0;
      stq_6_bits_uop_stq_idx <= 5'h0;
      stq_6_bits_uop_pdst <= 7'h0;
      stq_6_bits_uop_mem_cmd <= 5'h0;
      stq_6_bits_uop_mem_size <= 2'h0;
      stq_6_bits_uop_dst_rtype <= 2'h2;
      stq_7_bits_uop_br_mask <= 20'h0;
      stq_7_bits_uop_rob_idx <= 7'h0;
      stq_7_bits_uop_ldq_idx <= 5'h0;
      stq_7_bits_uop_stq_idx <= 5'h0;
      stq_7_bits_uop_pdst <= 7'h0;
      stq_7_bits_uop_mem_cmd <= 5'h0;
      stq_7_bits_uop_mem_size <= 2'h0;
      stq_7_bits_uop_dst_rtype <= 2'h2;
      stq_8_bits_uop_br_mask <= 20'h0;
      stq_8_bits_uop_rob_idx <= 7'h0;
      stq_8_bits_uop_ldq_idx <= 5'h0;
      stq_8_bits_uop_stq_idx <= 5'h0;
      stq_8_bits_uop_pdst <= 7'h0;
      stq_8_bits_uop_mem_cmd <= 5'h0;
      stq_8_bits_uop_mem_size <= 2'h0;
      stq_8_bits_uop_dst_rtype <= 2'h2;
      stq_9_bits_uop_br_mask <= 20'h0;
      stq_9_bits_uop_rob_idx <= 7'h0;
      stq_9_bits_uop_ldq_idx <= 5'h0;
      stq_9_bits_uop_stq_idx <= 5'h0;
      stq_9_bits_uop_pdst <= 7'h0;
      stq_9_bits_uop_mem_cmd <= 5'h0;
      stq_9_bits_uop_mem_size <= 2'h0;
      stq_9_bits_uop_dst_rtype <= 2'h2;
      stq_10_bits_uop_br_mask <= 20'h0;
      stq_10_bits_uop_rob_idx <= 7'h0;
      stq_10_bits_uop_ldq_idx <= 5'h0;
      stq_10_bits_uop_stq_idx <= 5'h0;
      stq_10_bits_uop_pdst <= 7'h0;
      stq_10_bits_uop_mem_cmd <= 5'h0;
      stq_10_bits_uop_mem_size <= 2'h0;
      stq_10_bits_uop_dst_rtype <= 2'h2;
      stq_11_bits_uop_br_mask <= 20'h0;
      stq_11_bits_uop_rob_idx <= 7'h0;
      stq_11_bits_uop_ldq_idx <= 5'h0;
      stq_11_bits_uop_stq_idx <= 5'h0;
      stq_11_bits_uop_pdst <= 7'h0;
      stq_11_bits_uop_mem_cmd <= 5'h0;
      stq_11_bits_uop_mem_size <= 2'h0;
      stq_11_bits_uop_dst_rtype <= 2'h2;
      stq_12_bits_uop_br_mask <= 20'h0;
      stq_12_bits_uop_rob_idx <= 7'h0;
      stq_12_bits_uop_ldq_idx <= 5'h0;
      stq_12_bits_uop_stq_idx <= 5'h0;
      stq_12_bits_uop_pdst <= 7'h0;
      stq_12_bits_uop_mem_cmd <= 5'h0;
      stq_12_bits_uop_mem_size <= 2'h0;
      stq_12_bits_uop_dst_rtype <= 2'h2;
      stq_13_bits_uop_br_mask <= 20'h0;
      stq_13_bits_uop_rob_idx <= 7'h0;
      stq_13_bits_uop_ldq_idx <= 5'h0;
      stq_13_bits_uop_stq_idx <= 5'h0;
      stq_13_bits_uop_pdst <= 7'h0;
      stq_13_bits_uop_mem_cmd <= 5'h0;
      stq_13_bits_uop_mem_size <= 2'h0;
      stq_13_bits_uop_dst_rtype <= 2'h2;
      stq_14_bits_uop_br_mask <= 20'h0;
      stq_14_bits_uop_rob_idx <= 7'h0;
      stq_14_bits_uop_ldq_idx <= 5'h0;
      stq_14_bits_uop_stq_idx <= 5'h0;
      stq_14_bits_uop_pdst <= 7'h0;
      stq_14_bits_uop_mem_cmd <= 5'h0;
      stq_14_bits_uop_mem_size <= 2'h0;
      stq_14_bits_uop_dst_rtype <= 2'h2;
      stq_15_bits_uop_br_mask <= 20'h0;
      stq_15_bits_uop_rob_idx <= 7'h0;
      stq_15_bits_uop_ldq_idx <= 5'h0;
      stq_15_bits_uop_stq_idx <= 5'h0;
      stq_15_bits_uop_pdst <= 7'h0;
      stq_15_bits_uop_mem_cmd <= 5'h0;
      stq_15_bits_uop_mem_size <= 2'h0;
      stq_15_bits_uop_dst_rtype <= 2'h2;
      stq_16_bits_uop_br_mask <= 20'h0;
      stq_16_bits_uop_rob_idx <= 7'h0;
      stq_16_bits_uop_ldq_idx <= 5'h0;
      stq_16_bits_uop_stq_idx <= 5'h0;
      stq_16_bits_uop_pdst <= 7'h0;
      stq_16_bits_uop_mem_cmd <= 5'h0;
      stq_16_bits_uop_mem_size <= 2'h0;
      stq_16_bits_uop_dst_rtype <= 2'h2;
      stq_17_bits_uop_br_mask <= 20'h0;
      stq_17_bits_uop_rob_idx <= 7'h0;
      stq_17_bits_uop_ldq_idx <= 5'h0;
      stq_17_bits_uop_stq_idx <= 5'h0;
      stq_17_bits_uop_pdst <= 7'h0;
      stq_17_bits_uop_mem_cmd <= 5'h0;
      stq_17_bits_uop_mem_size <= 2'h0;
      stq_17_bits_uop_dst_rtype <= 2'h2;
      stq_18_bits_uop_br_mask <= 20'h0;
      stq_18_bits_uop_rob_idx <= 7'h0;
      stq_18_bits_uop_ldq_idx <= 5'h0;
      stq_18_bits_uop_stq_idx <= 5'h0;
      stq_18_bits_uop_pdst <= 7'h0;
      stq_18_bits_uop_mem_cmd <= 5'h0;
      stq_18_bits_uop_mem_size <= 2'h0;
      stq_18_bits_uop_dst_rtype <= 2'h2;
      stq_19_bits_uop_br_mask <= 20'h0;
      stq_19_bits_uop_rob_idx <= 7'h0;
      stq_19_bits_uop_ldq_idx <= 5'h0;
      stq_19_bits_uop_stq_idx <= 5'h0;
      stq_19_bits_uop_pdst <= 7'h0;
      stq_19_bits_uop_mem_cmd <= 5'h0;
      stq_19_bits_uop_mem_size <= 2'h0;
      stq_19_bits_uop_dst_rtype <= 2'h2;
      stq_20_bits_uop_br_mask <= 20'h0;
      stq_20_bits_uop_rob_idx <= 7'h0;
      stq_20_bits_uop_ldq_idx <= 5'h0;
      stq_20_bits_uop_stq_idx <= 5'h0;
      stq_20_bits_uop_pdst <= 7'h0;
      stq_20_bits_uop_mem_cmd <= 5'h0;
      stq_20_bits_uop_mem_size <= 2'h0;
      stq_20_bits_uop_dst_rtype <= 2'h2;
      stq_21_bits_uop_br_mask <= 20'h0;
      stq_21_bits_uop_rob_idx <= 7'h0;
      stq_21_bits_uop_ldq_idx <= 5'h0;
      stq_21_bits_uop_stq_idx <= 5'h0;
      stq_21_bits_uop_pdst <= 7'h0;
      stq_21_bits_uop_mem_cmd <= 5'h0;
      stq_21_bits_uop_mem_size <= 2'h0;
      stq_21_bits_uop_dst_rtype <= 2'h2;
      stq_22_bits_uop_br_mask <= 20'h0;
      stq_22_bits_uop_rob_idx <= 7'h0;
      stq_22_bits_uop_ldq_idx <= 5'h0;
      stq_22_bits_uop_stq_idx <= 5'h0;
      stq_22_bits_uop_pdst <= 7'h0;
      stq_22_bits_uop_mem_cmd <= 5'h0;
      stq_22_bits_uop_mem_size <= 2'h0;
      stq_22_bits_uop_dst_rtype <= 2'h2;
      stq_23_bits_uop_br_mask <= 20'h0;
      stq_23_bits_uop_rob_idx <= 7'h0;
      stq_23_bits_uop_ldq_idx <= 5'h0;
      stq_23_bits_uop_stq_idx <= 5'h0;
      stq_23_bits_uop_pdst <= 7'h0;
      stq_23_bits_uop_mem_cmd <= 5'h0;
      stq_23_bits_uop_mem_size <= 2'h0;
      stq_23_bits_uop_dst_rtype <= 2'h2;
      stq_24_bits_uop_br_mask <= 20'h0;
      stq_24_bits_uop_rob_idx <= 7'h0;
      stq_24_bits_uop_ldq_idx <= 5'h0;
      stq_24_bits_uop_stq_idx <= 5'h0;
      stq_24_bits_uop_pdst <= 7'h0;
      stq_24_bits_uop_mem_cmd <= 5'h0;
      stq_24_bits_uop_mem_size <= 2'h0;
      stq_24_bits_uop_dst_rtype <= 2'h2;
      stq_25_bits_uop_br_mask <= 20'h0;
      stq_25_bits_uop_rob_idx <= 7'h0;
      stq_25_bits_uop_ldq_idx <= 5'h0;
      stq_25_bits_uop_stq_idx <= 5'h0;
      stq_25_bits_uop_pdst <= 7'h0;
      stq_25_bits_uop_mem_cmd <= 5'h0;
      stq_25_bits_uop_mem_size <= 2'h0;
      stq_25_bits_uop_dst_rtype <= 2'h2;
      stq_26_bits_uop_br_mask <= 20'h0;
      stq_26_bits_uop_rob_idx <= 7'h0;
      stq_26_bits_uop_ldq_idx <= 5'h0;
      stq_26_bits_uop_stq_idx <= 5'h0;
      stq_26_bits_uop_pdst <= 7'h0;
      stq_26_bits_uop_mem_cmd <= 5'h0;
      stq_26_bits_uop_mem_size <= 2'h0;
      stq_26_bits_uop_dst_rtype <= 2'h2;
      stq_27_bits_uop_br_mask <= 20'h0;
      stq_27_bits_uop_rob_idx <= 7'h0;
      stq_27_bits_uop_ldq_idx <= 5'h0;
      stq_27_bits_uop_stq_idx <= 5'h0;
      stq_27_bits_uop_pdst <= 7'h0;
      stq_27_bits_uop_mem_cmd <= 5'h0;
      stq_27_bits_uop_mem_size <= 2'h0;
      stq_27_bits_uop_dst_rtype <= 2'h2;
      stq_28_bits_uop_br_mask <= 20'h0;
      stq_28_bits_uop_rob_idx <= 7'h0;
      stq_28_bits_uop_ldq_idx <= 5'h0;
      stq_28_bits_uop_stq_idx <= 5'h0;
      stq_28_bits_uop_pdst <= 7'h0;
      stq_28_bits_uop_mem_cmd <= 5'h0;
      stq_28_bits_uop_mem_size <= 2'h0;
      stq_28_bits_uop_dst_rtype <= 2'h2;
      stq_29_bits_uop_br_mask <= 20'h0;
      stq_29_bits_uop_rob_idx <= 7'h0;
      stq_29_bits_uop_ldq_idx <= 5'h0;
      stq_29_bits_uop_stq_idx <= 5'h0;
      stq_29_bits_uop_pdst <= 7'h0;
      stq_29_bits_uop_mem_cmd <= 5'h0;
      stq_29_bits_uop_mem_size <= 2'h0;
      stq_29_bits_uop_dst_rtype <= 2'h2;
      stq_30_bits_uop_br_mask <= 20'h0;
      stq_30_bits_uop_rob_idx <= 7'h0;
      stq_30_bits_uop_ldq_idx <= 5'h0;
      stq_30_bits_uop_stq_idx <= 5'h0;
      stq_30_bits_uop_pdst <= 7'h0;
      stq_30_bits_uop_mem_cmd <= 5'h0;
      stq_30_bits_uop_mem_size <= 2'h0;
      stq_30_bits_uop_dst_rtype <= 2'h2;
      stq_31_bits_uop_br_mask <= 20'h0;
      stq_31_bits_uop_rob_idx <= 7'h0;
      stq_31_bits_uop_ldq_idx <= 5'h0;
      stq_31_bits_uop_stq_idx <= 5'h0;
      stq_31_bits_uop_pdst <= 7'h0;
      stq_31_bits_uop_mem_cmd <= 5'h0;
      stq_31_bits_uop_mem_size <= 2'h0;
      stq_31_bits_uop_dst_rtype <= 2'h2;
      stq_head <= 5'h0;
      stq_commit_head <= 5'h0;
      stq_execute_head <= 5'h0;
    end
    else begin
      if (stq_0_valid)
        stq_0_bits_uop_br_mask <= stq_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1428) begin
        if (_GEN_1364) begin
          if (_GEN_1332) begin
            if (_GEN_1268) begin
            end
            else
              stq_0_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_0_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_0_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_0_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1428) begin
        if (_GEN_1364) begin
          if (_GEN_1332) begin
            if (_GEN_1268) begin
            end
            else begin
              stq_0_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_0_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_0_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_0_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_0_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_0_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_0_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_0_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_0_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_0_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_0_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_0_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1680) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_0_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_0_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_0_bits_uop_pdst <= casez_tmp_60;
        else
          stq_0_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1585) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_0_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_0_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_0_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1428) begin
        if (_GEN_1364) begin
          if (_GEN_1332) begin
            if (_GEN_1268) begin
            end
            else
              stq_0_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_0_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_0_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_0_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1428) begin
        if (_GEN_1364) begin
          if (_GEN_1332) begin
            if (_GEN_1268) begin
            end
            else begin
              stq_0_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_0_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_0_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_0_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_0_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_0_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_0_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_0_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_0_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_0_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_0_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_0_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_1_valid)
        stq_1_bits_uop_br_mask <= stq_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1429) begin
        if (_GEN_1365) begin
          if (_GEN_1333) begin
            if (_GEN_1269) begin
            end
            else
              stq_1_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_1_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_1_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_1_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1429) begin
        if (_GEN_1365) begin
          if (_GEN_1333) begin
            if (_GEN_1269) begin
            end
            else begin
              stq_1_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_1_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_1_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_1_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_1_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_1_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_1_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_1_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_1_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_1_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_1_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_1_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1681) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_1_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_1_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_1_bits_uop_pdst <= casez_tmp_60;
        else
          stq_1_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1586) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_1_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_1_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_1_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1429) begin
        if (_GEN_1365) begin
          if (_GEN_1333) begin
            if (_GEN_1269) begin
            end
            else
              stq_1_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_1_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_1_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_1_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1429) begin
        if (_GEN_1365) begin
          if (_GEN_1333) begin
            if (_GEN_1269) begin
            end
            else begin
              stq_1_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_1_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_1_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_1_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_1_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_1_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_1_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_1_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_1_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_1_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_1_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_1_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_2_valid)
        stq_2_bits_uop_br_mask <= stq_2_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1430) begin
        if (_GEN_1366) begin
          if (_GEN_1334) begin
            if (_GEN_1270) begin
            end
            else
              stq_2_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_2_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_2_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_2_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1430) begin
        if (_GEN_1366) begin
          if (_GEN_1334) begin
            if (_GEN_1270) begin
            end
            else begin
              stq_2_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_2_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_2_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_2_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_2_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_2_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_2_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_2_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_2_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_2_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_2_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_2_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1682) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_2_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_2_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_2_bits_uop_pdst <= casez_tmp_60;
        else
          stq_2_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1587) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_2_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_2_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_2_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1430) begin
        if (_GEN_1366) begin
          if (_GEN_1334) begin
            if (_GEN_1270) begin
            end
            else
              stq_2_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_2_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_2_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_2_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1430) begin
        if (_GEN_1366) begin
          if (_GEN_1334) begin
            if (_GEN_1270) begin
            end
            else begin
              stq_2_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_2_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_2_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_2_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_2_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_2_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_2_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_2_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_2_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_2_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_2_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_2_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_3_valid)
        stq_3_bits_uop_br_mask <= stq_3_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1431) begin
        if (_GEN_1367) begin
          if (_GEN_1335) begin
            if (_GEN_1271) begin
            end
            else
              stq_3_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_3_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_3_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_3_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1431) begin
        if (_GEN_1367) begin
          if (_GEN_1335) begin
            if (_GEN_1271) begin
            end
            else begin
              stq_3_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_3_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_3_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_3_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_3_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_3_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_3_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_3_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_3_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_3_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_3_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_3_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1683) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_3_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_3_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_3_bits_uop_pdst <= casez_tmp_60;
        else
          stq_3_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1588) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_3_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_3_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_3_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1431) begin
        if (_GEN_1367) begin
          if (_GEN_1335) begin
            if (_GEN_1271) begin
            end
            else
              stq_3_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_3_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_3_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_3_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1431) begin
        if (_GEN_1367) begin
          if (_GEN_1335) begin
            if (_GEN_1271) begin
            end
            else begin
              stq_3_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_3_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_3_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_3_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_3_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_3_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_3_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_3_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_3_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_3_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_3_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_3_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_4_valid)
        stq_4_bits_uop_br_mask <= stq_4_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1432) begin
        if (_GEN_1368) begin
          if (_GEN_1336) begin
            if (_GEN_1272) begin
            end
            else
              stq_4_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_4_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_4_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_4_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1432) begin
        if (_GEN_1368) begin
          if (_GEN_1336) begin
            if (_GEN_1272) begin
            end
            else begin
              stq_4_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_4_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_4_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_4_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_4_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_4_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_4_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_4_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_4_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_4_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_4_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_4_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1684) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_4_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_4_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_4_bits_uop_pdst <= casez_tmp_60;
        else
          stq_4_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1589) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_4_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_4_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_4_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1432) begin
        if (_GEN_1368) begin
          if (_GEN_1336) begin
            if (_GEN_1272) begin
            end
            else
              stq_4_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_4_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_4_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_4_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1432) begin
        if (_GEN_1368) begin
          if (_GEN_1336) begin
            if (_GEN_1272) begin
            end
            else begin
              stq_4_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_4_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_4_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_4_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_4_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_4_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_4_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_4_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_4_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_4_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_4_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_4_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_5_valid)
        stq_5_bits_uop_br_mask <= stq_5_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1433) begin
        if (_GEN_1369) begin
          if (_GEN_1337) begin
            if (_GEN_1273) begin
            end
            else
              stq_5_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_5_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_5_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_5_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1433) begin
        if (_GEN_1369) begin
          if (_GEN_1337) begin
            if (_GEN_1273) begin
            end
            else begin
              stq_5_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_5_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_5_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_5_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_5_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_5_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_5_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_5_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_5_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_5_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_5_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_5_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1685) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_5_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_5_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_5_bits_uop_pdst <= casez_tmp_60;
        else
          stq_5_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1590) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_5_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_5_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_5_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1433) begin
        if (_GEN_1369) begin
          if (_GEN_1337) begin
            if (_GEN_1273) begin
            end
            else
              stq_5_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_5_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_5_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_5_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1433) begin
        if (_GEN_1369) begin
          if (_GEN_1337) begin
            if (_GEN_1273) begin
            end
            else begin
              stq_5_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_5_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_5_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_5_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_5_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_5_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_5_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_5_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_5_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_5_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_5_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_5_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_6_valid)
        stq_6_bits_uop_br_mask <= stq_6_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1434) begin
        if (_GEN_1370) begin
          if (_GEN_1338) begin
            if (_GEN_1274) begin
            end
            else
              stq_6_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_6_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_6_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_6_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1434) begin
        if (_GEN_1370) begin
          if (_GEN_1338) begin
            if (_GEN_1274) begin
            end
            else begin
              stq_6_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_6_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_6_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_6_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_6_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_6_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_6_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_6_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_6_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_6_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_6_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_6_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1686) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_6_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_6_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_6_bits_uop_pdst <= casez_tmp_60;
        else
          stq_6_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1591) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_6_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_6_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_6_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1434) begin
        if (_GEN_1370) begin
          if (_GEN_1338) begin
            if (_GEN_1274) begin
            end
            else
              stq_6_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_6_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_6_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_6_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1434) begin
        if (_GEN_1370) begin
          if (_GEN_1338) begin
            if (_GEN_1274) begin
            end
            else begin
              stq_6_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_6_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_6_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_6_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_6_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_6_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_6_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_6_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_6_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_6_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_6_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_6_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_7_valid)
        stq_7_bits_uop_br_mask <= stq_7_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1435) begin
        if (_GEN_1371) begin
          if (_GEN_1339) begin
            if (_GEN_1275) begin
            end
            else
              stq_7_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_7_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_7_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_7_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1435) begin
        if (_GEN_1371) begin
          if (_GEN_1339) begin
            if (_GEN_1275) begin
            end
            else begin
              stq_7_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_7_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_7_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_7_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_7_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_7_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_7_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_7_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_7_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_7_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_7_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_7_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1687) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_7_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_7_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_7_bits_uop_pdst <= casez_tmp_60;
        else
          stq_7_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1592) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_7_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_7_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_7_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1435) begin
        if (_GEN_1371) begin
          if (_GEN_1339) begin
            if (_GEN_1275) begin
            end
            else
              stq_7_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_7_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_7_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_7_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1435) begin
        if (_GEN_1371) begin
          if (_GEN_1339) begin
            if (_GEN_1275) begin
            end
            else begin
              stq_7_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_7_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_7_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_7_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_7_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_7_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_7_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_7_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_7_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_7_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_7_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_7_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_8_valid)
        stq_8_bits_uop_br_mask <= stq_8_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1436) begin
        if (_GEN_1372) begin
          if (_GEN_1340) begin
            if (_GEN_1276) begin
            end
            else
              stq_8_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_8_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_8_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_8_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1436) begin
        if (_GEN_1372) begin
          if (_GEN_1340) begin
            if (_GEN_1276) begin
            end
            else begin
              stq_8_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_8_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_8_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_8_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_8_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_8_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_8_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_8_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_8_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_8_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_8_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_8_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1688) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_8_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_8_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_8_bits_uop_pdst <= casez_tmp_60;
        else
          stq_8_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1593) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_8_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_8_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_8_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1436) begin
        if (_GEN_1372) begin
          if (_GEN_1340) begin
            if (_GEN_1276) begin
            end
            else
              stq_8_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_8_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_8_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_8_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1436) begin
        if (_GEN_1372) begin
          if (_GEN_1340) begin
            if (_GEN_1276) begin
            end
            else begin
              stq_8_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_8_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_8_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_8_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_8_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_8_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_8_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_8_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_8_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_8_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_8_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_8_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_9_valid)
        stq_9_bits_uop_br_mask <= stq_9_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1437) begin
        if (_GEN_1373) begin
          if (_GEN_1341) begin
            if (_GEN_1277) begin
            end
            else
              stq_9_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_9_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_9_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_9_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1437) begin
        if (_GEN_1373) begin
          if (_GEN_1341) begin
            if (_GEN_1277) begin
            end
            else begin
              stq_9_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_9_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_9_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_9_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_9_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_9_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_9_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_9_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_9_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_9_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_9_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_9_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1689) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_9_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_9_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_9_bits_uop_pdst <= casez_tmp_60;
        else
          stq_9_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1594) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_9_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_9_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_9_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1437) begin
        if (_GEN_1373) begin
          if (_GEN_1341) begin
            if (_GEN_1277) begin
            end
            else
              stq_9_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_9_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_9_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_9_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1437) begin
        if (_GEN_1373) begin
          if (_GEN_1341) begin
            if (_GEN_1277) begin
            end
            else begin
              stq_9_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_9_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_9_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_9_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_9_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_9_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_9_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_9_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_9_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_9_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_9_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_9_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_10_valid)
        stq_10_bits_uop_br_mask <= stq_10_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1438) begin
        if (_GEN_1374) begin
          if (_GEN_1342) begin
            if (_GEN_1278) begin
            end
            else
              stq_10_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_10_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_10_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_10_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1438) begin
        if (_GEN_1374) begin
          if (_GEN_1342) begin
            if (_GEN_1278) begin
            end
            else begin
              stq_10_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_10_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_10_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_10_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_10_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_10_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_10_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_10_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_10_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_10_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_10_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_10_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1690) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_10_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_10_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_10_bits_uop_pdst <= casez_tmp_60;
        else
          stq_10_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1595) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_10_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_10_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_10_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1438) begin
        if (_GEN_1374) begin
          if (_GEN_1342) begin
            if (_GEN_1278) begin
            end
            else
              stq_10_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_10_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_10_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_10_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1438) begin
        if (_GEN_1374) begin
          if (_GEN_1342) begin
            if (_GEN_1278) begin
            end
            else begin
              stq_10_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_10_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_10_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_10_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_10_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_10_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_10_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_10_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_10_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_10_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_10_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_10_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_11_valid)
        stq_11_bits_uop_br_mask <= stq_11_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1439) begin
        if (_GEN_1375) begin
          if (_GEN_1343) begin
            if (_GEN_1279) begin
            end
            else
              stq_11_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_11_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_11_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_11_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1439) begin
        if (_GEN_1375) begin
          if (_GEN_1343) begin
            if (_GEN_1279) begin
            end
            else begin
              stq_11_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_11_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_11_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_11_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_11_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_11_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_11_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_11_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_11_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_11_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_11_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_11_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1691) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_11_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_11_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_11_bits_uop_pdst <= casez_tmp_60;
        else
          stq_11_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1596) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_11_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_11_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_11_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1439) begin
        if (_GEN_1375) begin
          if (_GEN_1343) begin
            if (_GEN_1279) begin
            end
            else
              stq_11_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_11_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_11_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_11_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1439) begin
        if (_GEN_1375) begin
          if (_GEN_1343) begin
            if (_GEN_1279) begin
            end
            else begin
              stq_11_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_11_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_11_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_11_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_11_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_11_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_11_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_11_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_11_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_11_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_11_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_11_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_12_valid)
        stq_12_bits_uop_br_mask <= stq_12_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1440) begin
        if (_GEN_1376) begin
          if (_GEN_1344) begin
            if (_GEN_1280) begin
            end
            else
              stq_12_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_12_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_12_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_12_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1440) begin
        if (_GEN_1376) begin
          if (_GEN_1344) begin
            if (_GEN_1280) begin
            end
            else begin
              stq_12_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_12_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_12_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_12_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_12_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_12_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_12_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_12_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_12_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_12_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_12_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_12_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1692) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_12_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_12_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_12_bits_uop_pdst <= casez_tmp_60;
        else
          stq_12_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1597) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_12_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_12_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_12_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1440) begin
        if (_GEN_1376) begin
          if (_GEN_1344) begin
            if (_GEN_1280) begin
            end
            else
              stq_12_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_12_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_12_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_12_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1440) begin
        if (_GEN_1376) begin
          if (_GEN_1344) begin
            if (_GEN_1280) begin
            end
            else begin
              stq_12_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_12_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_12_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_12_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_12_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_12_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_12_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_12_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_12_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_12_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_12_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_12_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_13_valid)
        stq_13_bits_uop_br_mask <= stq_13_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1441) begin
        if (_GEN_1377) begin
          if (_GEN_1345) begin
            if (_GEN_1281) begin
            end
            else
              stq_13_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_13_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_13_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_13_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1441) begin
        if (_GEN_1377) begin
          if (_GEN_1345) begin
            if (_GEN_1281) begin
            end
            else begin
              stq_13_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_13_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_13_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_13_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_13_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_13_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_13_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_13_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_13_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_13_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_13_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_13_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1693) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_13_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_13_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_13_bits_uop_pdst <= casez_tmp_60;
        else
          stq_13_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1598) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_13_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_13_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_13_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1441) begin
        if (_GEN_1377) begin
          if (_GEN_1345) begin
            if (_GEN_1281) begin
            end
            else
              stq_13_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_13_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_13_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_13_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1441) begin
        if (_GEN_1377) begin
          if (_GEN_1345) begin
            if (_GEN_1281) begin
            end
            else begin
              stq_13_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_13_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_13_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_13_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_13_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_13_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_13_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_13_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_13_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_13_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_13_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_13_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_14_valid)
        stq_14_bits_uop_br_mask <= stq_14_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1442) begin
        if (_GEN_1378) begin
          if (_GEN_1346) begin
            if (_GEN_1282) begin
            end
            else
              stq_14_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_14_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_14_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_14_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1442) begin
        if (_GEN_1378) begin
          if (_GEN_1346) begin
            if (_GEN_1282) begin
            end
            else begin
              stq_14_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_14_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_14_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_14_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_14_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_14_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_14_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_14_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_14_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_14_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_14_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_14_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1694) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_14_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_14_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_14_bits_uop_pdst <= casez_tmp_60;
        else
          stq_14_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1599) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_14_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_14_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_14_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1442) begin
        if (_GEN_1378) begin
          if (_GEN_1346) begin
            if (_GEN_1282) begin
            end
            else
              stq_14_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_14_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_14_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_14_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1442) begin
        if (_GEN_1378) begin
          if (_GEN_1346) begin
            if (_GEN_1282) begin
            end
            else begin
              stq_14_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_14_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_14_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_14_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_14_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_14_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_14_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_14_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_14_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_14_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_14_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_14_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_15_valid)
        stq_15_bits_uop_br_mask <= stq_15_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1443) begin
        if (_GEN_1379) begin
          if (_GEN_1347) begin
            if (_GEN_1283) begin
            end
            else
              stq_15_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_15_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_15_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_15_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1443) begin
        if (_GEN_1379) begin
          if (_GEN_1347) begin
            if (_GEN_1283) begin
            end
            else begin
              stq_15_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_15_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_15_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_15_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_15_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_15_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_15_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_15_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_15_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_15_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_15_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_15_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1695) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_15_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_15_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_15_bits_uop_pdst <= casez_tmp_60;
        else
          stq_15_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1600) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_15_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_15_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_15_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1443) begin
        if (_GEN_1379) begin
          if (_GEN_1347) begin
            if (_GEN_1283) begin
            end
            else
              stq_15_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_15_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_15_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_15_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1443) begin
        if (_GEN_1379) begin
          if (_GEN_1347) begin
            if (_GEN_1283) begin
            end
            else begin
              stq_15_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_15_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_15_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_15_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_15_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_15_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_15_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_15_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_15_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_15_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_15_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_15_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_16_valid)
        stq_16_bits_uop_br_mask <= stq_16_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1444) begin
        if (_GEN_1380) begin
          if (_GEN_1348) begin
            if (_GEN_1284) begin
            end
            else
              stq_16_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_16_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_16_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_16_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1444) begin
        if (_GEN_1380) begin
          if (_GEN_1348) begin
            if (_GEN_1284) begin
            end
            else begin
              stq_16_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_16_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_16_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_16_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_16_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_16_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_16_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_16_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_16_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_16_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_16_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_16_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1696) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_16_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_16_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_16_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_16_bits_uop_pdst <= casez_tmp_60;
        else
          stq_16_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1601) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_16_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_16_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_16_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1444) begin
        if (_GEN_1380) begin
          if (_GEN_1348) begin
            if (_GEN_1284) begin
            end
            else
              stq_16_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_16_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_16_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_16_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1444) begin
        if (_GEN_1380) begin
          if (_GEN_1348) begin
            if (_GEN_1284) begin
            end
            else begin
              stq_16_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_16_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_16_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_16_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_16_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_16_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_16_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_16_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_16_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_16_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_16_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_16_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_17_valid)
        stq_17_bits_uop_br_mask <= stq_17_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1445) begin
        if (_GEN_1381) begin
          if (_GEN_1349) begin
            if (_GEN_1285) begin
            end
            else
              stq_17_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_17_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_17_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_17_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1445) begin
        if (_GEN_1381) begin
          if (_GEN_1349) begin
            if (_GEN_1285) begin
            end
            else begin
              stq_17_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_17_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_17_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_17_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_17_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_17_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_17_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_17_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_17_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_17_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_17_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_17_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1697) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_17_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_17_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_17_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_17_bits_uop_pdst <= casez_tmp_60;
        else
          stq_17_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1602) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_17_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_17_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_17_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1445) begin
        if (_GEN_1381) begin
          if (_GEN_1349) begin
            if (_GEN_1285) begin
            end
            else
              stq_17_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_17_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_17_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_17_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1445) begin
        if (_GEN_1381) begin
          if (_GEN_1349) begin
            if (_GEN_1285) begin
            end
            else begin
              stq_17_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_17_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_17_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_17_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_17_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_17_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_17_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_17_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_17_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_17_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_17_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_17_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_18_valid)
        stq_18_bits_uop_br_mask <= stq_18_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1446) begin
        if (_GEN_1382) begin
          if (_GEN_1350) begin
            if (_GEN_1286) begin
            end
            else
              stq_18_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_18_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_18_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_18_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1446) begin
        if (_GEN_1382) begin
          if (_GEN_1350) begin
            if (_GEN_1286) begin
            end
            else begin
              stq_18_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_18_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_18_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_18_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_18_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_18_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_18_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_18_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_18_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_18_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_18_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_18_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1698) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_18_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_18_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_18_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_18_bits_uop_pdst <= casez_tmp_60;
        else
          stq_18_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1603) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_18_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_18_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_18_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1446) begin
        if (_GEN_1382) begin
          if (_GEN_1350) begin
            if (_GEN_1286) begin
            end
            else
              stq_18_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_18_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_18_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_18_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1446) begin
        if (_GEN_1382) begin
          if (_GEN_1350) begin
            if (_GEN_1286) begin
            end
            else begin
              stq_18_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_18_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_18_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_18_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_18_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_18_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_18_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_18_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_18_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_18_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_18_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_18_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_19_valid)
        stq_19_bits_uop_br_mask <= stq_19_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1447) begin
        if (_GEN_1383) begin
          if (_GEN_1351) begin
            if (_GEN_1287) begin
            end
            else
              stq_19_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_19_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_19_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_19_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1447) begin
        if (_GEN_1383) begin
          if (_GEN_1351) begin
            if (_GEN_1287) begin
            end
            else begin
              stq_19_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_19_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_19_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_19_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_19_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_19_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_19_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_19_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_19_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_19_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_19_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_19_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1699) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_19_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_19_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_19_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_19_bits_uop_pdst <= casez_tmp_60;
        else
          stq_19_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1604) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_19_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_19_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_19_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1447) begin
        if (_GEN_1383) begin
          if (_GEN_1351) begin
            if (_GEN_1287) begin
            end
            else
              stq_19_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_19_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_19_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_19_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1447) begin
        if (_GEN_1383) begin
          if (_GEN_1351) begin
            if (_GEN_1287) begin
            end
            else begin
              stq_19_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_19_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_19_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_19_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_19_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_19_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_19_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_19_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_19_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_19_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_19_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_19_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_20_valid)
        stq_20_bits_uop_br_mask <= stq_20_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1448) begin
        if (_GEN_1384) begin
          if (_GEN_1352) begin
            if (_GEN_1288) begin
            end
            else
              stq_20_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_20_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_20_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_20_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1448) begin
        if (_GEN_1384) begin
          if (_GEN_1352) begin
            if (_GEN_1288) begin
            end
            else begin
              stq_20_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_20_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_20_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_20_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_20_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_20_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_20_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_20_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_20_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_20_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_20_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_20_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1700) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_20_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_20_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_20_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_20_bits_uop_pdst <= casez_tmp_60;
        else
          stq_20_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1605) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_20_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_20_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_20_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1448) begin
        if (_GEN_1384) begin
          if (_GEN_1352) begin
            if (_GEN_1288) begin
            end
            else
              stq_20_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_20_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_20_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_20_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1448) begin
        if (_GEN_1384) begin
          if (_GEN_1352) begin
            if (_GEN_1288) begin
            end
            else begin
              stq_20_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_20_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_20_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_20_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_20_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_20_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_20_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_20_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_20_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_20_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_20_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_20_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_21_valid)
        stq_21_bits_uop_br_mask <= stq_21_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1449) begin
        if (_GEN_1385) begin
          if (_GEN_1353) begin
            if (_GEN_1289) begin
            end
            else
              stq_21_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_21_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_21_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_21_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1449) begin
        if (_GEN_1385) begin
          if (_GEN_1353) begin
            if (_GEN_1289) begin
            end
            else begin
              stq_21_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_21_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_21_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_21_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_21_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_21_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_21_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_21_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_21_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_21_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_21_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_21_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1701) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_21_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_21_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_21_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_21_bits_uop_pdst <= casez_tmp_60;
        else
          stq_21_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1606) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_21_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_21_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_21_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1449) begin
        if (_GEN_1385) begin
          if (_GEN_1353) begin
            if (_GEN_1289) begin
            end
            else
              stq_21_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_21_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_21_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_21_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1449) begin
        if (_GEN_1385) begin
          if (_GEN_1353) begin
            if (_GEN_1289) begin
            end
            else begin
              stq_21_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_21_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_21_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_21_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_21_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_21_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_21_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_21_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_21_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_21_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_21_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_21_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_22_valid)
        stq_22_bits_uop_br_mask <= stq_22_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1450) begin
        if (_GEN_1386) begin
          if (_GEN_1354) begin
            if (_GEN_1290) begin
            end
            else
              stq_22_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_22_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_22_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_22_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1450) begin
        if (_GEN_1386) begin
          if (_GEN_1354) begin
            if (_GEN_1290) begin
            end
            else begin
              stq_22_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_22_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_22_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_22_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_22_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_22_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_22_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_22_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_22_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_22_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_22_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_22_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1702) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_22_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_22_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_22_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_22_bits_uop_pdst <= casez_tmp_60;
        else
          stq_22_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1607) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_22_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_22_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_22_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1450) begin
        if (_GEN_1386) begin
          if (_GEN_1354) begin
            if (_GEN_1290) begin
            end
            else
              stq_22_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_22_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_22_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_22_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1450) begin
        if (_GEN_1386) begin
          if (_GEN_1354) begin
            if (_GEN_1290) begin
            end
            else begin
              stq_22_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_22_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_22_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_22_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_22_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_22_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_22_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_22_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_22_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_22_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_22_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_22_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_23_valid)
        stq_23_bits_uop_br_mask <= stq_23_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1451) begin
        if (_GEN_1387) begin
          if (_GEN_1355) begin
            if (_GEN_1291) begin
            end
            else
              stq_23_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_23_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_23_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_23_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1451) begin
        if (_GEN_1387) begin
          if (_GEN_1355) begin
            if (_GEN_1291) begin
            end
            else begin
              stq_23_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_23_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_23_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_23_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_23_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_23_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_23_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_23_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_23_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_23_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_23_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_23_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1703) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_23_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_23_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_23_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_23_bits_uop_pdst <= casez_tmp_60;
        else
          stq_23_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1608) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_23_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_23_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_23_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1451) begin
        if (_GEN_1387) begin
          if (_GEN_1355) begin
            if (_GEN_1291) begin
            end
            else
              stq_23_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_23_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_23_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_23_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1451) begin
        if (_GEN_1387) begin
          if (_GEN_1355) begin
            if (_GEN_1291) begin
            end
            else begin
              stq_23_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_23_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_23_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_23_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_23_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_23_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_23_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_23_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_23_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_23_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_23_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_23_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_24_valid)
        stq_24_bits_uop_br_mask <= stq_24_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1452) begin
        if (_GEN_1388) begin
          if (_GEN_1356) begin
            if (_GEN_1292) begin
            end
            else
              stq_24_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_24_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_24_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_24_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1452) begin
        if (_GEN_1388) begin
          if (_GEN_1356) begin
            if (_GEN_1292) begin
            end
            else begin
              stq_24_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_24_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_24_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_24_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_24_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_24_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_24_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_24_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_24_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_24_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_24_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_24_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1704) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_24_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_24_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_24_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_24_bits_uop_pdst <= casez_tmp_60;
        else
          stq_24_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1609) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_24_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_24_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_24_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1452) begin
        if (_GEN_1388) begin
          if (_GEN_1356) begin
            if (_GEN_1292) begin
            end
            else
              stq_24_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_24_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_24_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_24_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1452) begin
        if (_GEN_1388) begin
          if (_GEN_1356) begin
            if (_GEN_1292) begin
            end
            else begin
              stq_24_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_24_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_24_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_24_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_24_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_24_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_24_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_24_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_24_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_24_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_24_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_24_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_25_valid)
        stq_25_bits_uop_br_mask <= stq_25_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1453) begin
        if (_GEN_1389) begin
          if (_GEN_1357) begin
            if (_GEN_1293) begin
            end
            else
              stq_25_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_25_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_25_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_25_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1453) begin
        if (_GEN_1389) begin
          if (_GEN_1357) begin
            if (_GEN_1293) begin
            end
            else begin
              stq_25_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_25_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_25_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_25_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_25_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_25_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_25_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_25_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_25_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_25_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_25_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_25_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1705) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_25_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_25_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_25_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_25_bits_uop_pdst <= casez_tmp_60;
        else
          stq_25_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1610) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_25_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_25_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_25_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1453) begin
        if (_GEN_1389) begin
          if (_GEN_1357) begin
            if (_GEN_1293) begin
            end
            else
              stq_25_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_25_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_25_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_25_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1453) begin
        if (_GEN_1389) begin
          if (_GEN_1357) begin
            if (_GEN_1293) begin
            end
            else begin
              stq_25_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_25_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_25_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_25_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_25_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_25_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_25_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_25_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_25_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_25_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_25_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_25_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_26_valid)
        stq_26_bits_uop_br_mask <= stq_26_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1454) begin
        if (_GEN_1390) begin
          if (_GEN_1358) begin
            if (_GEN_1294) begin
            end
            else
              stq_26_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_26_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_26_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_26_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1454) begin
        if (_GEN_1390) begin
          if (_GEN_1358) begin
            if (_GEN_1294) begin
            end
            else begin
              stq_26_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_26_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_26_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_26_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_26_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_26_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_26_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_26_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_26_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_26_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_26_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_26_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1706) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_26_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_26_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_26_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_26_bits_uop_pdst <= casez_tmp_60;
        else
          stq_26_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1611) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_26_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_26_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_26_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1454) begin
        if (_GEN_1390) begin
          if (_GEN_1358) begin
            if (_GEN_1294) begin
            end
            else
              stq_26_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_26_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_26_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_26_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1454) begin
        if (_GEN_1390) begin
          if (_GEN_1358) begin
            if (_GEN_1294) begin
            end
            else begin
              stq_26_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_26_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_26_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_26_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_26_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_26_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_26_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_26_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_26_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_26_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_26_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_26_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_27_valid)
        stq_27_bits_uop_br_mask <= stq_27_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1455) begin
        if (_GEN_1391) begin
          if (_GEN_1359) begin
            if (_GEN_1295) begin
            end
            else
              stq_27_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_27_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_27_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_27_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1455) begin
        if (_GEN_1391) begin
          if (_GEN_1359) begin
            if (_GEN_1295) begin
            end
            else begin
              stq_27_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_27_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_27_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_27_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_27_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_27_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_27_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_27_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_27_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_27_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_27_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_27_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1707) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_27_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_27_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_27_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_27_bits_uop_pdst <= casez_tmp_60;
        else
          stq_27_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1612) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_27_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_27_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_27_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1455) begin
        if (_GEN_1391) begin
          if (_GEN_1359) begin
            if (_GEN_1295) begin
            end
            else
              stq_27_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_27_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_27_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_27_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1455) begin
        if (_GEN_1391) begin
          if (_GEN_1359) begin
            if (_GEN_1295) begin
            end
            else begin
              stq_27_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_27_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_27_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_27_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_27_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_27_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_27_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_27_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_27_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_27_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_27_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_27_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_28_valid)
        stq_28_bits_uop_br_mask <= stq_28_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1456) begin
        if (_GEN_1392) begin
          if (_GEN_1360) begin
            if (_GEN_1296) begin
            end
            else
              stq_28_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_28_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_28_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_28_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1456) begin
        if (_GEN_1392) begin
          if (_GEN_1360) begin
            if (_GEN_1296) begin
            end
            else begin
              stq_28_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_28_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_28_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_28_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_28_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_28_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_28_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_28_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_28_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_28_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_28_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_28_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1708) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_28_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_28_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_28_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_28_bits_uop_pdst <= casez_tmp_60;
        else
          stq_28_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1613) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_28_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_28_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_28_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1456) begin
        if (_GEN_1392) begin
          if (_GEN_1360) begin
            if (_GEN_1296) begin
            end
            else
              stq_28_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_28_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_28_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_28_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1456) begin
        if (_GEN_1392) begin
          if (_GEN_1360) begin
            if (_GEN_1296) begin
            end
            else begin
              stq_28_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_28_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_28_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_28_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_28_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_28_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_28_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_28_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_28_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_28_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_28_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_28_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_29_valid)
        stq_29_bits_uop_br_mask <= stq_29_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1457) begin
        if (_GEN_1393) begin
          if (_GEN_1361) begin
            if (_GEN_1297) begin
            end
            else
              stq_29_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_29_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_29_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_29_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1457) begin
        if (_GEN_1393) begin
          if (_GEN_1361) begin
            if (_GEN_1297) begin
            end
            else begin
              stq_29_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_29_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_29_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_29_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_29_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_29_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_29_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_29_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_29_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_29_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_29_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_29_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1709) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_29_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_29_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_29_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_29_bits_uop_pdst <= casez_tmp_60;
        else
          stq_29_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1614) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_29_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_29_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_29_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1457) begin
        if (_GEN_1393) begin
          if (_GEN_1361) begin
            if (_GEN_1297) begin
            end
            else
              stq_29_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_29_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_29_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_29_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1457) begin
        if (_GEN_1393) begin
          if (_GEN_1361) begin
            if (_GEN_1297) begin
            end
            else begin
              stq_29_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_29_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_29_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_29_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_29_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_29_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_29_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_29_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_29_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_29_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_29_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_29_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_30_valid)
        stq_30_bits_uop_br_mask <= stq_30_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1458) begin
        if (_GEN_1394) begin
          if (_GEN_1362) begin
            if (_GEN_1298) begin
            end
            else
              stq_30_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_30_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_30_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_30_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1458) begin
        if (_GEN_1394) begin
          if (_GEN_1362) begin
            if (_GEN_1298) begin
            end
            else begin
              stq_30_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_30_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_30_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_30_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_30_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_30_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_30_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_30_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_30_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_30_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_30_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_30_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1710) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_30_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_30_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_30_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_30_bits_uop_pdst <= casez_tmp_60;
        else
          stq_30_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1615) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_30_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_30_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_30_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1458) begin
        if (_GEN_1394) begin
          if (_GEN_1362) begin
            if (_GEN_1298) begin
            end
            else
              stq_30_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_30_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_30_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_30_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1458) begin
        if (_GEN_1394) begin
          if (_GEN_1362) begin
            if (_GEN_1298) begin
            end
            else begin
              stq_30_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_30_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_30_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_30_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_30_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_30_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_30_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_30_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_30_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_30_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_30_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_30_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (stq_31_valid)
        stq_31_bits_uop_br_mask <= stq_31_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
      else if (_GEN_1459) begin
        if (_GEN_1395) begin
          if (_GEN_1363) begin
            if (_GEN_1299) begin
            end
            else
              stq_31_bits_uop_br_mask <= io_core_dis_uops_0_bits_br_mask;
          end
          else
            stq_31_bits_uop_br_mask <= io_core_dis_uops_1_bits_br_mask;
        end
        else
          stq_31_bits_uop_br_mask <= io_core_dis_uops_2_bits_br_mask;
      end
      else
        stq_31_bits_uop_br_mask <= io_core_dis_uops_3_bits_br_mask;
      if (_GEN_1459) begin
        if (_GEN_1395) begin
          if (_GEN_1363) begin
            if (_GEN_1299) begin
            end
            else begin
              stq_31_bits_uop_rob_idx <= io_core_dis_uops_0_bits_rob_idx;
              stq_31_bits_uop_ldq_idx <= io_core_dis_uops_0_bits_ldq_idx;
              stq_31_bits_uop_stq_idx <= io_core_dis_uops_0_bits_stq_idx;
            end
          end
          else begin
            stq_31_bits_uop_rob_idx <= io_core_dis_uops_1_bits_rob_idx;
            stq_31_bits_uop_ldq_idx <= io_core_dis_uops_1_bits_ldq_idx;
            stq_31_bits_uop_stq_idx <= io_core_dis_uops_1_bits_stq_idx;
          end
        end
        else begin
          stq_31_bits_uop_rob_idx <= io_core_dis_uops_2_bits_rob_idx;
          stq_31_bits_uop_ldq_idx <= io_core_dis_uops_2_bits_ldq_idx;
          stq_31_bits_uop_stq_idx <= io_core_dis_uops_2_bits_stq_idx;
        end
      end
      else begin
        stq_31_bits_uop_rob_idx <= io_core_dis_uops_3_bits_rob_idx;
        stq_31_bits_uop_ldq_idx <= io_core_dis_uops_3_bits_ldq_idx;
        stq_31_bits_uop_stq_idx <= io_core_dis_uops_3_bits_stq_idx;
      end
      if (_GEN_1711) begin
        if (_exe_tlb_uop_T_9) begin
          if (_GEN_329)
            stq_31_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_31_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else if (will_fire_load_retry_1)
          stq_31_bits_uop_pdst <= casez_tmp_71;
        else if (will_fire_sta_retry_1)
          stq_31_bits_uop_pdst <= casez_tmp_60;
        else
          stq_31_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1616) begin
        if (_exe_tlb_uop_T_2) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_31_bits_uop_pdst <= io_core_exe_1_req_bits_uop_pdst;
          else
            stq_31_bits_uop_pdst <= io_core_exe_0_req_bits_uop_pdst;
        end
        else
          stq_31_bits_uop_pdst <= 7'h0;
      end
      else if (_GEN_1459) begin
        if (_GEN_1395) begin
          if (_GEN_1363) begin
            if (_GEN_1299) begin
            end
            else
              stq_31_bits_uop_pdst <= io_core_dis_uops_0_bits_pdst;
          end
          else
            stq_31_bits_uop_pdst <= io_core_dis_uops_1_bits_pdst;
        end
        else
          stq_31_bits_uop_pdst <= io_core_dis_uops_2_bits_pdst;
      end
      else
        stq_31_bits_uop_pdst <= io_core_dis_uops_3_bits_pdst;
      if (_GEN_1459) begin
        if (_GEN_1395) begin
          if (_GEN_1363) begin
            if (_GEN_1299) begin
            end
            else begin
              stq_31_bits_uop_mem_cmd <= io_core_dis_uops_0_bits_mem_cmd;
              stq_31_bits_uop_mem_size <= io_core_dis_uops_0_bits_mem_size;
              stq_31_bits_uop_dst_rtype <= io_core_dis_uops_0_bits_dst_rtype;
            end
          end
          else begin
            stq_31_bits_uop_mem_cmd <= io_core_dis_uops_1_bits_mem_cmd;
            stq_31_bits_uop_mem_size <= io_core_dis_uops_1_bits_mem_size;
            stq_31_bits_uop_dst_rtype <= io_core_dis_uops_1_bits_dst_rtype;
          end
        end
        else begin
          stq_31_bits_uop_mem_cmd <= io_core_dis_uops_2_bits_mem_cmd;
          stq_31_bits_uop_mem_size <= io_core_dis_uops_2_bits_mem_size;
          stq_31_bits_uop_dst_rtype <= io_core_dis_uops_2_bits_dst_rtype;
        end
      end
      else begin
        stq_31_bits_uop_mem_cmd <= io_core_dis_uops_3_bits_mem_cmd;
        stq_31_bits_uop_mem_size <= io_core_dis_uops_3_bits_mem_size;
        stq_31_bits_uop_dst_rtype <= io_core_dis_uops_3_bits_dst_rtype;
      end
      if (clear_store)
        stq_head <= stq_head + 5'h1;
      if (commit_store_3)
        stq_commit_head <= _GEN_1227 + 5'h1;
      else if (commit_store_2)
        stq_commit_head <= _GEN_1226;
      else if (commit_store_1)
        stq_commit_head <= _GEN_1222;
      else if (commit_store)
        stq_commit_head <= _GEN_1218;
      if (clear_store & casez_tmp_2)
        stq_execute_head <= _stq_execute_head_T_8;
      else if (~io_dmem_nack_1_valid | io_dmem_nack_1_bits_is_hella | io_dmem_nack_1_bits_uop_uses_ldq | io_dmem_nack_1_bits_uop_stq_idx < stq_head ^ _GEN_1236 ^ io_dmem_nack_1_bits_uop_stq_idx >= stq_execute_head) begin
        if (~io_dmem_nack_0_valid | io_dmem_nack_0_bits_is_hella | io_dmem_nack_0_bits_uop_uses_ldq | io_dmem_nack_0_bits_uop_stq_idx < stq_head ^ _GEN_1236 ^ io_dmem_nack_0_bits_uop_stq_idx >= stq_execute_head) begin
          if (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & dmem_req_fire_0)) begin
          end
          else
            stq_execute_head <= _stq_execute_head_T_8;
        end
        else
          stq_execute_head <= io_dmem_nack_0_bits_uop_stq_idx;
      end
      else
        stq_execute_head <= io_dmem_nack_1_bits_uop_stq_idx;
    end
    stq_0_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h0 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h0 | (_GEN_1428 ? (_GEN_1364 ? (_GEN_1332 ? (_GEN_1268 ? stq_0_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_0_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1428 ? (_GEN_1364 ? (_GEN_1332 ? (_GEN_1268 ? stq_0_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_0_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1428 ? (_GEN_1364 ? (_GEN_1332 ? (_GEN_1268 ? stq_0_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_0_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1428 ? (_GEN_1364 ? (_GEN_1332 ? (_GEN_1268 ? stq_0_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_0_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1428 ? (_GEN_1364 ? (_GEN_1332 ? (_GEN_1268 ? stq_0_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_0_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1428 ? (_GEN_1364 ? (_GEN_1332 ? (_GEN_1268 ? stq_0_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_0_bits_addr_valid <= ~_GEN_2479 & (clear_store ? ~_GEN_2411 & _GEN_82006 : ~_GEN_1997 & _GEN_82006);
    if (_GEN_1680) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_0_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_0_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_0_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_0_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_0_bits_addr_bits <= hella_req_addr;
        else
          stq_0_bits_addr_bits <= 40'h0;
      end
      else
        stq_0_bits_addr_bits <= _GEN_338;
      stq_0_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1585) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_0_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_0_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_0_bits_addr_bits <= _GEN_332;
        else
          stq_0_bits_addr_bits <= 40'h0;
      end
      else
        stq_0_bits_addr_bits <= _GEN_334;
      stq_0_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_0_bits_data_valid <= ~_GEN_2479 & (clear_store ? ~_GEN_2411 & _GEN_82230 : ~_GEN_1997 & _GEN_82230);
    if (_stq_bits_data_bits_T_2 & _GEN_1712) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_0_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_0_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_0_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1617) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_0_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_0_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_0_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_0_bits_committed <= ~_GEN_2443 & (commit_store_3 ? _GEN_2347 | _GEN_2283 | _GEN_137950 : _GEN_2283 | _GEN_137950);
    stq_0_bits_succeeded <= ~_GEN_2443 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h0 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h0 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h0)) & _GEN_1428 & _GEN_1364 & _GEN_1332 & _GEN_1268 & stq_0_bits_succeeded);
    stq_1_valid <= ~_GEN_2480 & (clear_store ? ~_GEN_2412 & _GEN_52417 : ~_GEN_1998 & _GEN_52417);
    stq_1_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1 | (_GEN_1429 ? (_GEN_1365 ? (_GEN_1333 ? (_GEN_1269 ? stq_1_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_1_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1429 ? (_GEN_1365 ? (_GEN_1333 ? (_GEN_1269 ? stq_1_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_1_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1429 ? (_GEN_1365 ? (_GEN_1333 ? (_GEN_1269 ? stq_1_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_1_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1429 ? (_GEN_1365 ? (_GEN_1333 ? (_GEN_1269 ? stq_1_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_1_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1429 ? (_GEN_1365 ? (_GEN_1333 ? (_GEN_1269 ? stq_1_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_1_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1429 ? (_GEN_1365 ? (_GEN_1333 ? (_GEN_1269 ? stq_1_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_1_bits_addr_valid <= ~_GEN_2480 & (clear_store ? ~_GEN_2412 & _GEN_82007 : ~_GEN_1998 & _GEN_82007);
    if (_GEN_1681) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_1_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_1_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_1_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_1_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_1_bits_addr_bits <= hella_req_addr;
        else
          stq_1_bits_addr_bits <= 40'h0;
      end
      else
        stq_1_bits_addr_bits <= _GEN_338;
      stq_1_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1586) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_1_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_1_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_1_bits_addr_bits <= _GEN_332;
        else
          stq_1_bits_addr_bits <= 40'h0;
      end
      else
        stq_1_bits_addr_bits <= _GEN_334;
      stq_1_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_1_bits_data_valid <= ~_GEN_2480 & (clear_store ? ~_GEN_2412 & _GEN_82231 : ~_GEN_1998 & _GEN_82231);
    if (_stq_bits_data_bits_T_2 & _GEN_1713) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_1_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_1_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_1_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1618) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_1_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_1_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_1_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_1_bits_committed <= ~_GEN_2444 & (commit_store_3 ? _GEN_2348 | _GEN_2284 | _GEN_137951 : _GEN_2284 | _GEN_137951);
    stq_1_bits_succeeded <= ~_GEN_2444 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h1)) & _GEN_1429 & _GEN_1365 & _GEN_1333 & _GEN_1269 & stq_1_bits_succeeded);
    stq_2_valid <= ~_GEN_2481 & (clear_store ? ~_GEN_2413 & _GEN_52418 : ~_GEN_1999 & _GEN_52418);
    stq_2_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h2 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h2 | (_GEN_1430 ? (_GEN_1366 ? (_GEN_1334 ? (_GEN_1270 ? stq_2_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_2_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1430 ? (_GEN_1366 ? (_GEN_1334 ? (_GEN_1270 ? stq_2_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_2_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1430 ? (_GEN_1366 ? (_GEN_1334 ? (_GEN_1270 ? stq_2_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_2_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1430 ? (_GEN_1366 ? (_GEN_1334 ? (_GEN_1270 ? stq_2_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_2_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1430 ? (_GEN_1366 ? (_GEN_1334 ? (_GEN_1270 ? stq_2_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_2_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1430 ? (_GEN_1366 ? (_GEN_1334 ? (_GEN_1270 ? stq_2_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_2_bits_addr_valid <= ~_GEN_2481 & (clear_store ? ~_GEN_2413 & _GEN_82008 : ~_GEN_1999 & _GEN_82008);
    if (_GEN_1682) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_2_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_2_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_2_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_2_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_2_bits_addr_bits <= hella_req_addr;
        else
          stq_2_bits_addr_bits <= 40'h0;
      end
      else
        stq_2_bits_addr_bits <= _GEN_338;
      stq_2_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1587) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_2_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_2_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_2_bits_addr_bits <= _GEN_332;
        else
          stq_2_bits_addr_bits <= 40'h0;
      end
      else
        stq_2_bits_addr_bits <= _GEN_334;
      stq_2_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_2_bits_data_valid <= ~_GEN_2481 & (clear_store ? ~_GEN_2413 & _GEN_82232 : ~_GEN_1999 & _GEN_82232);
    if (_stq_bits_data_bits_T_2 & _GEN_1714) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_2_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_2_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_2_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1619) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_2_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_2_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_2_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_2_bits_committed <= ~_GEN_2445 & (commit_store_3 ? _GEN_2349 | _GEN_2285 | _GEN_137952 : _GEN_2285 | _GEN_137952);
    stq_2_bits_succeeded <= ~_GEN_2445 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h2 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h2 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h2)) & _GEN_1430 & _GEN_1366 & _GEN_1334 & _GEN_1270 & stq_2_bits_succeeded);
    stq_3_valid <= ~_GEN_2482 & (clear_store ? ~_GEN_2414 & _GEN_52419 : ~_GEN_2000 & _GEN_52419);
    stq_3_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h3 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h3 | (_GEN_1431 ? (_GEN_1367 ? (_GEN_1335 ? (_GEN_1271 ? stq_3_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_3_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1431 ? (_GEN_1367 ? (_GEN_1335 ? (_GEN_1271 ? stq_3_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_3_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1431 ? (_GEN_1367 ? (_GEN_1335 ? (_GEN_1271 ? stq_3_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_3_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1431 ? (_GEN_1367 ? (_GEN_1335 ? (_GEN_1271 ? stq_3_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_3_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1431 ? (_GEN_1367 ? (_GEN_1335 ? (_GEN_1271 ? stq_3_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_3_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1431 ? (_GEN_1367 ? (_GEN_1335 ? (_GEN_1271 ? stq_3_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_3_bits_addr_valid <= ~_GEN_2482 & (clear_store ? ~_GEN_2414 & _GEN_82009 : ~_GEN_2000 & _GEN_82009);
    if (_GEN_1683) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_3_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_3_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_3_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_3_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_3_bits_addr_bits <= hella_req_addr;
        else
          stq_3_bits_addr_bits <= 40'h0;
      end
      else
        stq_3_bits_addr_bits <= _GEN_338;
      stq_3_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1588) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_3_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_3_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_3_bits_addr_bits <= _GEN_332;
        else
          stq_3_bits_addr_bits <= 40'h0;
      end
      else
        stq_3_bits_addr_bits <= _GEN_334;
      stq_3_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_3_bits_data_valid <= ~_GEN_2482 & (clear_store ? ~_GEN_2414 & _GEN_82233 : ~_GEN_2000 & _GEN_82233);
    if (_stq_bits_data_bits_T_2 & _GEN_1715) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_3_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_3_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_3_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1620) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_3_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_3_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_3_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_3_bits_committed <= ~_GEN_2446 & (commit_store_3 ? _GEN_2350 | _GEN_2286 | _GEN_137953 : _GEN_2286 | _GEN_137953);
    stq_3_bits_succeeded <= ~_GEN_2446 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h3 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h3 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h3)) & _GEN_1431 & _GEN_1367 & _GEN_1335 & _GEN_1271 & stq_3_bits_succeeded);
    stq_4_valid <= ~_GEN_2483 & (clear_store ? ~_GEN_2415 & _GEN_52420 : ~_GEN_2001 & _GEN_52420);
    stq_4_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h4 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h4 | (_GEN_1432 ? (_GEN_1368 ? (_GEN_1336 ? (_GEN_1272 ? stq_4_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_4_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1432 ? (_GEN_1368 ? (_GEN_1336 ? (_GEN_1272 ? stq_4_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_4_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1432 ? (_GEN_1368 ? (_GEN_1336 ? (_GEN_1272 ? stq_4_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_4_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1432 ? (_GEN_1368 ? (_GEN_1336 ? (_GEN_1272 ? stq_4_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_4_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1432 ? (_GEN_1368 ? (_GEN_1336 ? (_GEN_1272 ? stq_4_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_4_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1432 ? (_GEN_1368 ? (_GEN_1336 ? (_GEN_1272 ? stq_4_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_4_bits_addr_valid <= ~_GEN_2483 & (clear_store ? ~_GEN_2415 & _GEN_82010 : ~_GEN_2001 & _GEN_82010);
    if (_GEN_1684) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_4_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_4_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_4_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_4_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_4_bits_addr_bits <= hella_req_addr;
        else
          stq_4_bits_addr_bits <= 40'h0;
      end
      else
        stq_4_bits_addr_bits <= _GEN_338;
      stq_4_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1589) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_4_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_4_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_4_bits_addr_bits <= _GEN_332;
        else
          stq_4_bits_addr_bits <= 40'h0;
      end
      else
        stq_4_bits_addr_bits <= _GEN_334;
      stq_4_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_4_bits_data_valid <= ~_GEN_2483 & (clear_store ? ~_GEN_2415 & _GEN_82234 : ~_GEN_2001 & _GEN_82234);
    if (_stq_bits_data_bits_T_2 & _GEN_1716) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_4_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_4_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_4_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1621) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_4_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_4_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_4_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_4_bits_committed <= ~_GEN_2447 & (commit_store_3 ? _GEN_2351 | _GEN_2287 | _GEN_137954 : _GEN_2287 | _GEN_137954);
    stq_4_bits_succeeded <= ~_GEN_2447 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h4 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h4 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h4)) & _GEN_1432 & _GEN_1368 & _GEN_1336 & _GEN_1272 & stq_4_bits_succeeded);
    stq_5_valid <= ~_GEN_2484 & (clear_store ? ~_GEN_2416 & _GEN_52421 : ~_GEN_2002 & _GEN_52421);
    stq_5_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h5 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h5 | (_GEN_1433 ? (_GEN_1369 ? (_GEN_1337 ? (_GEN_1273 ? stq_5_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_5_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1433 ? (_GEN_1369 ? (_GEN_1337 ? (_GEN_1273 ? stq_5_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_5_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1433 ? (_GEN_1369 ? (_GEN_1337 ? (_GEN_1273 ? stq_5_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_5_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1433 ? (_GEN_1369 ? (_GEN_1337 ? (_GEN_1273 ? stq_5_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_5_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1433 ? (_GEN_1369 ? (_GEN_1337 ? (_GEN_1273 ? stq_5_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_5_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1433 ? (_GEN_1369 ? (_GEN_1337 ? (_GEN_1273 ? stq_5_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_5_bits_addr_valid <= ~_GEN_2484 & (clear_store ? ~_GEN_2416 & _GEN_82011 : ~_GEN_2002 & _GEN_82011);
    if (_GEN_1685) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_5_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_5_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_5_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_5_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_5_bits_addr_bits <= hella_req_addr;
        else
          stq_5_bits_addr_bits <= 40'h0;
      end
      else
        stq_5_bits_addr_bits <= _GEN_338;
      stq_5_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1590) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_5_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_5_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_5_bits_addr_bits <= _GEN_332;
        else
          stq_5_bits_addr_bits <= 40'h0;
      end
      else
        stq_5_bits_addr_bits <= _GEN_334;
      stq_5_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_5_bits_data_valid <= ~_GEN_2484 & (clear_store ? ~_GEN_2416 & _GEN_82235 : ~_GEN_2002 & _GEN_82235);
    if (_stq_bits_data_bits_T_2 & _GEN_1717) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_5_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_5_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_5_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1622) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_5_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_5_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_5_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_5_bits_committed <= ~_GEN_2448 & (commit_store_3 ? _GEN_2352 | _GEN_2288 | _GEN_137955 : _GEN_2288 | _GEN_137955);
    stq_5_bits_succeeded <= ~_GEN_2448 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h5 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h5 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h5)) & _GEN_1433 & _GEN_1369 & _GEN_1337 & _GEN_1273 & stq_5_bits_succeeded);
    stq_6_valid <= ~_GEN_2485 & (clear_store ? ~_GEN_2417 & _GEN_52422 : ~_GEN_2003 & _GEN_52422);
    stq_6_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h6 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h6 | (_GEN_1434 ? (_GEN_1370 ? (_GEN_1338 ? (_GEN_1274 ? stq_6_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_6_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1434 ? (_GEN_1370 ? (_GEN_1338 ? (_GEN_1274 ? stq_6_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_6_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1434 ? (_GEN_1370 ? (_GEN_1338 ? (_GEN_1274 ? stq_6_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_6_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1434 ? (_GEN_1370 ? (_GEN_1338 ? (_GEN_1274 ? stq_6_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_6_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1434 ? (_GEN_1370 ? (_GEN_1338 ? (_GEN_1274 ? stq_6_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_6_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1434 ? (_GEN_1370 ? (_GEN_1338 ? (_GEN_1274 ? stq_6_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_6_bits_addr_valid <= ~_GEN_2485 & (clear_store ? ~_GEN_2417 & _GEN_82012 : ~_GEN_2003 & _GEN_82012);
    if (_GEN_1686) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_6_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_6_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_6_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_6_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_6_bits_addr_bits <= hella_req_addr;
        else
          stq_6_bits_addr_bits <= 40'h0;
      end
      else
        stq_6_bits_addr_bits <= _GEN_338;
      stq_6_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1591) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_6_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_6_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_6_bits_addr_bits <= _GEN_332;
        else
          stq_6_bits_addr_bits <= 40'h0;
      end
      else
        stq_6_bits_addr_bits <= _GEN_334;
      stq_6_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_6_bits_data_valid <= ~_GEN_2485 & (clear_store ? ~_GEN_2417 & _GEN_82236 : ~_GEN_2003 & _GEN_82236);
    if (_stq_bits_data_bits_T_2 & _GEN_1718) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_6_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_6_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_6_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1623) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_6_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_6_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_6_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_6_bits_committed <= ~_GEN_2449 & (commit_store_3 ? _GEN_2353 | _GEN_2289 | _GEN_137956 : _GEN_2289 | _GEN_137956);
    stq_6_bits_succeeded <= ~_GEN_2449 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h6 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h6 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h6)) & _GEN_1434 & _GEN_1370 & _GEN_1338 & _GEN_1274 & stq_6_bits_succeeded);
    stq_7_valid <= ~_GEN_2486 & (clear_store ? ~_GEN_2418 & _GEN_52423 : ~_GEN_2004 & _GEN_52423);
    stq_7_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h7 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h7 | (_GEN_1435 ? (_GEN_1371 ? (_GEN_1339 ? (_GEN_1275 ? stq_7_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_7_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1435 ? (_GEN_1371 ? (_GEN_1339 ? (_GEN_1275 ? stq_7_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_7_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1435 ? (_GEN_1371 ? (_GEN_1339 ? (_GEN_1275 ? stq_7_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_7_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1435 ? (_GEN_1371 ? (_GEN_1339 ? (_GEN_1275 ? stq_7_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_7_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1435 ? (_GEN_1371 ? (_GEN_1339 ? (_GEN_1275 ? stq_7_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_7_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1435 ? (_GEN_1371 ? (_GEN_1339 ? (_GEN_1275 ? stq_7_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_7_bits_addr_valid <= ~_GEN_2486 & (clear_store ? ~_GEN_2418 & _GEN_82013 : ~_GEN_2004 & _GEN_82013);
    if (_GEN_1687) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_7_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_7_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_7_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_7_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_7_bits_addr_bits <= hella_req_addr;
        else
          stq_7_bits_addr_bits <= 40'h0;
      end
      else
        stq_7_bits_addr_bits <= _GEN_338;
      stq_7_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1592) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_7_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_7_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_7_bits_addr_bits <= _GEN_332;
        else
          stq_7_bits_addr_bits <= 40'h0;
      end
      else
        stq_7_bits_addr_bits <= _GEN_334;
      stq_7_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_7_bits_data_valid <= ~_GEN_2486 & (clear_store ? ~_GEN_2418 & _GEN_82237 : ~_GEN_2004 & _GEN_82237);
    if (_stq_bits_data_bits_T_2 & _GEN_1719) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_7_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_7_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_7_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1624) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_7_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_7_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_7_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_7_bits_committed <= ~_GEN_2450 & (commit_store_3 ? _GEN_2354 | _GEN_2290 | _GEN_137957 : _GEN_2290 | _GEN_137957);
    stq_7_bits_succeeded <= ~_GEN_2450 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h7 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h7 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h7)) & _GEN_1435 & _GEN_1371 & _GEN_1339 & _GEN_1275 & stq_7_bits_succeeded);
    stq_8_valid <= ~_GEN_2487 & (clear_store ? ~_GEN_2419 & _GEN_52424 : ~_GEN_2005 & _GEN_52424);
    stq_8_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h8 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h8 | (_GEN_1436 ? (_GEN_1372 ? (_GEN_1340 ? (_GEN_1276 ? stq_8_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_8_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1436 ? (_GEN_1372 ? (_GEN_1340 ? (_GEN_1276 ? stq_8_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_8_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1436 ? (_GEN_1372 ? (_GEN_1340 ? (_GEN_1276 ? stq_8_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_8_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1436 ? (_GEN_1372 ? (_GEN_1340 ? (_GEN_1276 ? stq_8_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_8_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1436 ? (_GEN_1372 ? (_GEN_1340 ? (_GEN_1276 ? stq_8_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_8_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1436 ? (_GEN_1372 ? (_GEN_1340 ? (_GEN_1276 ? stq_8_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_8_bits_addr_valid <= ~_GEN_2487 & (clear_store ? ~_GEN_2419 & _GEN_82014 : ~_GEN_2005 & _GEN_82014);
    if (_GEN_1688) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_8_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_8_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_8_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_8_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_8_bits_addr_bits <= hella_req_addr;
        else
          stq_8_bits_addr_bits <= 40'h0;
      end
      else
        stq_8_bits_addr_bits <= _GEN_338;
      stq_8_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1593) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_8_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_8_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_8_bits_addr_bits <= _GEN_332;
        else
          stq_8_bits_addr_bits <= 40'h0;
      end
      else
        stq_8_bits_addr_bits <= _GEN_334;
      stq_8_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_8_bits_data_valid <= ~_GEN_2487 & (clear_store ? ~_GEN_2419 & _GEN_82238 : ~_GEN_2005 & _GEN_82238);
    if (_stq_bits_data_bits_T_2 & _GEN_1720) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_8_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_8_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_8_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1625) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_8_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_8_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_8_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_8_bits_committed <= ~_GEN_2451 & (commit_store_3 ? _GEN_2355 | _GEN_2291 | _GEN_137958 : _GEN_2291 | _GEN_137958);
    stq_8_bits_succeeded <= ~_GEN_2451 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h8 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h8 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h8)) & _GEN_1436 & _GEN_1372 & _GEN_1340 & _GEN_1276 & stq_8_bits_succeeded);
    stq_9_valid <= ~_GEN_2488 & (clear_store ? ~_GEN_2420 & _GEN_52425 : ~_GEN_2006 & _GEN_52425);
    stq_9_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h9 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h9 | (_GEN_1437 ? (_GEN_1373 ? (_GEN_1341 ? (_GEN_1277 ? stq_9_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_9_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1437 ? (_GEN_1373 ? (_GEN_1341 ? (_GEN_1277 ? stq_9_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_9_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1437 ? (_GEN_1373 ? (_GEN_1341 ? (_GEN_1277 ? stq_9_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_9_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1437 ? (_GEN_1373 ? (_GEN_1341 ? (_GEN_1277 ? stq_9_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_9_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1437 ? (_GEN_1373 ? (_GEN_1341 ? (_GEN_1277 ? stq_9_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_9_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1437 ? (_GEN_1373 ? (_GEN_1341 ? (_GEN_1277 ? stq_9_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_9_bits_addr_valid <= ~_GEN_2488 & (clear_store ? ~_GEN_2420 & _GEN_82015 : ~_GEN_2006 & _GEN_82015);
    if (_GEN_1689) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_9_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_9_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_9_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_9_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_9_bits_addr_bits <= hella_req_addr;
        else
          stq_9_bits_addr_bits <= 40'h0;
      end
      else
        stq_9_bits_addr_bits <= _GEN_338;
      stq_9_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1594) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_9_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_9_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_9_bits_addr_bits <= _GEN_332;
        else
          stq_9_bits_addr_bits <= 40'h0;
      end
      else
        stq_9_bits_addr_bits <= _GEN_334;
      stq_9_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_9_bits_data_valid <= ~_GEN_2488 & (clear_store ? ~_GEN_2420 & _GEN_82239 : ~_GEN_2006 & _GEN_82239);
    if (_stq_bits_data_bits_T_2 & _GEN_1721) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_9_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_9_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_9_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1626) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_9_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_9_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_9_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_9_bits_committed <= ~_GEN_2452 & (commit_store_3 ? _GEN_2356 | _GEN_2292 | _GEN_137959 : _GEN_2292 | _GEN_137959);
    stq_9_bits_succeeded <= ~_GEN_2452 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h9 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h9 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h9)) & _GEN_1437 & _GEN_1373 & _GEN_1341 & _GEN_1277 & stq_9_bits_succeeded);
    stq_10_valid <= ~_GEN_2489 & (clear_store ? ~_GEN_2421 & _GEN_52426 : ~_GEN_2007 & _GEN_52426);
    stq_10_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hA | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hA | (_GEN_1438 ? (_GEN_1374 ? (_GEN_1342 ? (_GEN_1278 ? stq_10_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_10_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1438 ? (_GEN_1374 ? (_GEN_1342 ? (_GEN_1278 ? stq_10_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_10_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1438 ? (_GEN_1374 ? (_GEN_1342 ? (_GEN_1278 ? stq_10_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_10_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1438 ? (_GEN_1374 ? (_GEN_1342 ? (_GEN_1278 ? stq_10_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_10_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1438 ? (_GEN_1374 ? (_GEN_1342 ? (_GEN_1278 ? stq_10_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_10_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1438 ? (_GEN_1374 ? (_GEN_1342 ? (_GEN_1278 ? stq_10_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_10_bits_addr_valid <= ~_GEN_2489 & (clear_store ? ~_GEN_2421 & _GEN_82016 : ~_GEN_2007 & _GEN_82016);
    if (_GEN_1690) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_10_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_10_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_10_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_10_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_10_bits_addr_bits <= hella_req_addr;
        else
          stq_10_bits_addr_bits <= 40'h0;
      end
      else
        stq_10_bits_addr_bits <= _GEN_338;
      stq_10_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1595) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_10_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_10_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_10_bits_addr_bits <= _GEN_332;
        else
          stq_10_bits_addr_bits <= 40'h0;
      end
      else
        stq_10_bits_addr_bits <= _GEN_334;
      stq_10_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_10_bits_data_valid <= ~_GEN_2489 & (clear_store ? ~_GEN_2421 & _GEN_82240 : ~_GEN_2007 & _GEN_82240);
    if (_stq_bits_data_bits_T_2 & _GEN_1722) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_10_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_10_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_10_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1627) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_10_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_10_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_10_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_10_bits_committed <= ~_GEN_2453 & (commit_store_3 ? _GEN_2357 | _GEN_2293 | _GEN_137960 : _GEN_2293 | _GEN_137960);
    stq_10_bits_succeeded <= ~_GEN_2453 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hA | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hA | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hA)) & _GEN_1438 & _GEN_1374 & _GEN_1342 & _GEN_1278 & stq_10_bits_succeeded);
    stq_11_valid <= ~_GEN_2490 & (clear_store ? ~_GEN_2422 & _GEN_52427 : ~_GEN_2008 & _GEN_52427);
    stq_11_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hB | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hB | (_GEN_1439 ? (_GEN_1375 ? (_GEN_1343 ? (_GEN_1279 ? stq_11_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_11_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1439 ? (_GEN_1375 ? (_GEN_1343 ? (_GEN_1279 ? stq_11_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_11_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1439 ? (_GEN_1375 ? (_GEN_1343 ? (_GEN_1279 ? stq_11_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_11_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1439 ? (_GEN_1375 ? (_GEN_1343 ? (_GEN_1279 ? stq_11_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_11_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1439 ? (_GEN_1375 ? (_GEN_1343 ? (_GEN_1279 ? stq_11_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_11_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1439 ? (_GEN_1375 ? (_GEN_1343 ? (_GEN_1279 ? stq_11_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_11_bits_addr_valid <= ~_GEN_2490 & (clear_store ? ~_GEN_2422 & _GEN_82017 : ~_GEN_2008 & _GEN_82017);
    if (_GEN_1691) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_11_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_11_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_11_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_11_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_11_bits_addr_bits <= hella_req_addr;
        else
          stq_11_bits_addr_bits <= 40'h0;
      end
      else
        stq_11_bits_addr_bits <= _GEN_338;
      stq_11_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1596) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_11_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_11_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_11_bits_addr_bits <= _GEN_332;
        else
          stq_11_bits_addr_bits <= 40'h0;
      end
      else
        stq_11_bits_addr_bits <= _GEN_334;
      stq_11_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_11_bits_data_valid <= ~_GEN_2490 & (clear_store ? ~_GEN_2422 & _GEN_82241 : ~_GEN_2008 & _GEN_82241);
    if (_stq_bits_data_bits_T_2 & _GEN_1723) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_11_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_11_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_11_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1628) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_11_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_11_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_11_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_11_bits_committed <= ~_GEN_2454 & (commit_store_3 ? _GEN_2358 | _GEN_2294 | _GEN_137961 : _GEN_2294 | _GEN_137961);
    stq_11_bits_succeeded <= ~_GEN_2454 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hB | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hB | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hB)) & _GEN_1439 & _GEN_1375 & _GEN_1343 & _GEN_1279 & stq_11_bits_succeeded);
    stq_12_valid <= ~_GEN_2491 & (clear_store ? ~_GEN_2423 & _GEN_52428 : ~_GEN_2009 & _GEN_52428);
    stq_12_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hC | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hC | (_GEN_1440 ? (_GEN_1376 ? (_GEN_1344 ? (_GEN_1280 ? stq_12_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_12_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1440 ? (_GEN_1376 ? (_GEN_1344 ? (_GEN_1280 ? stq_12_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_12_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1440 ? (_GEN_1376 ? (_GEN_1344 ? (_GEN_1280 ? stq_12_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_12_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1440 ? (_GEN_1376 ? (_GEN_1344 ? (_GEN_1280 ? stq_12_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_12_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1440 ? (_GEN_1376 ? (_GEN_1344 ? (_GEN_1280 ? stq_12_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_12_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1440 ? (_GEN_1376 ? (_GEN_1344 ? (_GEN_1280 ? stq_12_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_12_bits_addr_valid <= ~_GEN_2491 & (clear_store ? ~_GEN_2423 & _GEN_82018 : ~_GEN_2009 & _GEN_82018);
    if (_GEN_1692) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_12_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_12_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_12_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_12_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_12_bits_addr_bits <= hella_req_addr;
        else
          stq_12_bits_addr_bits <= 40'h0;
      end
      else
        stq_12_bits_addr_bits <= _GEN_338;
      stq_12_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1597) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_12_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_12_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_12_bits_addr_bits <= _GEN_332;
        else
          stq_12_bits_addr_bits <= 40'h0;
      end
      else
        stq_12_bits_addr_bits <= _GEN_334;
      stq_12_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_12_bits_data_valid <= ~_GEN_2491 & (clear_store ? ~_GEN_2423 & _GEN_82242 : ~_GEN_2009 & _GEN_82242);
    if (_stq_bits_data_bits_T_2 & _GEN_1724) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_12_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_12_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_12_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1629) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_12_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_12_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_12_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_12_bits_committed <= ~_GEN_2455 & (commit_store_3 ? _GEN_2359 | _GEN_2295 | _GEN_137962 : _GEN_2295 | _GEN_137962);
    stq_12_bits_succeeded <= ~_GEN_2455 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hC | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hC | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hC)) & _GEN_1440 & _GEN_1376 & _GEN_1344 & _GEN_1280 & stq_12_bits_succeeded);
    stq_13_valid <= ~_GEN_2492 & (clear_store ? ~_GEN_2424 & _GEN_52429 : ~_GEN_2010 & _GEN_52429);
    stq_13_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hD | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hD | (_GEN_1441 ? (_GEN_1377 ? (_GEN_1345 ? (_GEN_1281 ? stq_13_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_13_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1441 ? (_GEN_1377 ? (_GEN_1345 ? (_GEN_1281 ? stq_13_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_13_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1441 ? (_GEN_1377 ? (_GEN_1345 ? (_GEN_1281 ? stq_13_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_13_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1441 ? (_GEN_1377 ? (_GEN_1345 ? (_GEN_1281 ? stq_13_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_13_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1441 ? (_GEN_1377 ? (_GEN_1345 ? (_GEN_1281 ? stq_13_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_13_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1441 ? (_GEN_1377 ? (_GEN_1345 ? (_GEN_1281 ? stq_13_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_13_bits_addr_valid <= ~_GEN_2492 & (clear_store ? ~_GEN_2424 & _GEN_82019 : ~_GEN_2010 & _GEN_82019);
    if (_GEN_1693) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_13_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_13_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_13_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_13_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_13_bits_addr_bits <= hella_req_addr;
        else
          stq_13_bits_addr_bits <= 40'h0;
      end
      else
        stq_13_bits_addr_bits <= _GEN_338;
      stq_13_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1598) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_13_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_13_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_13_bits_addr_bits <= _GEN_332;
        else
          stq_13_bits_addr_bits <= 40'h0;
      end
      else
        stq_13_bits_addr_bits <= _GEN_334;
      stq_13_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_13_bits_data_valid <= ~_GEN_2492 & (clear_store ? ~_GEN_2424 & _GEN_82243 : ~_GEN_2010 & _GEN_82243);
    if (_stq_bits_data_bits_T_2 & _GEN_1725) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_13_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_13_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_13_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1630) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_13_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_13_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_13_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_13_bits_committed <= ~_GEN_2456 & (commit_store_3 ? _GEN_2360 | _GEN_2296 | _GEN_137963 : _GEN_2296 | _GEN_137963);
    stq_13_bits_succeeded <= ~_GEN_2456 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hD | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hD | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hD)) & _GEN_1441 & _GEN_1377 & _GEN_1345 & _GEN_1281 & stq_13_bits_succeeded);
    stq_14_valid <= ~_GEN_2493 & (clear_store ? ~_GEN_2425 & _GEN_52430 : ~_GEN_2011 & _GEN_52430);
    stq_14_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hE | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hE | (_GEN_1442 ? (_GEN_1378 ? (_GEN_1346 ? (_GEN_1282 ? stq_14_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_14_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1442 ? (_GEN_1378 ? (_GEN_1346 ? (_GEN_1282 ? stq_14_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_14_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1442 ? (_GEN_1378 ? (_GEN_1346 ? (_GEN_1282 ? stq_14_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_14_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1442 ? (_GEN_1378 ? (_GEN_1346 ? (_GEN_1282 ? stq_14_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_14_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1442 ? (_GEN_1378 ? (_GEN_1346 ? (_GEN_1282 ? stq_14_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_14_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1442 ? (_GEN_1378 ? (_GEN_1346 ? (_GEN_1282 ? stq_14_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_14_bits_addr_valid <= ~_GEN_2493 & (clear_store ? ~_GEN_2425 & _GEN_82020 : ~_GEN_2011 & _GEN_82020);
    if (_GEN_1694) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_14_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_14_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_14_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_14_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_14_bits_addr_bits <= hella_req_addr;
        else
          stq_14_bits_addr_bits <= 40'h0;
      end
      else
        stq_14_bits_addr_bits <= _GEN_338;
      stq_14_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1599) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_14_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_14_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_14_bits_addr_bits <= _GEN_332;
        else
          stq_14_bits_addr_bits <= 40'h0;
      end
      else
        stq_14_bits_addr_bits <= _GEN_334;
      stq_14_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_14_bits_data_valid <= ~_GEN_2493 & (clear_store ? ~_GEN_2425 & _GEN_82244 : ~_GEN_2011 & _GEN_82244);
    if (_stq_bits_data_bits_T_2 & _GEN_1726) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_14_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_14_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_14_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1631) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_14_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_14_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_14_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_14_bits_committed <= ~_GEN_2457 & (commit_store_3 ? _GEN_2361 | _GEN_2297 | _GEN_137964 : _GEN_2297 | _GEN_137964);
    stq_14_bits_succeeded <= ~_GEN_2457 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hE | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hE | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hE)) & _GEN_1442 & _GEN_1378 & _GEN_1346 & _GEN_1282 & stq_14_bits_succeeded);
    stq_15_valid <= ~_GEN_2494 & (clear_store ? ~_GEN_2426 & _GEN_52431 : ~_GEN_2012 & _GEN_52431);
    stq_15_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'hF | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'hF | (_GEN_1443 ? (_GEN_1379 ? (_GEN_1347 ? (_GEN_1283 ? stq_15_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_15_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1443 ? (_GEN_1379 ? (_GEN_1347 ? (_GEN_1283 ? stq_15_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_15_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1443 ? (_GEN_1379 ? (_GEN_1347 ? (_GEN_1283 ? stq_15_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_15_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1443 ? (_GEN_1379 ? (_GEN_1347 ? (_GEN_1283 ? stq_15_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_15_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1443 ? (_GEN_1379 ? (_GEN_1347 ? (_GEN_1283 ? stq_15_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_15_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1443 ? (_GEN_1379 ? (_GEN_1347 ? (_GEN_1283 ? stq_15_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_15_bits_addr_valid <= ~_GEN_2494 & (clear_store ? ~_GEN_2426 & _GEN_82021 : ~_GEN_2012 & _GEN_82021);
    if (_GEN_1695) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_15_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_15_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_15_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_15_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_15_bits_addr_bits <= hella_req_addr;
        else
          stq_15_bits_addr_bits <= 40'h0;
      end
      else
        stq_15_bits_addr_bits <= _GEN_338;
      stq_15_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1600) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_15_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_15_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_15_bits_addr_bits <= _GEN_332;
        else
          stq_15_bits_addr_bits <= 40'h0;
      end
      else
        stq_15_bits_addr_bits <= _GEN_334;
      stq_15_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_15_bits_data_valid <= ~_GEN_2494 & (clear_store ? ~_GEN_2426 & _GEN_82245 : ~_GEN_2012 & _GEN_82245);
    if (_stq_bits_data_bits_T_2 & _GEN_1727) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_15_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_15_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_15_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1632) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_15_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_15_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_15_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_15_bits_committed <= ~_GEN_2458 & (commit_store_3 ? _GEN_2362 | _GEN_2298 | _GEN_137965 : _GEN_2298 | _GEN_137965);
    stq_15_bits_succeeded <= ~_GEN_2458 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'hF | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'hF | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'hF)) & _GEN_1443 & _GEN_1379 & _GEN_1347 & _GEN_1283 & stq_15_bits_succeeded);
    stq_16_valid <= ~_GEN_2495 & (clear_store ? ~_GEN_2427 & _GEN_52432 : ~_GEN_2013 & _GEN_52432);
    stq_16_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h10 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h10 | (_GEN_1444 ? (_GEN_1380 ? (_GEN_1348 ? (_GEN_1284 ? stq_16_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_16_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1444 ? (_GEN_1380 ? (_GEN_1348 ? (_GEN_1284 ? stq_16_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_16_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1444 ? (_GEN_1380 ? (_GEN_1348 ? (_GEN_1284 ? stq_16_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_16_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1444 ? (_GEN_1380 ? (_GEN_1348 ? (_GEN_1284 ? stq_16_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_16_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1444 ? (_GEN_1380 ? (_GEN_1348 ? (_GEN_1284 ? stq_16_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_16_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1444 ? (_GEN_1380 ? (_GEN_1348 ? (_GEN_1284 ? stq_16_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_16_bits_addr_valid <= ~_GEN_2495 & (clear_store ? ~_GEN_2427 & _GEN_82022 : ~_GEN_2013 & _GEN_82022);
    if (_GEN_1696) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_16_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_16_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_16_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_16_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_16_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_16_bits_addr_bits <= hella_req_addr;
        else
          stq_16_bits_addr_bits <= 40'h0;
      end
      else
        stq_16_bits_addr_bits <= _GEN_338;
      stq_16_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1601) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_16_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_16_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_16_bits_addr_bits <= _GEN_332;
        else
          stq_16_bits_addr_bits <= 40'h0;
      end
      else
        stq_16_bits_addr_bits <= _GEN_334;
      stq_16_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_16_bits_data_valid <= ~_GEN_2495 & (clear_store ? ~_GEN_2427 & _GEN_82246 : ~_GEN_2013 & _GEN_82246);
    if (_stq_bits_data_bits_T_2 & _GEN_1728) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_16_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_16_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_16_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1633) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_16_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_16_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_16_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_16_bits_committed <= ~_GEN_2459 & (commit_store_3 ? _GEN_2363 | _GEN_2299 | _GEN_137966 : _GEN_2299 | _GEN_137966);
    stq_16_bits_succeeded <= ~_GEN_2459 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h10 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h10 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h10)) & _GEN_1444 & _GEN_1380 & _GEN_1348 & _GEN_1284 & stq_16_bits_succeeded);
    stq_17_valid <= ~_GEN_2496 & (clear_store ? ~_GEN_2428 & _GEN_52433 : ~_GEN_2014 & _GEN_52433);
    stq_17_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h11 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h11 | (_GEN_1445 ? (_GEN_1381 ? (_GEN_1349 ? (_GEN_1285 ? stq_17_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_17_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1445 ? (_GEN_1381 ? (_GEN_1349 ? (_GEN_1285 ? stq_17_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_17_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1445 ? (_GEN_1381 ? (_GEN_1349 ? (_GEN_1285 ? stq_17_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_17_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1445 ? (_GEN_1381 ? (_GEN_1349 ? (_GEN_1285 ? stq_17_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_17_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1445 ? (_GEN_1381 ? (_GEN_1349 ? (_GEN_1285 ? stq_17_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_17_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1445 ? (_GEN_1381 ? (_GEN_1349 ? (_GEN_1285 ? stq_17_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_17_bits_addr_valid <= ~_GEN_2496 & (clear_store ? ~_GEN_2428 & _GEN_82023 : ~_GEN_2014 & _GEN_82023);
    if (_GEN_1697) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_17_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_17_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_17_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_17_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_17_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_17_bits_addr_bits <= hella_req_addr;
        else
          stq_17_bits_addr_bits <= 40'h0;
      end
      else
        stq_17_bits_addr_bits <= _GEN_338;
      stq_17_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1602) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_17_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_17_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_17_bits_addr_bits <= _GEN_332;
        else
          stq_17_bits_addr_bits <= 40'h0;
      end
      else
        stq_17_bits_addr_bits <= _GEN_334;
      stq_17_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_17_bits_data_valid <= ~_GEN_2496 & (clear_store ? ~_GEN_2428 & _GEN_82247 : ~_GEN_2014 & _GEN_82247);
    if (_stq_bits_data_bits_T_2 & _GEN_1729) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_17_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_17_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_17_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1634) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_17_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_17_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_17_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_17_bits_committed <= ~_GEN_2460 & (commit_store_3 ? _GEN_2364 | _GEN_2300 | _GEN_137967 : _GEN_2300 | _GEN_137967);
    stq_17_bits_succeeded <= ~_GEN_2460 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h11 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h11 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h11)) & _GEN_1445 & _GEN_1381 & _GEN_1349 & _GEN_1285 & stq_17_bits_succeeded);
    stq_18_valid <= ~_GEN_2497 & (clear_store ? ~_GEN_2429 & _GEN_52434 : ~_GEN_2015 & _GEN_52434);
    stq_18_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h12 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h12 | (_GEN_1446 ? (_GEN_1382 ? (_GEN_1350 ? (_GEN_1286 ? stq_18_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_18_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1446 ? (_GEN_1382 ? (_GEN_1350 ? (_GEN_1286 ? stq_18_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_18_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1446 ? (_GEN_1382 ? (_GEN_1350 ? (_GEN_1286 ? stq_18_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_18_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1446 ? (_GEN_1382 ? (_GEN_1350 ? (_GEN_1286 ? stq_18_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_18_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1446 ? (_GEN_1382 ? (_GEN_1350 ? (_GEN_1286 ? stq_18_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_18_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1446 ? (_GEN_1382 ? (_GEN_1350 ? (_GEN_1286 ? stq_18_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_18_bits_addr_valid <= ~_GEN_2497 & (clear_store ? ~_GEN_2429 & _GEN_82024 : ~_GEN_2015 & _GEN_82024);
    if (_GEN_1698) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_18_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_18_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_18_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_18_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_18_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_18_bits_addr_bits <= hella_req_addr;
        else
          stq_18_bits_addr_bits <= 40'h0;
      end
      else
        stq_18_bits_addr_bits <= _GEN_338;
      stq_18_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1603) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_18_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_18_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_18_bits_addr_bits <= _GEN_332;
        else
          stq_18_bits_addr_bits <= 40'h0;
      end
      else
        stq_18_bits_addr_bits <= _GEN_334;
      stq_18_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_18_bits_data_valid <= ~_GEN_2497 & (clear_store ? ~_GEN_2429 & _GEN_82248 : ~_GEN_2015 & _GEN_82248);
    if (_stq_bits_data_bits_T_2 & _GEN_1730) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_18_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_18_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_18_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1635) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_18_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_18_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_18_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_18_bits_committed <= ~_GEN_2461 & (commit_store_3 ? _GEN_2365 | _GEN_2301 | _GEN_137968 : _GEN_2301 | _GEN_137968);
    stq_18_bits_succeeded <= ~_GEN_2461 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h12 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h12 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h12)) & _GEN_1446 & _GEN_1382 & _GEN_1350 & _GEN_1286 & stq_18_bits_succeeded);
    stq_19_valid <= ~_GEN_2498 & (clear_store ? ~_GEN_2430 & _GEN_52435 : ~_GEN_2016 & _GEN_52435);
    stq_19_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h13 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h13 | (_GEN_1447 ? (_GEN_1383 ? (_GEN_1351 ? (_GEN_1287 ? stq_19_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_19_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1447 ? (_GEN_1383 ? (_GEN_1351 ? (_GEN_1287 ? stq_19_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_19_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1447 ? (_GEN_1383 ? (_GEN_1351 ? (_GEN_1287 ? stq_19_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_19_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1447 ? (_GEN_1383 ? (_GEN_1351 ? (_GEN_1287 ? stq_19_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_19_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1447 ? (_GEN_1383 ? (_GEN_1351 ? (_GEN_1287 ? stq_19_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_19_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1447 ? (_GEN_1383 ? (_GEN_1351 ? (_GEN_1287 ? stq_19_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_19_bits_addr_valid <= ~_GEN_2498 & (clear_store ? ~_GEN_2430 & _GEN_82025 : ~_GEN_2016 & _GEN_82025);
    if (_GEN_1699) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_19_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_19_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_19_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_19_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_19_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_19_bits_addr_bits <= hella_req_addr;
        else
          stq_19_bits_addr_bits <= 40'h0;
      end
      else
        stq_19_bits_addr_bits <= _GEN_338;
      stq_19_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1604) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_19_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_19_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_19_bits_addr_bits <= _GEN_332;
        else
          stq_19_bits_addr_bits <= 40'h0;
      end
      else
        stq_19_bits_addr_bits <= _GEN_334;
      stq_19_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_19_bits_data_valid <= ~_GEN_2498 & (clear_store ? ~_GEN_2430 & _GEN_82249 : ~_GEN_2016 & _GEN_82249);
    if (_stq_bits_data_bits_T_2 & _GEN_1731) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_19_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_19_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_19_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1636) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_19_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_19_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_19_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_19_bits_committed <= ~_GEN_2462 & (commit_store_3 ? _GEN_2366 | _GEN_2302 | _GEN_137969 : _GEN_2302 | _GEN_137969);
    stq_19_bits_succeeded <= ~_GEN_2462 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h13 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h13 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h13)) & _GEN_1447 & _GEN_1383 & _GEN_1351 & _GEN_1287 & stq_19_bits_succeeded);
    stq_20_valid <= ~_GEN_2499 & (clear_store ? ~_GEN_2431 & _GEN_52436 : ~_GEN_2017 & _GEN_52436);
    stq_20_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h14 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h14 | (_GEN_1448 ? (_GEN_1384 ? (_GEN_1352 ? (_GEN_1288 ? stq_20_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_20_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1448 ? (_GEN_1384 ? (_GEN_1352 ? (_GEN_1288 ? stq_20_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_20_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1448 ? (_GEN_1384 ? (_GEN_1352 ? (_GEN_1288 ? stq_20_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_20_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1448 ? (_GEN_1384 ? (_GEN_1352 ? (_GEN_1288 ? stq_20_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_20_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1448 ? (_GEN_1384 ? (_GEN_1352 ? (_GEN_1288 ? stq_20_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_20_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1448 ? (_GEN_1384 ? (_GEN_1352 ? (_GEN_1288 ? stq_20_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_20_bits_addr_valid <= ~_GEN_2499 & (clear_store ? ~_GEN_2431 & _GEN_82026 : ~_GEN_2017 & _GEN_82026);
    if (_GEN_1700) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_20_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_20_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_20_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_20_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_20_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_20_bits_addr_bits <= hella_req_addr;
        else
          stq_20_bits_addr_bits <= 40'h0;
      end
      else
        stq_20_bits_addr_bits <= _GEN_338;
      stq_20_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1605) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_20_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_20_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_20_bits_addr_bits <= _GEN_332;
        else
          stq_20_bits_addr_bits <= 40'h0;
      end
      else
        stq_20_bits_addr_bits <= _GEN_334;
      stq_20_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_20_bits_data_valid <= ~_GEN_2499 & (clear_store ? ~_GEN_2431 & _GEN_82250 : ~_GEN_2017 & _GEN_82250);
    if (_stq_bits_data_bits_T_2 & _GEN_1732) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_20_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_20_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_20_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1637) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_20_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_20_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_20_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_20_bits_committed <= ~_GEN_2463 & (commit_store_3 ? _GEN_2367 | _GEN_2303 | _GEN_137970 : _GEN_2303 | _GEN_137970);
    stq_20_bits_succeeded <= ~_GEN_2463 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h14 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h14 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h14)) & _GEN_1448 & _GEN_1384 & _GEN_1352 & _GEN_1288 & stq_20_bits_succeeded);
    stq_21_valid <= ~_GEN_2500 & (clear_store ? ~_GEN_2432 & _GEN_52437 : ~_GEN_2018 & _GEN_52437);
    stq_21_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h15 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h15 | (_GEN_1449 ? (_GEN_1385 ? (_GEN_1353 ? (_GEN_1289 ? stq_21_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_21_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1449 ? (_GEN_1385 ? (_GEN_1353 ? (_GEN_1289 ? stq_21_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_21_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1449 ? (_GEN_1385 ? (_GEN_1353 ? (_GEN_1289 ? stq_21_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_21_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1449 ? (_GEN_1385 ? (_GEN_1353 ? (_GEN_1289 ? stq_21_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_21_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1449 ? (_GEN_1385 ? (_GEN_1353 ? (_GEN_1289 ? stq_21_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_21_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1449 ? (_GEN_1385 ? (_GEN_1353 ? (_GEN_1289 ? stq_21_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_21_bits_addr_valid <= ~_GEN_2500 & (clear_store ? ~_GEN_2432 & _GEN_82027 : ~_GEN_2018 & _GEN_82027);
    if (_GEN_1701) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_21_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_21_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_21_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_21_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_21_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_21_bits_addr_bits <= hella_req_addr;
        else
          stq_21_bits_addr_bits <= 40'h0;
      end
      else
        stq_21_bits_addr_bits <= _GEN_338;
      stq_21_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1606) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_21_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_21_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_21_bits_addr_bits <= _GEN_332;
        else
          stq_21_bits_addr_bits <= 40'h0;
      end
      else
        stq_21_bits_addr_bits <= _GEN_334;
      stq_21_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_21_bits_data_valid <= ~_GEN_2500 & (clear_store ? ~_GEN_2432 & _GEN_82251 : ~_GEN_2018 & _GEN_82251);
    if (_stq_bits_data_bits_T_2 & _GEN_1733) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_21_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_21_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_21_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1638) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_21_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_21_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_21_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_21_bits_committed <= ~_GEN_2464 & (commit_store_3 ? _GEN_2368 | _GEN_2304 | _GEN_137971 : _GEN_2304 | _GEN_137971);
    stq_21_bits_succeeded <= ~_GEN_2464 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h15 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h15 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h15)) & _GEN_1449 & _GEN_1385 & _GEN_1353 & _GEN_1289 & stq_21_bits_succeeded);
    stq_22_valid <= ~_GEN_2501 & (clear_store ? ~_GEN_2433 & _GEN_52438 : ~_GEN_2019 & _GEN_52438);
    stq_22_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h16 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h16 | (_GEN_1450 ? (_GEN_1386 ? (_GEN_1354 ? (_GEN_1290 ? stq_22_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_22_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1450 ? (_GEN_1386 ? (_GEN_1354 ? (_GEN_1290 ? stq_22_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_22_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1450 ? (_GEN_1386 ? (_GEN_1354 ? (_GEN_1290 ? stq_22_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_22_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1450 ? (_GEN_1386 ? (_GEN_1354 ? (_GEN_1290 ? stq_22_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_22_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1450 ? (_GEN_1386 ? (_GEN_1354 ? (_GEN_1290 ? stq_22_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_22_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1450 ? (_GEN_1386 ? (_GEN_1354 ? (_GEN_1290 ? stq_22_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_22_bits_addr_valid <= ~_GEN_2501 & (clear_store ? ~_GEN_2433 & _GEN_82028 : ~_GEN_2019 & _GEN_82028);
    if (_GEN_1702) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_22_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_22_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_22_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_22_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_22_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_22_bits_addr_bits <= hella_req_addr;
        else
          stq_22_bits_addr_bits <= 40'h0;
      end
      else
        stq_22_bits_addr_bits <= _GEN_338;
      stq_22_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1607) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_22_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_22_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_22_bits_addr_bits <= _GEN_332;
        else
          stq_22_bits_addr_bits <= 40'h0;
      end
      else
        stq_22_bits_addr_bits <= _GEN_334;
      stq_22_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_22_bits_data_valid <= ~_GEN_2501 & (clear_store ? ~_GEN_2433 & _GEN_82252 : ~_GEN_2019 & _GEN_82252);
    if (_stq_bits_data_bits_T_2 & _GEN_1734) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_22_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_22_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_22_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1639) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_22_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_22_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_22_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_22_bits_committed <= ~_GEN_2465 & (commit_store_3 ? _GEN_2369 | _GEN_2305 | _GEN_137972 : _GEN_2305 | _GEN_137972);
    stq_22_bits_succeeded <= ~_GEN_2465 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h16 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h16 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h16)) & _GEN_1450 & _GEN_1386 & _GEN_1354 & _GEN_1290 & stq_22_bits_succeeded);
    stq_23_valid <= ~_GEN_2502 & (clear_store ? ~_GEN_2434 & _GEN_52439 : ~_GEN_2020 & _GEN_52439);
    stq_23_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h17 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h17 | (_GEN_1451 ? (_GEN_1387 ? (_GEN_1355 ? (_GEN_1291 ? stq_23_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_23_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1451 ? (_GEN_1387 ? (_GEN_1355 ? (_GEN_1291 ? stq_23_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_23_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1451 ? (_GEN_1387 ? (_GEN_1355 ? (_GEN_1291 ? stq_23_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_23_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1451 ? (_GEN_1387 ? (_GEN_1355 ? (_GEN_1291 ? stq_23_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_23_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1451 ? (_GEN_1387 ? (_GEN_1355 ? (_GEN_1291 ? stq_23_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_23_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1451 ? (_GEN_1387 ? (_GEN_1355 ? (_GEN_1291 ? stq_23_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_23_bits_addr_valid <= ~_GEN_2502 & (clear_store ? ~_GEN_2434 & _GEN_82029 : ~_GEN_2020 & _GEN_82029);
    if (_GEN_1703) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_23_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_23_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_23_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_23_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_23_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_23_bits_addr_bits <= hella_req_addr;
        else
          stq_23_bits_addr_bits <= 40'h0;
      end
      else
        stq_23_bits_addr_bits <= _GEN_338;
      stq_23_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1608) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_23_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_23_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_23_bits_addr_bits <= _GEN_332;
        else
          stq_23_bits_addr_bits <= 40'h0;
      end
      else
        stq_23_bits_addr_bits <= _GEN_334;
      stq_23_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_23_bits_data_valid <= ~_GEN_2502 & (clear_store ? ~_GEN_2434 & _GEN_82253 : ~_GEN_2020 & _GEN_82253);
    if (_stq_bits_data_bits_T_2 & _GEN_1735) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_23_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_23_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_23_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1640) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_23_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_23_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_23_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_23_bits_committed <= ~_GEN_2466 & (commit_store_3 ? _GEN_2370 | _GEN_2306 | _GEN_137973 : _GEN_2306 | _GEN_137973);
    stq_23_bits_succeeded <= ~_GEN_2466 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h17 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h17 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h17)) & _GEN_1451 & _GEN_1387 & _GEN_1355 & _GEN_1291 & stq_23_bits_succeeded);
    stq_24_valid <= ~_GEN_2503 & (clear_store ? ~_GEN_2435 & _GEN_52440 : ~_GEN_2021 & _GEN_52440);
    stq_24_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h18 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h18 | (_GEN_1452 ? (_GEN_1388 ? (_GEN_1356 ? (_GEN_1292 ? stq_24_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_24_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1452 ? (_GEN_1388 ? (_GEN_1356 ? (_GEN_1292 ? stq_24_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_24_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1452 ? (_GEN_1388 ? (_GEN_1356 ? (_GEN_1292 ? stq_24_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_24_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1452 ? (_GEN_1388 ? (_GEN_1356 ? (_GEN_1292 ? stq_24_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_24_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1452 ? (_GEN_1388 ? (_GEN_1356 ? (_GEN_1292 ? stq_24_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_24_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1452 ? (_GEN_1388 ? (_GEN_1356 ? (_GEN_1292 ? stq_24_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_24_bits_addr_valid <= ~_GEN_2503 & (clear_store ? ~_GEN_2435 & _GEN_82030 : ~_GEN_2021 & _GEN_82030);
    if (_GEN_1704) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_24_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_24_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_24_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_24_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_24_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_24_bits_addr_bits <= hella_req_addr;
        else
          stq_24_bits_addr_bits <= 40'h0;
      end
      else
        stq_24_bits_addr_bits <= _GEN_338;
      stq_24_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1609) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_24_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_24_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_24_bits_addr_bits <= _GEN_332;
        else
          stq_24_bits_addr_bits <= 40'h0;
      end
      else
        stq_24_bits_addr_bits <= _GEN_334;
      stq_24_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_24_bits_data_valid <= ~_GEN_2503 & (clear_store ? ~_GEN_2435 & _GEN_82254 : ~_GEN_2021 & _GEN_82254);
    if (_stq_bits_data_bits_T_2 & _GEN_1736) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_24_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_24_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_24_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1641) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_24_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_24_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_24_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_24_bits_committed <= ~_GEN_2467 & (commit_store_3 ? _GEN_2371 | _GEN_2307 | _GEN_137974 : _GEN_2307 | _GEN_137974);
    stq_24_bits_succeeded <= ~_GEN_2467 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h18 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h18 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h18)) & _GEN_1452 & _GEN_1388 & _GEN_1356 & _GEN_1292 & stq_24_bits_succeeded);
    stq_25_valid <= ~_GEN_2504 & (clear_store ? ~_GEN_2436 & _GEN_52441 : ~_GEN_2022 & _GEN_52441);
    stq_25_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h19 | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h19 | (_GEN_1453 ? (_GEN_1389 ? (_GEN_1357 ? (_GEN_1293 ? stq_25_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_25_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1453 ? (_GEN_1389 ? (_GEN_1357 ? (_GEN_1293 ? stq_25_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_25_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1453 ? (_GEN_1389 ? (_GEN_1357 ? (_GEN_1293 ? stq_25_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_25_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1453 ? (_GEN_1389 ? (_GEN_1357 ? (_GEN_1293 ? stq_25_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_25_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1453 ? (_GEN_1389 ? (_GEN_1357 ? (_GEN_1293 ? stq_25_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_25_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1453 ? (_GEN_1389 ? (_GEN_1357 ? (_GEN_1293 ? stq_25_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_25_bits_addr_valid <= ~_GEN_2504 & (clear_store ? ~_GEN_2436 & _GEN_82031 : ~_GEN_2022 & _GEN_82031);
    if (_GEN_1705) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_25_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_25_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_25_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_25_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_25_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_25_bits_addr_bits <= hella_req_addr;
        else
          stq_25_bits_addr_bits <= 40'h0;
      end
      else
        stq_25_bits_addr_bits <= _GEN_338;
      stq_25_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1610) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_25_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_25_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_25_bits_addr_bits <= _GEN_332;
        else
          stq_25_bits_addr_bits <= 40'h0;
      end
      else
        stq_25_bits_addr_bits <= _GEN_334;
      stq_25_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_25_bits_data_valid <= ~_GEN_2504 & (clear_store ? ~_GEN_2436 & _GEN_82255 : ~_GEN_2022 & _GEN_82255);
    if (_stq_bits_data_bits_T_2 & _GEN_1737) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_25_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_25_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_25_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1642) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_25_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_25_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_25_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_25_bits_committed <= ~_GEN_2468 & (commit_store_3 ? _GEN_2372 | _GEN_2308 | _GEN_137975 : _GEN_2308 | _GEN_137975);
    stq_25_bits_succeeded <= ~_GEN_2468 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h19 | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h19 | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h19)) & _GEN_1453 & _GEN_1389 & _GEN_1357 & _GEN_1293 & stq_25_bits_succeeded);
    stq_26_valid <= ~_GEN_2505 & (clear_store ? ~_GEN_2437 & _GEN_52442 : ~_GEN_2023 & _GEN_52442);
    stq_26_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1A | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1A | (_GEN_1454 ? (_GEN_1390 ? (_GEN_1358 ? (_GEN_1294 ? stq_26_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_26_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1454 ? (_GEN_1390 ? (_GEN_1358 ? (_GEN_1294 ? stq_26_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_26_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1454 ? (_GEN_1390 ? (_GEN_1358 ? (_GEN_1294 ? stq_26_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_26_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1454 ? (_GEN_1390 ? (_GEN_1358 ? (_GEN_1294 ? stq_26_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_26_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1454 ? (_GEN_1390 ? (_GEN_1358 ? (_GEN_1294 ? stq_26_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_26_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1454 ? (_GEN_1390 ? (_GEN_1358 ? (_GEN_1294 ? stq_26_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_26_bits_addr_valid <= ~_GEN_2505 & (clear_store ? ~_GEN_2437 & _GEN_82032 : ~_GEN_2023 & _GEN_82032);
    if (_GEN_1706) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_26_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_26_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_26_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_26_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_26_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_26_bits_addr_bits <= hella_req_addr;
        else
          stq_26_bits_addr_bits <= 40'h0;
      end
      else
        stq_26_bits_addr_bits <= _GEN_338;
      stq_26_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1611) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_26_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_26_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_26_bits_addr_bits <= _GEN_332;
        else
          stq_26_bits_addr_bits <= 40'h0;
      end
      else
        stq_26_bits_addr_bits <= _GEN_334;
      stq_26_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_26_bits_data_valid <= ~_GEN_2505 & (clear_store ? ~_GEN_2437 & _GEN_82256 : ~_GEN_2023 & _GEN_82256);
    if (_stq_bits_data_bits_T_2 & _GEN_1738) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_26_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_26_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_26_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1643) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_26_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_26_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_26_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_26_bits_committed <= ~_GEN_2469 & (commit_store_3 ? _GEN_2373 | _GEN_2309 | _GEN_137976 : _GEN_2309 | _GEN_137976);
    stq_26_bits_succeeded <= ~_GEN_2469 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1A | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1A | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h1A)) & _GEN_1454 & _GEN_1390 & _GEN_1358 & _GEN_1294 & stq_26_bits_succeeded);
    stq_27_valid <= ~_GEN_2506 & (clear_store ? ~_GEN_2438 & _GEN_52443 : ~_GEN_2024 & _GEN_52443);
    stq_27_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1B | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1B | (_GEN_1455 ? (_GEN_1391 ? (_GEN_1359 ? (_GEN_1295 ? stq_27_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_27_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1455 ? (_GEN_1391 ? (_GEN_1359 ? (_GEN_1295 ? stq_27_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_27_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1455 ? (_GEN_1391 ? (_GEN_1359 ? (_GEN_1295 ? stq_27_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_27_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1455 ? (_GEN_1391 ? (_GEN_1359 ? (_GEN_1295 ? stq_27_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_27_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1455 ? (_GEN_1391 ? (_GEN_1359 ? (_GEN_1295 ? stq_27_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_27_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1455 ? (_GEN_1391 ? (_GEN_1359 ? (_GEN_1295 ? stq_27_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_27_bits_addr_valid <= ~_GEN_2506 & (clear_store ? ~_GEN_2438 & _GEN_82033 : ~_GEN_2024 & _GEN_82033);
    if (_GEN_1707) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_27_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_27_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_27_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_27_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_27_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_27_bits_addr_bits <= hella_req_addr;
        else
          stq_27_bits_addr_bits <= 40'h0;
      end
      else
        stq_27_bits_addr_bits <= _GEN_338;
      stq_27_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1612) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_27_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_27_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_27_bits_addr_bits <= _GEN_332;
        else
          stq_27_bits_addr_bits <= 40'h0;
      end
      else
        stq_27_bits_addr_bits <= _GEN_334;
      stq_27_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_27_bits_data_valid <= ~_GEN_2506 & (clear_store ? ~_GEN_2438 & _GEN_82257 : ~_GEN_2024 & _GEN_82257);
    if (_stq_bits_data_bits_T_2 & _GEN_1739) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_27_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_27_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_27_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1644) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_27_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_27_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_27_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_27_bits_committed <= ~_GEN_2470 & (commit_store_3 ? _GEN_2374 | _GEN_2310 | _GEN_137977 : _GEN_2310 | _GEN_137977);
    stq_27_bits_succeeded <= ~_GEN_2470 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1B | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1B | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h1B)) & _GEN_1455 & _GEN_1391 & _GEN_1359 & _GEN_1295 & stq_27_bits_succeeded);
    stq_28_valid <= ~_GEN_2507 & (clear_store ? ~_GEN_2439 & _GEN_52444 : ~_GEN_2025 & _GEN_52444);
    stq_28_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1C | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1C | (_GEN_1456 ? (_GEN_1392 ? (_GEN_1360 ? (_GEN_1296 ? stq_28_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_28_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1456 ? (_GEN_1392 ? (_GEN_1360 ? (_GEN_1296 ? stq_28_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_28_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1456 ? (_GEN_1392 ? (_GEN_1360 ? (_GEN_1296 ? stq_28_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_28_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1456 ? (_GEN_1392 ? (_GEN_1360 ? (_GEN_1296 ? stq_28_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_28_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1456 ? (_GEN_1392 ? (_GEN_1360 ? (_GEN_1296 ? stq_28_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_28_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1456 ? (_GEN_1392 ? (_GEN_1360 ? (_GEN_1296 ? stq_28_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_28_bits_addr_valid <= ~_GEN_2507 & (clear_store ? ~_GEN_2439 & _GEN_82034 : ~_GEN_2025 & _GEN_82034);
    if (_GEN_1708) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_28_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_28_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_28_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_28_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_28_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_28_bits_addr_bits <= hella_req_addr;
        else
          stq_28_bits_addr_bits <= 40'h0;
      end
      else
        stq_28_bits_addr_bits <= _GEN_338;
      stq_28_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1613) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_28_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_28_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_28_bits_addr_bits <= _GEN_332;
        else
          stq_28_bits_addr_bits <= 40'h0;
      end
      else
        stq_28_bits_addr_bits <= _GEN_334;
      stq_28_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_28_bits_data_valid <= ~_GEN_2507 & (clear_store ? ~_GEN_2439 & _GEN_82258 : ~_GEN_2025 & _GEN_82258);
    if (_stq_bits_data_bits_T_2 & _GEN_1740) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_28_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_28_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_28_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1645) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_28_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_28_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_28_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_28_bits_committed <= ~_GEN_2471 & (commit_store_3 ? _GEN_2375 | _GEN_2311 | _GEN_137978 : _GEN_2311 | _GEN_137978);
    stq_28_bits_succeeded <= ~_GEN_2471 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1C | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1C | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h1C)) & _GEN_1456 & _GEN_1392 & _GEN_1360 & _GEN_1296 & stq_28_bits_succeeded);
    stq_29_valid <= ~_GEN_2508 & (clear_store ? ~_GEN_2440 & _GEN_52445 : ~_GEN_2026 & _GEN_52445);
    stq_29_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1D | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1D | (_GEN_1457 ? (_GEN_1393 ? (_GEN_1361 ? (_GEN_1297 ? stq_29_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_29_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1457 ? (_GEN_1393 ? (_GEN_1361 ? (_GEN_1297 ? stq_29_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_29_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1457 ? (_GEN_1393 ? (_GEN_1361 ? (_GEN_1297 ? stq_29_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_29_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1457 ? (_GEN_1393 ? (_GEN_1361 ? (_GEN_1297 ? stq_29_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_29_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1457 ? (_GEN_1393 ? (_GEN_1361 ? (_GEN_1297 ? stq_29_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_29_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1457 ? (_GEN_1393 ? (_GEN_1361 ? (_GEN_1297 ? stq_29_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_29_bits_addr_valid <= ~_GEN_2508 & (clear_store ? ~_GEN_2440 & _GEN_82035 : ~_GEN_2026 & _GEN_82035);
    if (_GEN_1709) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_29_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_29_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_29_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_29_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_29_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_29_bits_addr_bits <= hella_req_addr;
        else
          stq_29_bits_addr_bits <= 40'h0;
      end
      else
        stq_29_bits_addr_bits <= _GEN_338;
      stq_29_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1614) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_29_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_29_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_29_bits_addr_bits <= _GEN_332;
        else
          stq_29_bits_addr_bits <= 40'h0;
      end
      else
        stq_29_bits_addr_bits <= _GEN_334;
      stq_29_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_29_bits_data_valid <= ~_GEN_2508 & (clear_store ? ~_GEN_2440 & _GEN_82259 : ~_GEN_2026 & _GEN_82259);
    if (_stq_bits_data_bits_T_2 & _GEN_1741) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_29_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_29_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_29_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1646) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_29_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_29_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_29_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_29_bits_committed <= ~_GEN_2472 & (commit_store_3 ? _GEN_2376 | _GEN_2312 | _GEN_137979 : _GEN_2312 | _GEN_137979);
    stq_29_bits_succeeded <= ~_GEN_2472 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1D | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1D | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h1D)) & _GEN_1457 & _GEN_1393 & _GEN_1361 & _GEN_1297 & stq_29_bits_succeeded);
    stq_30_valid <= ~_GEN_2509 & (clear_store ? ~_GEN_2441 & _GEN_52446 : ~_GEN_2027 & _GEN_52446);
    stq_30_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & mem_xcpt_uops_1_stq_idx == 5'h1E | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & mem_xcpt_uops_0_stq_idx == 5'h1E | (_GEN_1458 ? (_GEN_1394 ? (_GEN_1362 ? (_GEN_1298 ? stq_30_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_30_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1458 ? (_GEN_1394 ? (_GEN_1362 ? (_GEN_1298 ? stq_30_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_30_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1458 ? (_GEN_1394 ? (_GEN_1362 ? (_GEN_1298 ? stq_30_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_30_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1458 ? (_GEN_1394 ? (_GEN_1362 ? (_GEN_1298 ? stq_30_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_30_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1458 ? (_GEN_1394 ? (_GEN_1362 ? (_GEN_1298 ? stq_30_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_30_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1458 ? (_GEN_1394 ? (_GEN_1362 ? (_GEN_1298 ? stq_30_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_30_bits_addr_valid <= ~_GEN_2509 & (clear_store ? ~_GEN_2441 & _GEN_82036 : ~_GEN_2027 & _GEN_82036);
    if (_GEN_1710) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_30_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_30_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_30_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_30_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_30_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_30_bits_addr_bits <= hella_req_addr;
        else
          stq_30_bits_addr_bits <= 40'h0;
      end
      else
        stq_30_bits_addr_bits <= _GEN_338;
      stq_30_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1615) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_30_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_30_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_30_bits_addr_bits <= _GEN_332;
        else
          stq_30_bits_addr_bits <= 40'h0;
      end
      else
        stq_30_bits_addr_bits <= _GEN_334;
      stq_30_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_30_bits_data_valid <= ~_GEN_2509 & (clear_store ? ~_GEN_2441 & _GEN_82260 : ~_GEN_2027 & _GEN_82260);
    if (_stq_bits_data_bits_T_2 & _GEN_1742) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_30_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_30_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_30_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1647) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_30_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_30_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_30_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_30_bits_committed <= ~_GEN_2473 & (commit_store_3 ? _GEN_2377 | _GEN_2313 | _GEN_137980 : _GEN_2313 | _GEN_137980);
    stq_30_bits_succeeded <= ~_GEN_2473 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & io_dmem_resp_1_bits_uop_stq_idx == 5'h1E | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & io_dmem_resp_0_bits_uop_stq_idx == 5'h1E | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & stq_execute_head == 5'h1E)) & _GEN_1458 & _GEN_1394 & _GEN_1362 & _GEN_1298 & stq_30_bits_succeeded);
    stq_31_valid <= ~_GEN_2510 & (clear_store ? ~_GEN_2442 & _GEN_52447 : ~_GEN_2028 & _GEN_52447);
    stq_31_bits_uop_exception <= ~_GEN_1235 & (mem_xcpt_valids_1 & ~mem_xcpt_uops_1_uses_ldq & (&mem_xcpt_uops_1_stq_idx) | mem_xcpt_valids_0 & ~mem_xcpt_uops_0_uses_ldq & (&mem_xcpt_uops_0_stq_idx) | (_GEN_1459 ? (_GEN_1395 ? (_GEN_1363 ? (_GEN_1299 ? stq_31_bits_uop_exception : io_core_dis_uops_0_bits_exception) : io_core_dis_uops_1_bits_exception) : io_core_dis_uops_2_bits_exception) : io_core_dis_uops_3_bits_exception));
    stq_31_bits_uop_mem_signed <= ~_GEN_1235 & (_GEN_1459 ? (_GEN_1395 ? (_GEN_1363 ? (_GEN_1299 ? stq_31_bits_uop_mem_signed : io_core_dis_uops_0_bits_mem_signed) : io_core_dis_uops_1_bits_mem_signed) : io_core_dis_uops_2_bits_mem_signed) : io_core_dis_uops_3_bits_mem_signed);
    stq_31_bits_uop_is_fence <= ~_GEN_1235 & (_GEN_1459 ? (_GEN_1395 ? (_GEN_1363 ? (_GEN_1299 ? stq_31_bits_uop_is_fence : io_core_dis_uops_0_bits_is_fence) : io_core_dis_uops_1_bits_is_fence) : io_core_dis_uops_2_bits_is_fence) : io_core_dis_uops_3_bits_is_fence);
    stq_31_bits_uop_is_amo <= ~_GEN_1235 & (_GEN_1459 ? (_GEN_1395 ? (_GEN_1363 ? (_GEN_1299 ? stq_31_bits_uop_is_amo : io_core_dis_uops_0_bits_is_amo) : io_core_dis_uops_1_bits_is_amo) : io_core_dis_uops_2_bits_is_amo) : io_core_dis_uops_3_bits_is_amo);
    stq_31_bits_uop_uses_ldq <= ~_GEN_1235 & (_GEN_1459 ? (_GEN_1395 ? (_GEN_1363 ? (_GEN_1299 ? stq_31_bits_uop_uses_ldq : io_core_dis_uops_0_bits_uses_ldq) : io_core_dis_uops_1_bits_uses_ldq) : io_core_dis_uops_2_bits_uses_ldq) : io_core_dis_uops_3_bits_uses_ldq);
    stq_31_bits_uop_uses_stq <= ~_GEN_1235 & (_GEN_1459 ? (_GEN_1395 ? (_GEN_1363 ? (_GEN_1299 ? stq_31_bits_uop_uses_stq : io_core_dis_uops_0_bits_uses_stq) : io_core_dis_uops_1_bits_uses_stq) : io_core_dis_uops_2_bits_uses_stq) : io_core_dis_uops_3_bits_uses_stq);
    stq_31_bits_addr_valid <= ~_GEN_2510 & (clear_store ? ~_GEN_2442 & _GEN_82037 : ~_GEN_2028 & _GEN_82037);
    if (_GEN_1711) begin
      if (exe_tlb_miss_1) begin
        if (_exe_tlb_vaddr_T_8) begin
          if (_GEN_329)
            stq_31_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_31_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_1)
          stq_31_bits_addr_bits <= _GEN_333;
        else if (will_fire_load_retry_1)
          stq_31_bits_addr_bits <= casez_tmp_79;
        else if (will_fire_sta_retry_1)
          stq_31_bits_addr_bits <= casez_tmp_78;
        else if (will_fire_hella_incoming_1)
          stq_31_bits_addr_bits <= hella_req_addr;
        else
          stq_31_bits_addr_bits <= 40'h0;
      end
      else
        stq_31_bits_addr_bits <= _GEN_338;
      stq_31_bits_addr_is_virtual <= exe_tlb_miss_1;
    end
    else if (_GEN_1616) begin
      if (exe_tlb_miss_0) begin
        if (_exe_tlb_vaddr_T_1) begin
          if (io_core_exe_1_req_bits_sfence_valid)
            stq_31_bits_addr_bits <= io_core_exe_1_req_bits_addr;
          else
            stq_31_bits_addr_bits <= io_core_exe_0_req_bits_addr;
        end
        else if (will_fire_sfence_0)
          stq_31_bits_addr_bits <= _GEN_332;
        else
          stq_31_bits_addr_bits <= 40'h0;
      end
      else
        stq_31_bits_addr_bits <= _GEN_334;
      stq_31_bits_addr_is_virtual <= exe_tlb_miss_0;
    end
    stq_31_bits_data_valid <= ~_GEN_2510 & (clear_store ? ~_GEN_2442 & _GEN_82261 : ~_GEN_2028 & _GEN_82261);
    if (_stq_bits_data_bits_T_2 & (&sidx_1)) begin
      if (_stq_bits_data_bits_T_2) begin
        if (_GEN_329)
          stq_31_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_31_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_31_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    else if (_GEN_1648) begin
      if (_stq_bits_data_bits_T) begin
        if (io_core_exe_1_req_bits_sfence_valid)
          stq_31_bits_data_bits <= io_core_exe_1_req_bits_data;
        else
          stq_31_bits_data_bits <= io_core_exe_0_req_bits_data;
      end
      else
        stq_31_bits_data_bits <= io_core_fp_stdata_bits_data;
    end
    stq_31_bits_committed <= ~_GEN_2474 & (commit_store_3 ? (&idx_3) | _GEN_2314 | _GEN_137981 : _GEN_2314 | _GEN_137981);
    stq_31_bits_succeeded <= ~_GEN_2474 & (io_dmem_resp_1_valid & ~io_dmem_resp_1_bits_uop_uses_ldq & io_dmem_resp_1_bits_uop_uses_stq & (&io_dmem_resp_1_bits_uop_stq_idx) | io_dmem_resp_0_valid & ~io_dmem_resp_0_bits_uop_uses_ldq & io_dmem_resp_0_bits_uop_uses_stq & (&io_dmem_resp_0_bits_uop_stq_idx) | (can_fire_load_incoming_0 | ~(will_fire_store_commit_0 & (&stq_execute_head))) & _GEN_1459 & _GEN_1395 & _GEN_1363 & _GEN_1299 & stq_31_bits_succeeded);
    if (_GEN_1234) begin
      ldq_head <= 5'h0;
      ldq_tail <= 5'h0;
      if (reset)
        stq_tail <= 5'h0;
      else
        stq_tail <= stq_commit_head;
    end
    else begin
      if (commit_load_3)
        ldq_head <= _GEN_1229 + 5'h1;
      else if (commit_load_2)
        ldq_head <= _GEN_1228;
      else if (commit_load_1)
        ldq_head <= _GEN_1224;
      else if (commit_load)
        ldq_head <= _GEN_1220;
      if (io_core_brupdate_b2_mispredict & ~io_core_exception) begin
        ldq_tail <= io_core_brupdate_b2_uop_ldq_idx;
        stq_tail <= io_core_brupdate_b2_uop_stq_idx;
      end
      else begin
        if (dis_ld_val_3)
          ldq_tail <= _GEN_232;
        else if (dis_ld_val_2)
          ldq_tail <= _GEN_165;
        else if (dis_ld_val_1)
          ldq_tail <= _GEN_67;
        else if (dis_ld_val)
          ldq_tail <= _GEN_0;
        if (dis_st_val_3)
          stq_tail <= _GEN_233;
        else if (dis_st_val_2)
          stq_tail <= _GEN_166;
        else if (dis_st_val_1)
          stq_tail <= _GEN_68;
        else if (dis_st_val)
          stq_tail <= _GEN_1;
      end
    end
    if (_GEN_2476) begin
      hella_req_addr <= io_hellacache_req_bits_addr;
      hella_req_cmd <= 5'h0;
      hella_req_size <= 2'h3;
    end
    hella_req_signed <= ~_GEN_2476 & hella_req_signed;
    hella_req_phys <= _GEN_2476 | hella_req_phys;
    if (_GEN_2477)
      hella_data_data <= 64'h0;
    if (_GEN_340 | ~will_fire_hella_incoming_1) begin
    end
    else
      hella_paddr <= exe_tlb_paddr_1;
    if (_GEN_2477) begin
      hella_xcpt_ma_ld <= _dtlb_io_resp_1_ma_ld;
      hella_xcpt_ma_st <= _dtlb_io_resp_1_ma_st;
      hella_xcpt_pf_ld <= _dtlb_io_resp_1_pf_ld;
      hella_xcpt_pf_st <= _dtlb_io_resp_1_pf_st;
    end
    hella_xcpt_gf_ld <= _GEN_2478 & hella_xcpt_gf_ld;
    hella_xcpt_gf_st <= _GEN_2478 & hella_xcpt_gf_st;
    if (_GEN_2477) begin
      hella_xcpt_ae_ld <= _dtlb_io_resp_1_ae_ld;
      hella_xcpt_ae_st <= _dtlb_io_resp_1_ae_st;
    end
    if (will_fire_load_wakeup_1) begin
      p1_block_load_mask_0 <= _GEN_68532;
      p1_block_load_mask_1 <= _GEN_68533;
      p1_block_load_mask_2 <= _GEN_68534;
      p1_block_load_mask_3 <= _GEN_68535;
      p1_block_load_mask_4 <= _GEN_68536;
      p1_block_load_mask_5 <= _GEN_68537;
      p1_block_load_mask_6 <= _GEN_68538;
      p1_block_load_mask_7 <= _GEN_68539;
      p1_block_load_mask_8 <= _GEN_68540;
      p1_block_load_mask_9 <= _GEN_68541;
      p1_block_load_mask_10 <= _GEN_68542;
      p1_block_load_mask_11 <= _GEN_68543;
      p1_block_load_mask_12 <= _GEN_68544;
      p1_block_load_mask_13 <= _GEN_68545;
      p1_block_load_mask_14 <= _GEN_68546;
      p1_block_load_mask_15 <= _GEN_68547;
      p1_block_load_mask_16 <= _GEN_68548;
      p1_block_load_mask_17 <= _GEN_68549;
      p1_block_load_mask_18 <= _GEN_68550;
      p1_block_load_mask_19 <= _GEN_68551;
      p1_block_load_mask_20 <= _GEN_68552;
      p1_block_load_mask_21 <= _GEN_68553;
      p1_block_load_mask_22 <= _GEN_68554;
      p1_block_load_mask_23 <= _GEN_68555;
      p1_block_load_mask_24 <= _GEN_68556;
      p1_block_load_mask_25 <= _GEN_68557;
      p1_block_load_mask_26 <= _GEN_68558;
      p1_block_load_mask_27 <= _GEN_68559;
      p1_block_load_mask_28 <= _GEN_68560;
      p1_block_load_mask_29 <= _GEN_68561;
      p1_block_load_mask_30 <= _GEN_68562;
      p1_block_load_mask_31 <= _GEN_68563;
    end
    else if (can_fire_load_incoming_1) begin
      p1_block_load_mask_0 <= _GEN_68564;
      p1_block_load_mask_1 <= _GEN_68565;
      p1_block_load_mask_2 <= _GEN_68566;
      p1_block_load_mask_3 <= _GEN_68567;
      p1_block_load_mask_4 <= _GEN_68568;
      p1_block_load_mask_5 <= _GEN_68569;
      p1_block_load_mask_6 <= _GEN_68570;
      p1_block_load_mask_7 <= _GEN_68571;
      p1_block_load_mask_8 <= _GEN_68572;
      p1_block_load_mask_9 <= _GEN_68573;
      p1_block_load_mask_10 <= _GEN_68574;
      p1_block_load_mask_11 <= _GEN_68575;
      p1_block_load_mask_12 <= _GEN_68576;
      p1_block_load_mask_13 <= _GEN_68577;
      p1_block_load_mask_14 <= _GEN_68578;
      p1_block_load_mask_15 <= _GEN_68579;
      p1_block_load_mask_16 <= _GEN_68580;
      p1_block_load_mask_17 <= _GEN_68581;
      p1_block_load_mask_18 <= _GEN_68582;
      p1_block_load_mask_19 <= _GEN_68583;
      p1_block_load_mask_20 <= _GEN_68584;
      p1_block_load_mask_21 <= _GEN_68585;
      p1_block_load_mask_22 <= _GEN_68586;
      p1_block_load_mask_23 <= _GEN_68587;
      p1_block_load_mask_24 <= _GEN_68588;
      p1_block_load_mask_25 <= _GEN_68589;
      p1_block_load_mask_26 <= _GEN_68590;
      p1_block_load_mask_27 <= _GEN_68591;
      p1_block_load_mask_28 <= _GEN_68592;
      p1_block_load_mask_29 <= _GEN_68593;
      p1_block_load_mask_30 <= _GEN_68594;
      p1_block_load_mask_31 <= _GEN_68595;
    end
    else begin
      p1_block_load_mask_0 <= _GEN_68628;
      p1_block_load_mask_1 <= _GEN_68629;
      p1_block_load_mask_2 <= _GEN_68630;
      p1_block_load_mask_3 <= _GEN_68631;
      p1_block_load_mask_4 <= _GEN_68632;
      p1_block_load_mask_5 <= _GEN_68633;
      p1_block_load_mask_6 <= _GEN_68634;
      p1_block_load_mask_7 <= _GEN_68635;
      p1_block_load_mask_8 <= _GEN_68636;
      p1_block_load_mask_9 <= _GEN_68637;
      p1_block_load_mask_10 <= _GEN_68638;
      p1_block_load_mask_11 <= _GEN_68639;
      p1_block_load_mask_12 <= _GEN_68640;
      p1_block_load_mask_13 <= _GEN_68641;
      p1_block_load_mask_14 <= _GEN_68642;
      p1_block_load_mask_15 <= _GEN_68643;
      p1_block_load_mask_16 <= _GEN_68644;
      p1_block_load_mask_17 <= _GEN_68645;
      p1_block_load_mask_18 <= _GEN_68646;
      p1_block_load_mask_19 <= _GEN_68647;
      p1_block_load_mask_20 <= _GEN_68648;
      p1_block_load_mask_21 <= _GEN_68649;
      p1_block_load_mask_22 <= _GEN_68650;
      p1_block_load_mask_23 <= _GEN_68651;
      p1_block_load_mask_24 <= _GEN_68652;
      p1_block_load_mask_25 <= _GEN_68653;
      p1_block_load_mask_26 <= _GEN_68654;
      p1_block_load_mask_27 <= _GEN_68655;
      p1_block_load_mask_28 <= _GEN_68656;
      p1_block_load_mask_29 <= _GEN_68657;
      p1_block_load_mask_30 <= _GEN_68658;
      p1_block_load_mask_31 <= _GEN_68659;
    end
    p2_block_load_mask_0 <= p1_block_load_mask_0;
    p2_block_load_mask_1 <= p1_block_load_mask_1;
    p2_block_load_mask_2 <= p1_block_load_mask_2;
    p2_block_load_mask_3 <= p1_block_load_mask_3;
    p2_block_load_mask_4 <= p1_block_load_mask_4;
    p2_block_load_mask_5 <= p1_block_load_mask_5;
    p2_block_load_mask_6 <= p1_block_load_mask_6;
    p2_block_load_mask_7 <= p1_block_load_mask_7;
    p2_block_load_mask_8 <= p1_block_load_mask_8;
    p2_block_load_mask_9 <= p1_block_load_mask_9;
    p2_block_load_mask_10 <= p1_block_load_mask_10;
    p2_block_load_mask_11 <= p1_block_load_mask_11;
    p2_block_load_mask_12 <= p1_block_load_mask_12;
    p2_block_load_mask_13 <= p1_block_load_mask_13;
    p2_block_load_mask_14 <= p1_block_load_mask_14;
    p2_block_load_mask_15 <= p1_block_load_mask_15;
    p2_block_load_mask_16 <= p1_block_load_mask_16;
    p2_block_load_mask_17 <= p1_block_load_mask_17;
    p2_block_load_mask_18 <= p1_block_load_mask_18;
    p2_block_load_mask_19 <= p1_block_load_mask_19;
    p2_block_load_mask_20 <= p1_block_load_mask_20;
    p2_block_load_mask_21 <= p1_block_load_mask_21;
    p2_block_load_mask_22 <= p1_block_load_mask_22;
    p2_block_load_mask_23 <= p1_block_load_mask_23;
    p2_block_load_mask_24 <= p1_block_load_mask_24;
    p2_block_load_mask_25 <= p1_block_load_mask_25;
    p2_block_load_mask_26 <= p1_block_load_mask_26;
    p2_block_load_mask_27 <= p1_block_load_mask_27;
    p2_block_load_mask_28 <= p1_block_load_mask_28;
    p2_block_load_mask_29 <= p1_block_load_mask_29;
    p2_block_load_mask_30 <= p1_block_load_mask_30;
    p2_block_load_mask_31 <= p1_block_load_mask_31;
    ldq_wakeup_idx <= _ldq_wakeup_idx_T_7 & _temp_bits_T ? 5'h0 : _ldq_wakeup_idx_T_15 & _temp_bits_T_2 ? 5'h1 : _ldq_wakeup_idx_T_23 & _temp_bits_T_4 ? 5'h2 : _ldq_wakeup_idx_T_31 & _temp_bits_T_6 ? 5'h3 : _ldq_wakeup_idx_T_39 & _temp_bits_T_8 ? 5'h4 : _ldq_wakeup_idx_T_47 & _temp_bits_T_10 ? 5'h5 : _ldq_wakeup_idx_T_55 & _temp_bits_T_12 ? 5'h6 : _ldq_wakeup_idx_T_63 & _temp_bits_T_14 ? 5'h7 : _ldq_wakeup_idx_T_71 & _temp_bits_T_16 ? 5'h8 : _ldq_wakeup_idx_T_79 & _temp_bits_T_18 ? 5'h9 : _ldq_wakeup_idx_T_87 & _temp_bits_T_20 ? 5'hA : _ldq_wakeup_idx_T_95 & _temp_bits_T_22 ? 5'hB : _ldq_wakeup_idx_T_103 & _temp_bits_T_24 ? 5'hC : _ldq_wakeup_idx_T_111 & _temp_bits_T_26 ? 5'hD : _ldq_wakeup_idx_T_119 & _temp_bits_T_28 ? 5'hE : _ldq_wakeup_idx_T_127 & ~(ldq_head[4]) ? 5'hF : _ldq_wakeup_idx_T_135 & _temp_bits_T_32 ? 5'h10 : _ldq_wakeup_idx_T_143 & _temp_bits_T_34 ? 5'h11 : _ldq_wakeup_idx_T_151 & _temp_bits_T_36 ? 5'h12 : _ldq_wakeup_idx_T_159 & _temp_bits_T_38 ? 5'h13 : _ldq_wakeup_idx_idx_T_42[4:0];
    ldq_retry_idx <= _ldq_retry_idx_T_2 & _temp_bits_T ? 5'h0 : _ldq_retry_idx_T_5 & _temp_bits_T_2 ? 5'h1 : _ldq_retry_idx_T_8 & _temp_bits_T_4 ? 5'h2 : _ldq_retry_idx_T_11 & _temp_bits_T_6 ? 5'h3 : _ldq_retry_idx_T_14 & _temp_bits_T_8 ? 5'h4 : _ldq_retry_idx_T_17 & _temp_bits_T_10 ? 5'h5 : _ldq_retry_idx_T_20 & _temp_bits_T_12 ? 5'h6 : _ldq_retry_idx_T_23 & _temp_bits_T_14 ? 5'h7 : _ldq_retry_idx_T_26 & _temp_bits_T_16 ? 5'h8 : _ldq_retry_idx_T_29 & _temp_bits_T_18 ? 5'h9 : _ldq_retry_idx_T_32 & _temp_bits_T_20 ? 5'hA : _ldq_retry_idx_T_35 & _temp_bits_T_22 ? 5'hB : _ldq_retry_idx_T_38 & _temp_bits_T_24 ? 5'hC : _ldq_retry_idx_T_41 & _temp_bits_T_26 ? 5'hD : _ldq_retry_idx_T_44 & _temp_bits_T_28 ? 5'hE : _ldq_retry_idx_T_47 & ~(ldq_head[4]) ? 5'hF : _ldq_retry_idx_T_50 & _temp_bits_T_32 ? 5'h10 : _ldq_retry_idx_T_53 & _temp_bits_T_34 ? 5'h11 : _ldq_retry_idx_T_56 & _temp_bits_T_36 ? 5'h12 : _ldq_retry_idx_T_59 & _temp_bits_T_38 ? 5'h13 : _ldq_retry_idx_idx_T_42[4:0];
    can_fire_load_retry_REG_1 <= _dtlb_io_miss_rdy;
    stq_retry_idx <= _stq_retry_idx_T & stq_commit_head == 5'h0 ? 5'h0 : _stq_retry_idx_T_1 & stq_commit_head < 5'h2 ? 5'h1 : _stq_retry_idx_T_2 & stq_commit_head < 5'h3 ? 5'h2 : _stq_retry_idx_T_3 & stq_commit_head < 5'h4 ? 5'h3 : _stq_retry_idx_T_4 & stq_commit_head < 5'h5 ? 5'h4 : _stq_retry_idx_T_5 & stq_commit_head < 5'h6 ? 5'h5 : _stq_retry_idx_T_6 & stq_commit_head < 5'h7 ? 5'h6 : _stq_retry_idx_T_7 & stq_commit_head < 5'h8 ? 5'h7 : _stq_retry_idx_T_8 & stq_commit_head < 5'h9 ? 5'h8 : _stq_retry_idx_T_9 & stq_commit_head < 5'hA ? 5'h9 : _stq_retry_idx_T_10 & stq_commit_head < 5'hB ? 5'hA : _stq_retry_idx_T_11 & stq_commit_head < 5'hC ? 5'hB : _stq_retry_idx_T_12 & stq_commit_head < 5'hD ? 5'hC : _stq_retry_idx_T_13 & stq_commit_head < 5'hE ? 5'hD : _stq_retry_idx_T_14 & stq_commit_head < 5'hF ? 5'hE : _stq_retry_idx_T_15 & ~(stq_commit_head[4]) ? 5'hF : _stq_retry_idx_T_16 & stq_commit_head < 5'h11 ? 5'h10 : _stq_retry_idx_T_17 & stq_commit_head < 5'h12 ? 5'h11 : _stq_retry_idx_T_18 & stq_commit_head < 5'h13 ? 5'h12 : _stq_retry_idx_T_19 & stq_commit_head < 5'h14 ? 5'h13 : _stq_retry_idx_idx_T_42[4:0];
    can_fire_sta_retry_REG_1 <= _dtlb_io_miss_rdy;
    mem_xcpt_valids_0 <= (pf_ld_0 | pf_st_0 | ae_ld_0 | ~_will_fire_store_commit_0_T_2 & _dtlb_io_resp_0_ae_st & exe_tlb_uop_0_uses_stq | ma_ld_0 | ma_st_0) & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & exe_tlb_uop_0_br_mask) == 20'h0;
    mem_xcpt_valids_1 <= (pf_ld_1 | pf_st_1 | ae_ld_1 | ~_will_fire_store_commit_1_T_2 & _dtlb_io_resp_1_ae_st & exe_tlb_uop_1_uses_stq | ma_ld_1 | ma_st_1) & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & exe_tlb_uop_1_br_mask) == 20'h0;
    mem_xcpt_uops_0_br_mask <= exe_tlb_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask;
    if (_exe_tlb_uop_T_2) begin
      if (io_core_exe_1_req_bits_sfence_valid) begin
        mem_xcpt_uops_0_rob_idx <= io_core_exe_1_req_bits_uop_rob_idx;
        mem_xcpt_uops_0_stq_idx <= io_core_exe_1_req_bits_uop_stq_idx;
      end
      else begin
        mem_xcpt_uops_0_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;
        mem_xcpt_uops_0_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;
      end
    end
    else begin
      mem_xcpt_uops_0_rob_idx <= 7'h0;
      mem_xcpt_uops_0_stq_idx <= 5'h0;
    end
    mem_xcpt_uops_0_uses_ldq <= exe_tlb_uop_0_uses_ldq;
    mem_xcpt_uops_1_br_mask <= exe_tlb_uop_1_br_mask & ~io_core_brupdate_b1_resolve_mask;
    if (_exe_tlb_uop_T_9) begin
      if (_GEN_329) begin
        mem_xcpt_uops_1_rob_idx <= io_core_exe_1_req_bits_uop_rob_idx;
        mem_xcpt_uops_1_stq_idx <= io_core_exe_1_req_bits_uop_stq_idx;
        mem_xcpt_uops_1_uses_ldq <= io_core_exe_1_req_bits_uop_uses_ldq;
      end
      else begin
        mem_xcpt_uops_1_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;
        mem_xcpt_uops_1_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;
        mem_xcpt_uops_1_uses_ldq <= io_core_exe_0_req_bits_uop_uses_ldq;
      end
    end
    else if (will_fire_load_retry_1) begin
      mem_xcpt_uops_1_rob_idx <= casez_tmp_68;
      mem_xcpt_uops_1_stq_idx <= casez_tmp_70;
      mem_xcpt_uops_1_uses_ldq <= casez_tmp_76;
    end
    else begin
      if (will_fire_sta_retry_1) begin
        mem_xcpt_uops_1_rob_idx <= casez_tmp_57;
        mem_xcpt_uops_1_stq_idx <= casez_tmp_59;
      end
      else begin
        mem_xcpt_uops_1_rob_idx <= 7'h0;
        mem_xcpt_uops_1_stq_idx <= 5'h0;
      end
      mem_xcpt_uops_1_uses_ldq <= _exe_tlb_uop_T_11_uses_ldq;
    end
    if (ma_ld_0)
      mem_xcpt_causes_0 <= 4'h4;
    else if (ma_st_0)
      mem_xcpt_causes_0 <= 4'h6;
    else if (pf_ld_0)
      mem_xcpt_causes_0 <= 4'hD;
    else if (pf_st_0)
      mem_xcpt_causes_0 <= 4'hF;
    else
      mem_xcpt_causes_0 <= {2'h1, ~ae_ld_0, 1'h1};
    if (ma_ld_1)
      mem_xcpt_causes_1 <= 4'h4;
    else if (ma_st_1)
      mem_xcpt_causes_1 <= 4'h6;
    else if (pf_ld_1)
      mem_xcpt_causes_1 <= 4'hD;
    else if (pf_st_1)
      mem_xcpt_causes_1 <= 4'hF;
    else
      mem_xcpt_causes_1 <= {2'h1, ~ae_ld_1, 1'h1};
    if (_exe_tlb_vaddr_T_1) begin
      if (io_core_exe_1_req_bits_sfence_valid)
        mem_xcpt_vaddrs_0 <= io_core_exe_1_req_bits_addr;
      else
        mem_xcpt_vaddrs_0 <= io_core_exe_0_req_bits_addr;
    end
    else if (will_fire_sfence_0)
      mem_xcpt_vaddrs_0 <= _GEN_332;
    else
      mem_xcpt_vaddrs_0 <= 40'h0;
    if (_exe_tlb_vaddr_T_8) begin
      if (_GEN_329)
        mem_xcpt_vaddrs_1 <= io_core_exe_1_req_bits_addr;
      else
        mem_xcpt_vaddrs_1 <= io_core_exe_0_req_bits_addr;
    end
    else if (will_fire_sfence_1)
      mem_xcpt_vaddrs_1 <= _GEN_333;
    else if (will_fire_load_retry_1)
      mem_xcpt_vaddrs_1 <= casez_tmp_79;
    else if (will_fire_sta_retry_1)
      mem_xcpt_vaddrs_1 <= casez_tmp_78;
    else if (will_fire_hella_incoming_1)
      mem_xcpt_vaddrs_1 <= hella_req_addr;
    else
      mem_xcpt_vaddrs_1 <= 40'h0;
    fired_load_incoming_0 <= can_fire_load_incoming_0 & _fired_std_incoming_T;
    fired_load_incoming_1 <= can_fire_load_incoming_1 & _fired_std_incoming_T_2;
    fired_stad_incoming_0 <= will_fire_stad_incoming_0 & _fired_std_incoming_T;
    fired_stad_incoming_1 <= will_fire_stad_incoming_1 & _fired_std_incoming_T_2;
    fired_sta_incoming_0 <= will_fire_sta_incoming_0 & _fired_std_incoming_T;
    fired_sta_incoming_1 <= will_fire_sta_incoming_1 & _fired_std_incoming_T_2;
    fired_std_incoming_0 <= will_fire_std_incoming_0 & _fired_std_incoming_T;
    fired_std_incoming_1 <= will_fire_std_incoming_1 & _fired_std_incoming_T_2;
    fired_stdf_incoming <= fp_stdata_fire & (io_core_brupdate_b1_mispredict_mask & io_core_fp_stdata_bits_uop_br_mask) == 20'h0;
    fired_sfence_0 <= will_fire_sfence_0;
    fired_sfence_1 <= will_fire_sfence_1;
    fired_release_1 <= will_fire_release_1;
    fired_load_retry_1 <= will_fire_load_retry_1 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_67) == 20'h0;
    fired_sta_retry_1 <= will_fire_sta_retry_1 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_56) == 20'h0;
    fired_load_wakeup_1 <= will_fire_load_wakeup_1 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_92) == 20'h0;
    mem_incoming_uop_0_br_mask <= exe_req_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    if (io_core_exe_1_req_bits_sfence_valid) begin
      mem_incoming_uop_0_rob_idx <= io_core_exe_1_req_bits_uop_rob_idx;
      mem_incoming_uop_0_ldq_idx <= io_core_exe_1_req_bits_uop_ldq_idx;
      mem_incoming_uop_0_stq_idx <= io_core_exe_1_req_bits_uop_stq_idx;
      mem_incoming_uop_0_pdst <= io_core_exe_1_req_bits_uop_pdst;
      mem_incoming_uop_0_fp_val <= io_core_exe_1_req_bits_uop_fp_val;
    end
    else begin
      mem_incoming_uop_0_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;
      mem_incoming_uop_0_ldq_idx <= io_core_exe_0_req_bits_uop_ldq_idx;
      mem_incoming_uop_0_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;
      mem_incoming_uop_0_pdst <= io_core_exe_0_req_bits_uop_pdst;
      mem_incoming_uop_0_fp_val <= io_core_exe_0_req_bits_uop_fp_val;
    end
    mem_incoming_uop_1_br_mask <= exe_req_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    if (_GEN_329) begin
      mem_incoming_uop_1_rob_idx <= io_core_exe_1_req_bits_uop_rob_idx;
      mem_incoming_uop_1_ldq_idx <= io_core_exe_1_req_bits_uop_ldq_idx;
      mem_incoming_uop_1_stq_idx <= io_core_exe_1_req_bits_uop_stq_idx;
      mem_incoming_uop_1_pdst <= io_core_exe_1_req_bits_uop_pdst;
      mem_incoming_uop_1_fp_val <= io_core_exe_1_req_bits_uop_fp_val;
    end
    else begin
      mem_incoming_uop_1_rob_idx <= io_core_exe_0_req_bits_uop_rob_idx;
      mem_incoming_uop_1_ldq_idx <= io_core_exe_0_req_bits_uop_ldq_idx;
      mem_incoming_uop_1_stq_idx <= io_core_exe_0_req_bits_uop_stq_idx;
      mem_incoming_uop_1_pdst <= io_core_exe_0_req_bits_uop_pdst;
      mem_incoming_uop_1_fp_val <= io_core_exe_0_req_bits_uop_fp_val;
    end
    mem_ldq_incoming_e_0_bits_uop_br_mask <= casez_tmp_4 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_incoming_e_0_bits_uop_stq_idx <= casez_tmp_5;
    mem_ldq_incoming_e_0_bits_uop_mem_size <= casez_tmp_6;
    mem_ldq_incoming_e_0_bits_st_dep_mask <= casez_tmp_7;
    mem_ldq_incoming_e_1_bits_uop_br_mask <= casez_tmp_8 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_incoming_e_1_bits_uop_stq_idx <= casez_tmp_9;
    mem_ldq_incoming_e_1_bits_uop_mem_size <= casez_tmp_10;
    mem_ldq_incoming_e_1_bits_st_dep_mask <= casez_tmp_11;
    mem_stq_incoming_e_0_valid <= casez_tmp_12 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_13) == 20'h0;
    mem_stq_incoming_e_0_bits_uop_br_mask <= casez_tmp_13 & ~io_core_brupdate_b1_resolve_mask;
    mem_stq_incoming_e_0_bits_uop_rob_idx <= casez_tmp_14;
    mem_stq_incoming_e_0_bits_uop_stq_idx <= casez_tmp_15;
    mem_stq_incoming_e_0_bits_uop_mem_size <= casez_tmp_16;
    mem_stq_incoming_e_0_bits_uop_is_amo <= casez_tmp_17;
    mem_stq_incoming_e_0_bits_addr_valid <= casez_tmp_18;
    mem_stq_incoming_e_0_bits_addr_is_virtual <= casez_tmp_19;
    mem_stq_incoming_e_0_bits_data_valid <= casez_tmp_20;
    mem_stq_incoming_e_1_valid <= casez_tmp_21 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_22) == 20'h0;
    mem_stq_incoming_e_1_bits_uop_br_mask <= casez_tmp_22 & ~io_core_brupdate_b1_resolve_mask;
    mem_stq_incoming_e_1_bits_uop_rob_idx <= casez_tmp_23;
    mem_stq_incoming_e_1_bits_uop_stq_idx <= casez_tmp_24;
    mem_stq_incoming_e_1_bits_uop_mem_size <= casez_tmp_25;
    mem_stq_incoming_e_1_bits_uop_is_amo <= casez_tmp_26;
    mem_stq_incoming_e_1_bits_addr_valid <= casez_tmp_27;
    mem_stq_incoming_e_1_bits_addr_is_virtual <= casez_tmp_28;
    mem_stq_incoming_e_1_bits_data_valid <= casez_tmp_29;
    mem_ldq_wakeup_e_bits_uop_br_mask <= casez_tmp_92 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_wakeup_e_bits_uop_stq_idx <= casez_tmp_94;
    mem_ldq_wakeup_e_bits_uop_mem_size <= casez_tmp_96;
    mem_ldq_wakeup_e_bits_st_dep_mask <= casez_tmp_39;
    mem_ldq_retry_e_bits_uop_br_mask <= casez_tmp_67 & ~io_core_brupdate_b1_resolve_mask;
    mem_ldq_retry_e_bits_uop_stq_idx <= casez_tmp_70;
    mem_ldq_retry_e_bits_uop_mem_size <= casez_tmp_73;
    mem_ldq_retry_e_bits_st_dep_mask <= casez_tmp_102;
    mem_stq_retry_e_valid <= casez_tmp_46 & (io_core_brupdate_b1_mispredict_mask & casez_tmp_56) == 20'h0;
    mem_stq_retry_e_bits_uop_br_mask <= casez_tmp_56 & ~io_core_brupdate_b1_resolve_mask;
    mem_stq_retry_e_bits_uop_rob_idx <= casez_tmp_57;
    mem_stq_retry_e_bits_uop_stq_idx <= casez_tmp_59;
    mem_stq_retry_e_bits_uop_mem_size <= casez_tmp_62;
    mem_stq_retry_e_bits_uop_is_amo <= casez_tmp_64;
    mem_stq_retry_e_bits_data_valid <= casez_tmp_103;
    mem_stdf_uop_br_mask <= io_core_fp_stdata_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    mem_stdf_uop_rob_idx <= io_core_fp_stdata_bits_uop_rob_idx;
    mem_stdf_uop_stq_idx <= io_core_fp_stdata_bits_uop_stq_idx;
    mem_tlb_miss_0 <= exe_tlb_miss_0;
    mem_tlb_miss_1 <= exe_tlb_miss_1;
    mem_tlb_uncacheable_0 <= ~_dtlb_io_resp_0_cacheable;
    mem_tlb_uncacheable_1 <= ~_dtlb_io_resp_1_cacheable;
    if (can_fire_load_incoming_0)
      mem_paddr_0 <= _GEN_334;
    else if (will_fire_store_commit_0)
      mem_paddr_0 <= casez_tmp_80;
    else
      mem_paddr_0 <= 40'h0;
    if (_GEN_339)
      mem_paddr_1 <= _GEN_338;
    else if (will_fire_load_wakeup_1)
      mem_paddr_1 <= casez_tmp_91;
    else
      mem_paddr_1 <= _GEN_337;
    if (fired_stad_incoming_0 | fired_sta_incoming_0 | fired_std_incoming_0)
      clr_bsy_rob_idx_0 <= mem_stq_incoming_e_0_bits_uop_rob_idx;
    else if (fired_sfence_0)
      clr_bsy_rob_idx_0 <= mem_incoming_uop_0_rob_idx;
    else
      clr_bsy_rob_idx_0 <= 7'h0;
    if (fired_stad_incoming_1 | fired_sta_incoming_1 | fired_std_incoming_1)
      clr_bsy_rob_idx_1 <= mem_stq_incoming_e_1_bits_uop_rob_idx;
    else if (fired_sfence_1)
      clr_bsy_rob_idx_1 <= mem_incoming_uop_1_rob_idx;
    else if (fired_sta_retry_1)
      clr_bsy_rob_idx_1 <= mem_stq_retry_e_bits_uop_rob_idx;
    else
      clr_bsy_rob_idx_1 <= 7'h0;
    if (fired_stad_incoming_0)
      clr_bsy_brmask_0 <= mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (fired_sta_incoming_0)
      clr_bsy_brmask_0 <= mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (fired_std_incoming_0)
      clr_bsy_brmask_0 <= mem_stq_incoming_e_0_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (fired_sfence_0)
      clr_bsy_brmask_0 <= mem_incoming_uop_0_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else
      clr_bsy_brmask_0 <= 20'h0;
    if (fired_stad_incoming_1)
      clr_bsy_brmask_1 <= mem_stq_incoming_e_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (fired_sta_incoming_1)
      clr_bsy_brmask_1 <= mem_stq_incoming_e_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (fired_std_incoming_1)
      clr_bsy_brmask_1 <= mem_stq_incoming_e_1_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (fired_sfence_1)
      clr_bsy_brmask_1 <= mem_incoming_uop_1_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else if (fired_sta_retry_1)
      clr_bsy_brmask_1 <= mem_stq_retry_e_bits_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    else
      clr_bsy_brmask_1 <= 20'h0;
    io_core_clr_bsy_0_valid_REG <= io_core_exception;
    io_core_clr_bsy_0_valid_REG_1 <= io_core_exception;
    io_core_clr_bsy_0_valid_REG_2 <= io_core_clr_bsy_0_valid_REG_1;
    io_core_clr_bsy_1_valid_REG <= io_core_exception;
    io_core_clr_bsy_1_valid_REG_1 <= io_core_exception;
    io_core_clr_bsy_1_valid_REG_2 <= io_core_clr_bsy_1_valid_REG_1;
    if (fired_stdf_incoming) begin
      stdf_clr_bsy_rob_idx <= mem_stdf_uop_rob_idx;
      stdf_clr_bsy_brmask <= mem_stdf_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    end
    else begin
      stdf_clr_bsy_rob_idx <= 7'h0;
      stdf_clr_bsy_brmask <= 20'h0;
    end
    io_core_clr_bsy_2_valid_REG <= io_core_exception;
    io_core_clr_bsy_2_valid_REG_1 <= io_core_exception;
    io_core_clr_bsy_2_valid_REG_2 <= io_core_clr_bsy_2_valid_REG_1;
    lcam_addr_REG <= exe_tlb_paddr_0;
    lcam_addr_REG_2 <= exe_tlb_paddr_1;
    lcam_addr_REG_3 <= io_dmem_release_bits_address;
    lcam_ldq_idx_REG_2 <= ldq_wakeup_idx;
    lcam_ldq_idx_REG_3 <= ldq_retry_idx;
    lcam_stq_idx_REG_1 <= stq_retry_idx;
    if (can_fire_load_incoming_1 ? _GEN_1551 : will_fire_load_retry_1 ? _GEN_1552 : will_fire_load_wakeup_1 & _GEN_1550)
      s1_executing_loads_0 <= dmem_req_fire_1;
    else
      s1_executing_loads_0 <= can_fire_load_incoming_0 & ~(|ldq_incoming_idx_0) & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1460 : will_fire_load_retry_1 ? _GEN_1520 : will_fire_load_wakeup_1 & _GEN_1490)
      s1_executing_loads_1 <= dmem_req_fire_1;
    else
      s1_executing_loads_1 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1461 : will_fire_load_retry_1 ? _GEN_1521 : will_fire_load_wakeup_1 & _GEN_1491)
      s1_executing_loads_2 <= dmem_req_fire_1;
    else
      s1_executing_loads_2 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h2 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1462 : will_fire_load_retry_1 ? _GEN_1522 : will_fire_load_wakeup_1 & _GEN_1492)
      s1_executing_loads_3 <= dmem_req_fire_1;
    else
      s1_executing_loads_3 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h3 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1463 : will_fire_load_retry_1 ? _GEN_1523 : will_fire_load_wakeup_1 & _GEN_1493)
      s1_executing_loads_4 <= dmem_req_fire_1;
    else
      s1_executing_loads_4 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h4 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1464 : will_fire_load_retry_1 ? _GEN_1524 : will_fire_load_wakeup_1 & _GEN_1494)
      s1_executing_loads_5 <= dmem_req_fire_1;
    else
      s1_executing_loads_5 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h5 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1465 : will_fire_load_retry_1 ? _GEN_1525 : will_fire_load_wakeup_1 & _GEN_1495)
      s1_executing_loads_6 <= dmem_req_fire_1;
    else
      s1_executing_loads_6 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h6 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1466 : will_fire_load_retry_1 ? _GEN_1526 : will_fire_load_wakeup_1 & _GEN_1496)
      s1_executing_loads_7 <= dmem_req_fire_1;
    else
      s1_executing_loads_7 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h7 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1467 : will_fire_load_retry_1 ? _GEN_1527 : will_fire_load_wakeup_1 & _GEN_1497)
      s1_executing_loads_8 <= dmem_req_fire_1;
    else
      s1_executing_loads_8 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h8 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1468 : will_fire_load_retry_1 ? _GEN_1528 : will_fire_load_wakeup_1 & _GEN_1498)
      s1_executing_loads_9 <= dmem_req_fire_1;
    else
      s1_executing_loads_9 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h9 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1469 : will_fire_load_retry_1 ? _GEN_1529 : will_fire_load_wakeup_1 & _GEN_1499)
      s1_executing_loads_10 <= dmem_req_fire_1;
    else
      s1_executing_loads_10 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hA & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1470 : will_fire_load_retry_1 ? _GEN_1530 : will_fire_load_wakeup_1 & _GEN_1500)
      s1_executing_loads_11 <= dmem_req_fire_1;
    else
      s1_executing_loads_11 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hB & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1471 : will_fire_load_retry_1 ? _GEN_1531 : will_fire_load_wakeup_1 & _GEN_1501)
      s1_executing_loads_12 <= dmem_req_fire_1;
    else
      s1_executing_loads_12 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hC & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1472 : will_fire_load_retry_1 ? _GEN_1532 : will_fire_load_wakeup_1 & _GEN_1502)
      s1_executing_loads_13 <= dmem_req_fire_1;
    else
      s1_executing_loads_13 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hD & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1473 : will_fire_load_retry_1 ? _GEN_1533 : will_fire_load_wakeup_1 & _GEN_1503)
      s1_executing_loads_14 <= dmem_req_fire_1;
    else
      s1_executing_loads_14 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hE & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1474 : will_fire_load_retry_1 ? _GEN_1534 : will_fire_load_wakeup_1 & _GEN_1504)
      s1_executing_loads_15 <= dmem_req_fire_1;
    else
      s1_executing_loads_15 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'hF & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1475 : will_fire_load_retry_1 ? _GEN_1535 : will_fire_load_wakeup_1 & _GEN_1505)
      s1_executing_loads_16 <= dmem_req_fire_1;
    else
      s1_executing_loads_16 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h10 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1476 : will_fire_load_retry_1 ? _GEN_1536 : will_fire_load_wakeup_1 & _GEN_1506)
      s1_executing_loads_17 <= dmem_req_fire_1;
    else
      s1_executing_loads_17 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h11 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1477 : will_fire_load_retry_1 ? _GEN_1537 : will_fire_load_wakeup_1 & _GEN_1507)
      s1_executing_loads_18 <= dmem_req_fire_1;
    else
      s1_executing_loads_18 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h12 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1478 : will_fire_load_retry_1 ? _GEN_1538 : will_fire_load_wakeup_1 & _GEN_1508)
      s1_executing_loads_19 <= dmem_req_fire_1;
    else
      s1_executing_loads_19 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h13 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1479 : will_fire_load_retry_1 ? _GEN_1539 : will_fire_load_wakeup_1 & _GEN_1509)
      s1_executing_loads_20 <= dmem_req_fire_1;
    else
      s1_executing_loads_20 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h14 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1480 : will_fire_load_retry_1 ? _GEN_1540 : will_fire_load_wakeup_1 & _GEN_1510)
      s1_executing_loads_21 <= dmem_req_fire_1;
    else
      s1_executing_loads_21 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h15 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1481 : will_fire_load_retry_1 ? _GEN_1541 : will_fire_load_wakeup_1 & _GEN_1511)
      s1_executing_loads_22 <= dmem_req_fire_1;
    else
      s1_executing_loads_22 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h16 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1482 : will_fire_load_retry_1 ? _GEN_1542 : will_fire_load_wakeup_1 & _GEN_1512)
      s1_executing_loads_23 <= dmem_req_fire_1;
    else
      s1_executing_loads_23 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h17 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1483 : will_fire_load_retry_1 ? _GEN_1543 : will_fire_load_wakeup_1 & _GEN_1513)
      s1_executing_loads_24 <= dmem_req_fire_1;
    else
      s1_executing_loads_24 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h18 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1484 : will_fire_load_retry_1 ? _GEN_1544 : will_fire_load_wakeup_1 & _GEN_1514)
      s1_executing_loads_25 <= dmem_req_fire_1;
    else
      s1_executing_loads_25 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h19 & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1485 : will_fire_load_retry_1 ? _GEN_1545 : will_fire_load_wakeup_1 & _GEN_1515)
      s1_executing_loads_26 <= dmem_req_fire_1;
    else
      s1_executing_loads_26 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1A & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1486 : will_fire_load_retry_1 ? _GEN_1546 : will_fire_load_wakeup_1 & _GEN_1516)
      s1_executing_loads_27 <= dmem_req_fire_1;
    else
      s1_executing_loads_27 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1B & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1487 : will_fire_load_retry_1 ? _GEN_1547 : will_fire_load_wakeup_1 & _GEN_1517)
      s1_executing_loads_28 <= dmem_req_fire_1;
    else
      s1_executing_loads_28 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1C & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1488 : will_fire_load_retry_1 ? _GEN_1548 : will_fire_load_wakeup_1 & _GEN_1518)
      s1_executing_loads_29 <= dmem_req_fire_1;
    else
      s1_executing_loads_29 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1D & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? _GEN_1489 : will_fire_load_retry_1 ? _GEN_1549 : will_fire_load_wakeup_1 & _GEN_1519)
      s1_executing_loads_30 <= dmem_req_fire_1;
    else
      s1_executing_loads_30 <= can_fire_load_incoming_0 & ldq_incoming_idx_0 == 5'h1E & dmem_req_fire_0;
    if (can_fire_load_incoming_1 ? (&ldq_incoming_idx_1) : will_fire_load_retry_1 ? (&ldq_retry_idx) : will_fire_load_wakeup_1 & (&ldq_wakeup_idx))
      s1_executing_loads_31 <= dmem_req_fire_1;
    else
      s1_executing_loads_31 <= can_fire_load_incoming_0 & (&ldq_incoming_idx_0) & dmem_req_fire_0;
    wb_forward_valid_0 <= casez_tmp_176 & (io_core_brupdate_b1_mispredict_mask & (do_st_search_0 ? (_lcam_stq_idx_T ? mem_stq_incoming_e_0_bits_uop_br_mask : 20'h0) : _GEN_346 ? mem_ldq_incoming_e_0_bits_uop_br_mask : 20'h0)) == 20'h0 & ~io_core_exception & ~REG_2;
    wb_forward_valid_1 <= casez_tmp_177 & (io_core_brupdate_b1_mispredict_mask & (do_st_search_1 ? (_lcam_stq_idx_T_3 ? mem_stq_incoming_e_1_bits_uop_br_mask : fired_sta_retry_1 ? mem_stq_retry_e_bits_uop_br_mask : 20'h0) : do_ld_search_1 ? (fired_load_incoming_1 ? mem_ldq_incoming_e_1_bits_uop_br_mask : fired_load_retry_1 ? mem_ldq_retry_e_bits_uop_br_mask : fired_load_wakeup_1 ? mem_ldq_wakeup_e_bits_uop_br_mask : 20'h0) : 20'h0)) == 20'h0 & ~io_core_exception & ~REG_3;
    if (fired_load_incoming_0)
      wb_forward_ldq_idx_0 <= mem_incoming_uop_0_ldq_idx;
    else
      wb_forward_ldq_idx_0 <= 5'h0;
    if (fired_load_incoming_1)
      wb_forward_ldq_idx_1 <= mem_incoming_uop_1_ldq_idx;
    else if (fired_load_wakeup_1)
      wb_forward_ldq_idx_1 <= lcam_ldq_idx_REG_2;
    else if (fired_load_retry_1)
      wb_forward_ldq_idx_1 <= lcam_ldq_idx_REG_3;
    else
      wb_forward_ldq_idx_1 <= 5'h0;
    if (_lcam_stq_idx_T)
      wb_forward_ld_addr_0 <= _GEN_343;
    else
      wb_forward_ld_addr_0 <= mem_paddr_0;
    if (_lcam_addr_T_5)
      wb_forward_ld_addr_1 <= _GEN_345;
    else if (fired_release_1)
      wb_forward_ld_addr_1 <= _GEN_344;
    else
      wb_forward_ld_addr_1 <= mem_paddr_1;
    wb_forward_stq_idx_0 <= _forwarding_age_logic_0_io_forwarding_idx;
    wb_forward_stq_idx_1 <= _forwarding_age_logic_1_io_forwarding_idx;
    older_nacked_REG <= nacking_loads_0;
    io_dmem_s1_kill_0_REG <= dmem_req_fire_0;
    older_nacked_REG_1 <= nacking_loads_0;
    io_dmem_s1_kill_1_REG <= dmem_req_fire_1;
    older_nacked_REG_2 <= nacking_loads_1;
    io_dmem_s1_kill_0_REG_1 <= dmem_req_fire_0;
    older_nacked_REG_3 <= nacking_loads_1;
    io_dmem_s1_kill_1_REG_1 <= dmem_req_fire_1;
    older_nacked_REG_4 <= nacking_loads_2;
    io_dmem_s1_kill_0_REG_2 <= dmem_req_fire_0;
    older_nacked_REG_5 <= nacking_loads_2;
    io_dmem_s1_kill_1_REG_2 <= dmem_req_fire_1;
    older_nacked_REG_6 <= nacking_loads_3;
    io_dmem_s1_kill_0_REG_3 <= dmem_req_fire_0;
    older_nacked_REG_7 <= nacking_loads_3;
    io_dmem_s1_kill_1_REG_3 <= dmem_req_fire_1;
    older_nacked_REG_8 <= nacking_loads_4;
    io_dmem_s1_kill_0_REG_4 <= dmem_req_fire_0;
    older_nacked_REG_9 <= nacking_loads_4;
    io_dmem_s1_kill_1_REG_4 <= dmem_req_fire_1;
    older_nacked_REG_10 <= nacking_loads_5;
    io_dmem_s1_kill_0_REG_5 <= dmem_req_fire_0;
    older_nacked_REG_11 <= nacking_loads_5;
    io_dmem_s1_kill_1_REG_5 <= dmem_req_fire_1;
    older_nacked_REG_12 <= nacking_loads_6;
    io_dmem_s1_kill_0_REG_6 <= dmem_req_fire_0;
    older_nacked_REG_13 <= nacking_loads_6;
    io_dmem_s1_kill_1_REG_6 <= dmem_req_fire_1;
    older_nacked_REG_14 <= nacking_loads_7;
    io_dmem_s1_kill_0_REG_7 <= dmem_req_fire_0;
    older_nacked_REG_15 <= nacking_loads_7;
    io_dmem_s1_kill_1_REG_7 <= dmem_req_fire_1;
    older_nacked_REG_16 <= nacking_loads_8;
    io_dmem_s1_kill_0_REG_8 <= dmem_req_fire_0;
    older_nacked_REG_17 <= nacking_loads_8;
    io_dmem_s1_kill_1_REG_8 <= dmem_req_fire_1;
    older_nacked_REG_18 <= nacking_loads_9;
    io_dmem_s1_kill_0_REG_9 <= dmem_req_fire_0;
    older_nacked_REG_19 <= nacking_loads_9;
    io_dmem_s1_kill_1_REG_9 <= dmem_req_fire_1;
    older_nacked_REG_20 <= nacking_loads_10;
    io_dmem_s1_kill_0_REG_10 <= dmem_req_fire_0;
    older_nacked_REG_21 <= nacking_loads_10;
    io_dmem_s1_kill_1_REG_10 <= dmem_req_fire_1;
    older_nacked_REG_22 <= nacking_loads_11;
    io_dmem_s1_kill_0_REG_11 <= dmem_req_fire_0;
    older_nacked_REG_23 <= nacking_loads_11;
    io_dmem_s1_kill_1_REG_11 <= dmem_req_fire_1;
    older_nacked_REG_24 <= nacking_loads_12;
    io_dmem_s1_kill_0_REG_12 <= dmem_req_fire_0;
    older_nacked_REG_25 <= nacking_loads_12;
    io_dmem_s1_kill_1_REG_12 <= dmem_req_fire_1;
    older_nacked_REG_26 <= nacking_loads_13;
    io_dmem_s1_kill_0_REG_13 <= dmem_req_fire_0;
    older_nacked_REG_27 <= nacking_loads_13;
    io_dmem_s1_kill_1_REG_13 <= dmem_req_fire_1;
    older_nacked_REG_28 <= nacking_loads_14;
    io_dmem_s1_kill_0_REG_14 <= dmem_req_fire_0;
    older_nacked_REG_29 <= nacking_loads_14;
    io_dmem_s1_kill_1_REG_14 <= dmem_req_fire_1;
    older_nacked_REG_30 <= nacking_loads_15;
    io_dmem_s1_kill_0_REG_15 <= dmem_req_fire_0;
    older_nacked_REG_31 <= nacking_loads_15;
    io_dmem_s1_kill_1_REG_15 <= dmem_req_fire_1;
    older_nacked_REG_32 <= nacking_loads_16;
    io_dmem_s1_kill_0_REG_16 <= dmem_req_fire_0;
    older_nacked_REG_33 <= nacking_loads_16;
    io_dmem_s1_kill_1_REG_16 <= dmem_req_fire_1;
    older_nacked_REG_34 <= nacking_loads_17;
    io_dmem_s1_kill_0_REG_17 <= dmem_req_fire_0;
    older_nacked_REG_35 <= nacking_loads_17;
    io_dmem_s1_kill_1_REG_17 <= dmem_req_fire_1;
    older_nacked_REG_36 <= nacking_loads_18;
    io_dmem_s1_kill_0_REG_18 <= dmem_req_fire_0;
    older_nacked_REG_37 <= nacking_loads_18;
    io_dmem_s1_kill_1_REG_18 <= dmem_req_fire_1;
    older_nacked_REG_38 <= nacking_loads_19;
    io_dmem_s1_kill_0_REG_19 <= dmem_req_fire_0;
    older_nacked_REG_39 <= nacking_loads_19;
    io_dmem_s1_kill_1_REG_19 <= dmem_req_fire_1;
    older_nacked_REG_40 <= nacking_loads_20;
    io_dmem_s1_kill_0_REG_20 <= dmem_req_fire_0;
    older_nacked_REG_41 <= nacking_loads_20;
    io_dmem_s1_kill_1_REG_20 <= dmem_req_fire_1;
    older_nacked_REG_42 <= nacking_loads_21;
    io_dmem_s1_kill_0_REG_21 <= dmem_req_fire_0;
    older_nacked_REG_43 <= nacking_loads_21;
    io_dmem_s1_kill_1_REG_21 <= dmem_req_fire_1;
    older_nacked_REG_44 <= nacking_loads_22;
    io_dmem_s1_kill_0_REG_22 <= dmem_req_fire_0;
    older_nacked_REG_45 <= nacking_loads_22;
    io_dmem_s1_kill_1_REG_22 <= dmem_req_fire_1;
    older_nacked_REG_46 <= nacking_loads_23;
    io_dmem_s1_kill_0_REG_23 <= dmem_req_fire_0;
    older_nacked_REG_47 <= nacking_loads_23;
    io_dmem_s1_kill_1_REG_23 <= dmem_req_fire_1;
    older_nacked_REG_48 <= nacking_loads_24;
    io_dmem_s1_kill_0_REG_24 <= dmem_req_fire_0;
    older_nacked_REG_49 <= nacking_loads_24;
    io_dmem_s1_kill_1_REG_24 <= dmem_req_fire_1;
    older_nacked_REG_50 <= nacking_loads_25;
    io_dmem_s1_kill_0_REG_25 <= dmem_req_fire_0;
    older_nacked_REG_51 <= nacking_loads_25;
    io_dmem_s1_kill_1_REG_25 <= dmem_req_fire_1;
    older_nacked_REG_52 <= nacking_loads_26;
    io_dmem_s1_kill_0_REG_26 <= dmem_req_fire_0;
    older_nacked_REG_53 <= nacking_loads_26;
    io_dmem_s1_kill_1_REG_26 <= dmem_req_fire_1;
    older_nacked_REG_54 <= nacking_loads_27;
    io_dmem_s1_kill_0_REG_27 <= dmem_req_fire_0;
    older_nacked_REG_55 <= nacking_loads_27;
    io_dmem_s1_kill_1_REG_27 <= dmem_req_fire_1;
    older_nacked_REG_56 <= nacking_loads_28;
    io_dmem_s1_kill_0_REG_28 <= dmem_req_fire_0;
    older_nacked_REG_57 <= nacking_loads_28;
    io_dmem_s1_kill_1_REG_28 <= dmem_req_fire_1;
    older_nacked_REG_58 <= nacking_loads_29;
    io_dmem_s1_kill_0_REG_29 <= dmem_req_fire_0;
    older_nacked_REG_59 <= nacking_loads_29;
    io_dmem_s1_kill_1_REG_29 <= dmem_req_fire_1;
    older_nacked_REG_60 <= nacking_loads_30;
    io_dmem_s1_kill_0_REG_30 <= dmem_req_fire_0;
    older_nacked_REG_61 <= nacking_loads_30;
    io_dmem_s1_kill_1_REG_30 <= dmem_req_fire_1;
    older_nacked_REG_62 <= nacking_loads_31;
    io_dmem_s1_kill_0_REG_31 <= dmem_req_fire_0;
    older_nacked_REG_63 <= nacking_loads_31;
    io_dmem_s1_kill_1_REG_31 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_32 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_33 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_34 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_32 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_33 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_34 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_35 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_36 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_37 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_35 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_36 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_37 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_38 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_39 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_40 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_38 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_39 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_40 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_41 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_42 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_43 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_41 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_42 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_43 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_44 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_45 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_46 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_44 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_45 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_46 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_47 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_48 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_49 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_47 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_48 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_49 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_50 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_51 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_52 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_50 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_51 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_52 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_53 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_54 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_55 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_53 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_54 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_55 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_56 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_57 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_58 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_56 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_57 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_58 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_59 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_60 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_61 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_59 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_60 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_61 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_62 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_63 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_64 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_62 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_63 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_64 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_65 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_66 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_67 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_65 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_66 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_67 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_68 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_69 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_70 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_68 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_69 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_70 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_71 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_72 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_73 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_71 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_72 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_73 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_74 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_75 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_76 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_74 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_75 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_76 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_77 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_78 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_79 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_77 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_78 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_79 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_80 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_81 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_82 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_80 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_81 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_82 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_83 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_84 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_85 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_83 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_84 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_85 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_86 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_87 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_88 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_86 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_87 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_88 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_89 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_90 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_91 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_89 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_90 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_91 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_92 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_93 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_94 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_92 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_93 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_94 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_95 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_96 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_97 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_95 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_96 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_97 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_98 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_99 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_100 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_98 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_99 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_100 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_101 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_102 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_103 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_101 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_102 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_103 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_104 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_105 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_106 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_104 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_105 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_106 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_107 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_108 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_109 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_107 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_108 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_109 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_110 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_111 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_112 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_110 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_111 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_112 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_113 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_114 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_115 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_113 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_114 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_115 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_116 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_117 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_118 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_116 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_117 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_118 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_119 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_120 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_121 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_119 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_120 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_121 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_122 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_123 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_124 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_122 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_123 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_124 <= dmem_req_fire_1;
    io_dmem_s1_kill_0_REG_125 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_126 <= dmem_req_fire_0;
    io_dmem_s1_kill_0_REG_127 <= dmem_req_fire_0;
    io_dmem_s1_kill_1_REG_125 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_126 <= dmem_req_fire_1;
    io_dmem_s1_kill_1_REG_127 <= dmem_req_fire_1;
    REG_2 <= io_core_exception;
    REG_3 <= io_core_exception;
    r_xcpt_uop_br_mask <= xcpt_uop_br_mask & ~io_core_brupdate_b1_resolve_mask;
    if (use_mem_xcpt) begin
      if (is_older)
        r_xcpt_uop_rob_idx <= mem_xcpt_uops_1_rob_idx;
      else
        r_xcpt_uop_rob_idx <= mem_xcpt_uops_0_rob_idx;
      r_xcpt_cause <= {1'h0, is_older ? mem_xcpt_causes_1 : mem_xcpt_causes_0};
    end
    else begin
      r_xcpt_uop_rob_idx <= casez_tmp_178;
      r_xcpt_cause <= 5'h10;
    end
    if (is_older)
      r_xcpt_badvaddr <= mem_xcpt_vaddrs_1;
    else
      r_xcpt_badvaddr <= mem_xcpt_vaddrs_0;
    io_core_ld_miss_REG <= _io_core_spec_ld_wakeup_0_valid_output | _io_core_spec_ld_wakeup_1_valid_output;
    spec_ld_succeed_REG <= _io_core_spec_ld_wakeup_0_valid_output;
    spec_ld_succeed_REG_1 <= mem_incoming_uop_0_ldq_idx;
    spec_ld_succeed_REG_2 <= _io_core_spec_ld_wakeup_1_valid_output;
    spec_ld_succeed_REG_3 <= mem_incoming_uop_1_ldq_idx;
    if (reset) begin
      hella_state <= 3'h0;
      live_store_mask <= 32'h0;
      clr_bsy_valid_0 <= 1'h0;
      clr_bsy_valid_1 <= 1'h0;
      stdf_clr_bsy_valid <= 1'h0;
      r_xcpt_valid <= 1'h0;
    end
    else begin
      if (|hella_state)
        hella_state <= casez_tmp_246;
      else if (_GEN_2475)
        hella_state <= 3'h1;
      live_store_mask <=
        ({32{dis_st_val_3}} & 32'h1 << _ldq_T_115_bits_youngest_stq_idx | _ldq_T_115_bits_st_dep_mask) & ~{stq_31_valid & (|_GEN_1217), stq_30_valid & (|_GEN_1216), stq_29_valid & (|_GEN_1215), stq_28_valid & (|_GEN_1214), stq_27_valid & (|_GEN_1213), stq_26_valid & (|_GEN_1212), stq_25_valid & (|_GEN_1211), stq_24_valid & (|_GEN_1210), stq_23_valid & (|_GEN_1209), stq_22_valid & (|_GEN_1208), stq_21_valid & (|_GEN_1207), stq_20_valid & (|_GEN_1206), stq_19_valid & (|_GEN_1205), stq_18_valid & (|_GEN_1204), stq_17_valid & (|_GEN_1203), stq_16_valid & (|_GEN_1202), stq_15_valid & (|_GEN_1201), stq_14_valid & (|_GEN_1200), stq_13_valid & (|_GEN_1199), stq_12_valid & (|_GEN_1198), stq_11_valid & (|_GEN_1197), stq_10_valid & (|_GEN_1196), stq_9_valid & (|_GEN_1195), stq_8_valid & (|_GEN_1194), stq_7_valid & (|_GEN_1193), stq_6_valid & (|_GEN_1192), stq_5_valid & (|_GEN_1191), stq_4_valid & (|_GEN_1190), stq_3_valid & (|_GEN_1189), stq_2_valid & (|_GEN_1188), stq_1_valid & (|_GEN_1187), stq_0_valid & (|_GEN_1186)}
        & ~{_GEN_1234 & ~reset & _GEN_140449, _GEN_1234 & ~reset & _GEN_140445, _GEN_1234 & ~reset & _GEN_140441, _GEN_1234 & ~reset & _GEN_140437, _GEN_1234 & ~reset & _GEN_140433, _GEN_1234 & ~reset & _GEN_140429, _GEN_1234 & ~reset & _GEN_140425, _GEN_1234 & ~reset & _GEN_140421, _GEN_1234 & ~reset & _GEN_140417, _GEN_1234 & ~reset & _GEN_140413, _GEN_1234 & ~reset & _GEN_140409, _GEN_1234 & ~reset & _GEN_140405, _GEN_1234 & ~reset & _GEN_140401, _GEN_1234 & ~reset & _GEN_140397, _GEN_1234 & ~reset & _GEN_140393, _GEN_1234 & ~reset & _GEN_140389, _GEN_1234 & ~reset & _GEN_140385, _GEN_1234 & ~reset & _GEN_140381, _GEN_1234 & ~reset & _GEN_140377, _GEN_1234 & ~reset & _GEN_140373, _GEN_1234 & ~reset & _GEN_140369, _GEN_1234 & ~reset & _GEN_140365, _GEN_1234 & ~reset & _GEN_140361, _GEN_1234 & ~reset & _GEN_140357, _GEN_1234 & ~reset & _GEN_140353, _GEN_1234 & ~reset & _GEN_140349, _GEN_1234 & ~reset & _GEN_140345, _GEN_1234 & ~reset & _GEN_140341, _GEN_1234 & ~reset & _GEN_140337, _GEN_1234 & ~reset & _GEN_140333, _GEN_1234 & ~reset & _GEN_140329, _GEN_1234 & ~reset & _GEN_140325};
      if (fired_stad_incoming_0)
        clr_bsy_valid_0 <= mem_stq_incoming_e_0_valid & ~mem_tlb_miss_0 & ~mem_stq_incoming_e_0_bits_uop_is_amo & _clr_bsy_valid_0_T_22 == 20'h0;
      else if (fired_sta_incoming_0)
        clr_bsy_valid_0 <= mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_data_valid & ~mem_tlb_miss_0 & ~mem_stq_incoming_e_0_bits_uop_is_amo & _clr_bsy_valid_0_T_22 == 20'h0;
      else if (fired_std_incoming_0)
        clr_bsy_valid_0 <= mem_stq_incoming_e_0_valid & mem_stq_incoming_e_0_bits_addr_valid & ~mem_stq_incoming_e_0_bits_addr_is_virtual & ~mem_stq_incoming_e_0_bits_uop_is_amo & _clr_bsy_valid_0_T_22 == 20'h0;
      else
        clr_bsy_valid_0 <= fired_sfence_0;
      if (fired_stad_incoming_1)
        clr_bsy_valid_1 <= mem_stq_incoming_e_1_valid & ~mem_tlb_miss_1 & ~mem_stq_incoming_e_1_bits_uop_is_amo & _clr_bsy_valid_1_T_22 == 20'h0;
      else if (fired_sta_incoming_1)
        clr_bsy_valid_1 <= mem_stq_incoming_e_1_valid & mem_stq_incoming_e_1_bits_data_valid & ~mem_tlb_miss_1 & ~mem_stq_incoming_e_1_bits_uop_is_amo & _clr_bsy_valid_1_T_22 == 20'h0;
      else if (fired_std_incoming_1)
        clr_bsy_valid_1 <= mem_stq_incoming_e_1_valid & mem_stq_incoming_e_1_bits_addr_valid & ~mem_stq_incoming_e_1_bits_addr_is_virtual & ~mem_stq_incoming_e_1_bits_uop_is_amo & _clr_bsy_valid_1_T_22 == 20'h0;
      else
        clr_bsy_valid_1 <= ~fired_sfence_1 & fired_sta_retry_1 & mem_stq_retry_e_valid & mem_stq_retry_e_bits_data_valid & ~mem_tlb_miss_1 & ~mem_stq_retry_e_bits_uop_is_amo & (io_core_brupdate_b1_mispredict_mask & mem_stq_retry_e_bits_uop_br_mask) == 20'h0;
      stdf_clr_bsy_valid <= fired_stdf_incoming & casez_tmp_104 & casez_tmp_105 & ~casez_tmp_106 & ~casez_tmp_107 & (io_core_brupdate_b1_mispredict_mask & mem_stdf_uop_br_mask) == 20'h0;
      r_xcpt_valid <= (ld_xcpt_valid | mem_xcpt_valid) & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & xcpt_uop_br_mask) == 20'h0;
    end
  end // always @(posedge)
  NBDTLB dtlb (
    .clock                        (clock),
    .reset                        (reset),
    .io_req_0_valid               (~_will_fire_store_commit_0_T_2),
    .io_req_0_bits_vaddr          (exe_tlb_vaddr_0),
    .io_req_0_bits_size           ((_exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0) & _exe_tlb_uop_T_2 ? mem_incoming_uop_out_mem_size : 2'h0),
    .io_req_0_bits_cmd            ((_exe_cmd_T | will_fire_sta_incoming_0 | will_fire_sfence_0) & _exe_tlb_uop_T_2 ? mem_incoming_uop_out_mem_cmd : 5'h0),
    .io_req_1_valid               (~_will_fire_store_commit_1_T_2),
    .io_req_1_bits_vaddr          (exe_tlb_vaddr_1),
    .io_req_1_bits_passthrough    (will_fire_hella_incoming_1 & hella_req_phys),
    .io_req_1_bits_size           (_exe_cmd_T_7 | will_fire_sta_incoming_1 | will_fire_sfence_1 | will_fire_load_retry_1 | will_fire_sta_retry_1 ? exe_tlb_uop_1_mem_size : will_fire_hella_incoming_1 ? hella_req_size : 2'h0),
    .io_req_1_bits_cmd            (_exe_cmd_T_7 | will_fire_sta_incoming_1 | will_fire_sfence_1 | will_fire_load_retry_1 | will_fire_sta_retry_1 ? exe_tlb_uop_1_mem_cmd : will_fire_hella_incoming_1 ? hella_req_cmd : 5'h0),
    .io_sfence_valid              (will_fire_sfence_1 ? exe_req_1_bits_sfence_valid : will_fire_sfence_0 & exe_req_0_bits_sfence_valid),
    .io_sfence_bits_rs1           (will_fire_sfence_1 ? (_GEN_329 ? io_core_exe_1_req_bits_sfence_bits_rs1 : io_core_exe_0_req_bits_sfence_bits_rs1) : will_fire_sfence_0 & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_bits_rs1 : io_core_exe_0_req_bits_sfence_bits_rs1)),
    .io_sfence_bits_rs2           (will_fire_sfence_1 ? (_GEN_329 ? io_core_exe_1_req_bits_sfence_bits_rs2 : io_core_exe_0_req_bits_sfence_bits_rs2) : will_fire_sfence_0 & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_sfence_bits_rs2 : io_core_exe_0_req_bits_sfence_bits_rs2)),
    .io_sfence_bits_addr          (will_fire_sfence_1 ? exe_req_1_bits_sfence_bits_addr : will_fire_sfence_0 ? exe_req_0_bits_sfence_bits_addr : 39'h0),
    .io_ptw_req_ready             (io_ptw_req_ready),
    .io_ptw_resp_valid            (io_ptw_resp_valid),
    .io_ptw_resp_bits_ae_final    (io_ptw_resp_bits_ae_final),
    .io_ptw_resp_bits_pte_ppn     (io_ptw_resp_bits_pte_ppn),
    .io_ptw_resp_bits_pte_d       (io_ptw_resp_bits_pte_d),
    .io_ptw_resp_bits_pte_a       (io_ptw_resp_bits_pte_a),
    .io_ptw_resp_bits_pte_g       (io_ptw_resp_bits_pte_g),
    .io_ptw_resp_bits_pte_u       (io_ptw_resp_bits_pte_u),
    .io_ptw_resp_bits_pte_x       (io_ptw_resp_bits_pte_x),
    .io_ptw_resp_bits_pte_w       (io_ptw_resp_bits_pte_w),
    .io_ptw_resp_bits_pte_r       (io_ptw_resp_bits_pte_r),
    .io_ptw_resp_bits_pte_v       (io_ptw_resp_bits_pte_v),
    .io_ptw_resp_bits_level       (io_ptw_resp_bits_level),
    .io_ptw_resp_bits_homogeneous (io_ptw_resp_bits_homogeneous),
    .io_ptw_ptbr_mode             (io_ptw_ptbr_mode),
    .io_ptw_status_dprv           (io_ptw_status_dprv),
    .io_ptw_status_mxr            (io_ptw_status_mxr),
    .io_ptw_status_sum            (io_ptw_status_sum),
    .io_ptw_pmp_0_cfg_l           (io_ptw_pmp_0_cfg_l),
    .io_ptw_pmp_0_cfg_a           (io_ptw_pmp_0_cfg_a),
    .io_ptw_pmp_0_cfg_x           (io_ptw_pmp_0_cfg_x),
    .io_ptw_pmp_0_cfg_w           (io_ptw_pmp_0_cfg_w),
    .io_ptw_pmp_0_cfg_r           (io_ptw_pmp_0_cfg_r),
    .io_ptw_pmp_0_addr            (io_ptw_pmp_0_addr),
    .io_ptw_pmp_0_mask            (io_ptw_pmp_0_mask),
    .io_ptw_pmp_1_cfg_l           (io_ptw_pmp_1_cfg_l),
    .io_ptw_pmp_1_cfg_a           (io_ptw_pmp_1_cfg_a),
    .io_ptw_pmp_1_cfg_x           (io_ptw_pmp_1_cfg_x),
    .io_ptw_pmp_1_cfg_w           (io_ptw_pmp_1_cfg_w),
    .io_ptw_pmp_1_cfg_r           (io_ptw_pmp_1_cfg_r),
    .io_ptw_pmp_1_addr            (io_ptw_pmp_1_addr),
    .io_ptw_pmp_1_mask            (io_ptw_pmp_1_mask),
    .io_ptw_pmp_2_cfg_l           (io_ptw_pmp_2_cfg_l),
    .io_ptw_pmp_2_cfg_a           (io_ptw_pmp_2_cfg_a),
    .io_ptw_pmp_2_cfg_x           (io_ptw_pmp_2_cfg_x),
    .io_ptw_pmp_2_cfg_w           (io_ptw_pmp_2_cfg_w),
    .io_ptw_pmp_2_cfg_r           (io_ptw_pmp_2_cfg_r),
    .io_ptw_pmp_2_addr            (io_ptw_pmp_2_addr),
    .io_ptw_pmp_2_mask            (io_ptw_pmp_2_mask),
    .io_ptw_pmp_3_cfg_l           (io_ptw_pmp_3_cfg_l),
    .io_ptw_pmp_3_cfg_a           (io_ptw_pmp_3_cfg_a),
    .io_ptw_pmp_3_cfg_x           (io_ptw_pmp_3_cfg_x),
    .io_ptw_pmp_3_cfg_w           (io_ptw_pmp_3_cfg_w),
    .io_ptw_pmp_3_cfg_r           (io_ptw_pmp_3_cfg_r),
    .io_ptw_pmp_3_addr            (io_ptw_pmp_3_addr),
    .io_ptw_pmp_3_mask            (io_ptw_pmp_3_mask),
    .io_ptw_pmp_4_cfg_l           (io_ptw_pmp_4_cfg_l),
    .io_ptw_pmp_4_cfg_a           (io_ptw_pmp_4_cfg_a),
    .io_ptw_pmp_4_cfg_x           (io_ptw_pmp_4_cfg_x),
    .io_ptw_pmp_4_cfg_w           (io_ptw_pmp_4_cfg_w),
    .io_ptw_pmp_4_cfg_r           (io_ptw_pmp_4_cfg_r),
    .io_ptw_pmp_4_addr            (io_ptw_pmp_4_addr),
    .io_ptw_pmp_4_mask            (io_ptw_pmp_4_mask),
    .io_ptw_pmp_5_cfg_l           (io_ptw_pmp_5_cfg_l),
    .io_ptw_pmp_5_cfg_a           (io_ptw_pmp_5_cfg_a),
    .io_ptw_pmp_5_cfg_x           (io_ptw_pmp_5_cfg_x),
    .io_ptw_pmp_5_cfg_w           (io_ptw_pmp_5_cfg_w),
    .io_ptw_pmp_5_cfg_r           (io_ptw_pmp_5_cfg_r),
    .io_ptw_pmp_5_addr            (io_ptw_pmp_5_addr),
    .io_ptw_pmp_5_mask            (io_ptw_pmp_5_mask),
    .io_ptw_pmp_6_cfg_l           (io_ptw_pmp_6_cfg_l),
    .io_ptw_pmp_6_cfg_a           (io_ptw_pmp_6_cfg_a),
    .io_ptw_pmp_6_cfg_x           (io_ptw_pmp_6_cfg_x),
    .io_ptw_pmp_6_cfg_w           (io_ptw_pmp_6_cfg_w),
    .io_ptw_pmp_6_cfg_r           (io_ptw_pmp_6_cfg_r),
    .io_ptw_pmp_6_addr            (io_ptw_pmp_6_addr),
    .io_ptw_pmp_6_mask            (io_ptw_pmp_6_mask),
    .io_ptw_pmp_7_cfg_l           (io_ptw_pmp_7_cfg_l),
    .io_ptw_pmp_7_cfg_a           (io_ptw_pmp_7_cfg_a),
    .io_ptw_pmp_7_cfg_x           (io_ptw_pmp_7_cfg_x),
    .io_ptw_pmp_7_cfg_w           (io_ptw_pmp_7_cfg_w),
    .io_ptw_pmp_7_cfg_r           (io_ptw_pmp_7_cfg_r),
    .io_ptw_pmp_7_addr            (io_ptw_pmp_7_addr),
    .io_ptw_pmp_7_mask            (io_ptw_pmp_7_mask),
    .io_kill                      (will_fire_hella_incoming_1 & io_hellacache_s1_kill),
    .io_miss_rdy                  (_dtlb_io_miss_rdy),
    .io_resp_0_miss               (_dtlb_io_resp_0_miss),
    .io_resp_0_paddr              (_dtlb_io_resp_0_paddr),
    .io_resp_0_pf_ld              (_dtlb_io_resp_0_pf_ld),
    .io_resp_0_pf_st              (_dtlb_io_resp_0_pf_st),
    .io_resp_0_ae_ld              (_dtlb_io_resp_0_ae_ld),
    .io_resp_0_ae_st              (_dtlb_io_resp_0_ae_st),
    .io_resp_0_cacheable          (_dtlb_io_resp_0_cacheable),
    .io_resp_1_miss               (_dtlb_io_resp_1_miss),
    .io_resp_1_paddr              (_dtlb_io_resp_1_paddr),
    .io_resp_1_pf_ld              (_dtlb_io_resp_1_pf_ld),
    .io_resp_1_pf_st              (_dtlb_io_resp_1_pf_st),
    .io_resp_1_ae_ld              (_dtlb_io_resp_1_ae_ld),
    .io_resp_1_ae_st              (_dtlb_io_resp_1_ae_st),
    .io_resp_1_ma_ld              (_dtlb_io_resp_1_ma_ld),
    .io_resp_1_ma_st              (_dtlb_io_resp_1_ma_st),
    .io_resp_1_cacheable          (_dtlb_io_resp_1_cacheable),
    .io_ptw_req_valid             (io_ptw_req_valid),
    .io_ptw_req_bits_valid        (io_ptw_req_bits_valid),
    .io_ptw_req_bits_bits_addr    (io_ptw_req_bits_bits_addr)
  );
  ForwardingAgeLogic forwarding_age_logic_0 (
    .io_addr_matches    ({_GEN_1171 & (_GEN_113704 | _GEN_1173 | _GEN_113869), _GEN_1165 & (_GEN_113236 | _GEN_1167 | _GEN_113401), _GEN_1159 & (_GEN_112768 | _GEN_1161 | _GEN_112933), _GEN_1153 & (_GEN_112300 | _GEN_1155 | _GEN_112465), _GEN_1147 & (_GEN_111832 | _GEN_1149 | _GEN_111997), _GEN_1141 & (_GEN_111364 | _GEN_1143 | _GEN_111529), _GEN_1135 & (_GEN_110896 | _GEN_1137 | _GEN_111061), _GEN_1129 & (_GEN_110428 | _GEN_1131 | _GEN_110593), _GEN_1123 & (_GEN_109960 | _GEN_1125 | _GEN_110125), _GEN_1117 & (_GEN_109492 | _GEN_1119 | _GEN_109657), _GEN_1111 & (_GEN_109024 | _GEN_1113 | _GEN_109189), _GEN_1105 & (_GEN_108556 | _GEN_1107 | _GEN_108721), _GEN_1099 & (_GEN_108088 | _GEN_1101 | _GEN_108253), _GEN_1093 & (_GEN_107620 | _GEN_1095 | _GEN_107785), _GEN_1087 & (_GEN_107152 | _GEN_1089 | _GEN_107317), _GEN_1081 & (_GEN_106684 | _GEN_1083 | _GEN_106849), _GEN_1075 & (_GEN_106216 | _GEN_1077 | _GEN_106381), _GEN_1069 & (_GEN_105748 | _GEN_1071 | _GEN_105913), _GEN_1063 & (_GEN_105280 | _GEN_1065 | _GEN_105445), _GEN_1057 & (_GEN_104812 | _GEN_1059 | _GEN_104977), _GEN_1051 & (_GEN_104344 | _GEN_1053 | _GEN_104509), _GEN_1045 & (_GEN_103876 | _GEN_1047 | _GEN_104041), _GEN_1039 & (_GEN_103408 | _GEN_1041 | _GEN_103573), _GEN_1033 & (_GEN_102940 | _GEN_1035 | _GEN_103105), _GEN_1027 & (_GEN_102472 | _GEN_1029 | _GEN_102637), _GEN_1021 & (_GEN_102004 | _GEN_1023 | _GEN_102169), _GEN_1015 & (_GEN_101536 | _GEN_1017 | _GEN_101701), _GEN_1009 & (_GEN_101068 | _GEN_1011 | _GEN_101233), _GEN_1003 & (_GEN_100600 | _GEN_1005 | _GEN_100765), _GEN_997 & (_GEN_100132 | _GEN_999 | _GEN_100297), _GEN_991 & (_GEN_99664 | _GEN_993 | _GEN_99829), _GEN_985 & (_GEN_99196 | _GEN_987 | _GEN_99361)}),
    .io_youngest_st_idx (do_st_search_0 ? (_lcam_stq_idx_T ? mem_stq_incoming_e_0_bits_uop_stq_idx : 5'h0) : _GEN_346 ? mem_ldq_incoming_e_0_bits_uop_stq_idx : 5'h0),
    .io_forwarding_idx  (_forwarding_age_logic_0_io_forwarding_idx)
  );
  ForwardingAgeLogic forwarding_age_logic_1 (
    .io_addr_matches    ({_GEN_1174 & (_GEN_113938 | _GEN_1176 | _GEN_113869), _GEN_1168 & (_GEN_113470 | _GEN_1170 | _GEN_113401), _GEN_1162 & (_GEN_113002 | _GEN_1164 | _GEN_112933), _GEN_1156 & (_GEN_112534 | _GEN_1158 | _GEN_112465), _GEN_1150 & (_GEN_112066 | _GEN_1152 | _GEN_111997), _GEN_1144 & (_GEN_111598 | _GEN_1146 | _GEN_111529), _GEN_1138 & (_GEN_111130 | _GEN_1140 | _GEN_111061), _GEN_1132 & (_GEN_110662 | _GEN_1134 | _GEN_110593), _GEN_1126 & (_GEN_110194 | _GEN_1128 | _GEN_110125), _GEN_1120 & (_GEN_109726 | _GEN_1122 | _GEN_109657), _GEN_1114 & (_GEN_109258 | _GEN_1116 | _GEN_109189), _GEN_1108 & (_GEN_108790 | _GEN_1110 | _GEN_108721), _GEN_1102 & (_GEN_108322 | _GEN_1104 | _GEN_108253), _GEN_1096 & (_GEN_107854 | _GEN_1098 | _GEN_107785), _GEN_1090 & (_GEN_107386 | _GEN_1092 | _GEN_107317), _GEN_1084 & (_GEN_106918 | _GEN_1086 | _GEN_106849), _GEN_1078 & (_GEN_106450 | _GEN_1080 | _GEN_106381), _GEN_1072 & (_GEN_105982 | _GEN_1074 | _GEN_105913), _GEN_1066 & (_GEN_105514 | _GEN_1068 | _GEN_105445), _GEN_1060 & (_GEN_105046 | _GEN_1062 | _GEN_104977), _GEN_1054 & (_GEN_104578 | _GEN_1056 | _GEN_104509), _GEN_1048 & (_GEN_104110 | _GEN_1050 | _GEN_104041), _GEN_1042 & (_GEN_103642 | _GEN_1044 | _GEN_103573), _GEN_1036 & (_GEN_103174 | _GEN_1038 | _GEN_103105), _GEN_1030 & (_GEN_102706 | _GEN_1032 | _GEN_102637), _GEN_1024 & (_GEN_102238 | _GEN_1026 | _GEN_102169), _GEN_1018 & (_GEN_101770 | _GEN_1020 | _GEN_101701), _GEN_1012 & (_GEN_101302 | _GEN_1014 | _GEN_101233), _GEN_1006 & (_GEN_100834 | _GEN_1008 | _GEN_100765), _GEN_1000 & (_GEN_100366 | _GEN_1002 | _GEN_100297), _GEN_994 & (_GEN_99898 | _GEN_996 | _GEN_99829), _GEN_988 & (_GEN_99430 | _GEN_990 | _GEN_99361)}),
    .io_youngest_st_idx (do_st_search_1 ? (_lcam_stq_idx_T_3 ? mem_stq_incoming_e_1_bits_uop_stq_idx : fired_sta_retry_1 ? mem_stq_retry_e_bits_uop_stq_idx : 5'h0) : do_ld_search_1 ? (fired_load_incoming_1 ? mem_ldq_incoming_e_1_bits_uop_stq_idx : fired_load_retry_1 ? mem_ldq_retry_e_bits_uop_stq_idx : fired_load_wakeup_1 ? mem_ldq_wakeup_e_bits_uop_stq_idx : 5'h0) : 5'h0),
    .io_forwarding_idx  (_forwarding_age_logic_1_io_forwarding_idx)
  );
  assign io_core_exe_0_iresp_valid = _io_core_exe_0_iresp_valid_output;
  assign io_core_exe_0_iresp_bits_uop_rob_idx = _GEN_1181 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_183 : casez_tmp_191) : casez_tmp_205;
  assign io_core_exe_0_iresp_bits_uop_pdst = _GEN_1181 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_186 : casez_tmp_193) : casez_tmp_208;
  assign io_core_exe_0_iresp_bits_uop_is_amo = _GEN_1181 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_188 : casez_tmp_194) : casez_tmp_210;
  assign io_core_exe_0_iresp_bits_uop_uses_stq = _GEN_1181 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_189 : casez_tmp_195) : casez_tmp_211;
  assign io_core_exe_0_iresp_bits_uop_dst_rtype = _GEN_1181 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_180 : casez_tmp_196) : casez_tmp_202;
  assign io_core_exe_0_iresp_bits_data = _GEN_1181 ? io_dmem_resp_0_bits_data : {_ldq_bits_debug_wb_data_T_19 ? {56{casez_tmp_209 & io_core_exe_0_iresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_10 ? {48{casez_tmp_209 & io_core_exe_0_iresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_1 ? {32{casez_tmp_209 & io_core_exe_0_iresp_bits_data_zeroed[31]}} : casez_tmp_200[63:32], io_core_exe_0_iresp_bits_data_zeroed[31:16]}, io_core_exe_0_iresp_bits_data_zeroed_1[15:8]}, io_core_exe_0_iresp_bits_data_zeroed_2};
  assign io_core_exe_0_fresp_valid = _io_core_exe_0_fresp_valid_output;
  assign io_core_exe_0_fresp_bits_uop_uopc = _GEN_1181 ? casez_tmp_181 : casez_tmp_204;
  assign io_core_exe_0_fresp_bits_uop_br_mask = _GEN_1181 ? casez_tmp_182 : casez_tmp_197;
  assign io_core_exe_0_fresp_bits_uop_rob_idx = _GEN_1181 ? casez_tmp_183 : casez_tmp_205;
  assign io_core_exe_0_fresp_bits_uop_stq_idx = _GEN_1181 ? casez_tmp_185 : casez_tmp_207;
  assign io_core_exe_0_fresp_bits_uop_pdst = _GEN_1181 ? casez_tmp_186 : casez_tmp_208;
  assign io_core_exe_0_fresp_bits_uop_mem_size = _GEN_1181 ? casez_tmp_187 : casez_tmp_201;
  assign io_core_exe_0_fresp_bits_uop_is_amo = _GEN_1181 ? casez_tmp_188 : casez_tmp_210;
  assign io_core_exe_0_fresp_bits_uop_uses_stq = _GEN_1181 ? casez_tmp_189 : casez_tmp_211;
  assign io_core_exe_0_fresp_bits_uop_dst_rtype = _GEN_1181 ? casez_tmp_180 : casez_tmp_202;
  assign io_core_exe_0_fresp_bits_uop_fp_val = _GEN_1181 ? casez_tmp_190 : casez_tmp_212;
  assign io_core_exe_0_fresp_bits_data = {1'h0, _GEN_1181 ? io_dmem_resp_0_bits_data : {_ldq_bits_debug_wb_data_T_19 ? {56{casez_tmp_209 & io_core_exe_0_fresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_10 ? {48{casez_tmp_209 & io_core_exe_0_fresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_1 ? {32{casez_tmp_209 & io_core_exe_0_fresp_bits_data_zeroed[31]}} : casez_tmp_200[63:32], io_core_exe_0_fresp_bits_data_zeroed[31:16]}, io_core_exe_0_fresp_bits_data_zeroed_1[15:8]}, io_core_exe_0_fresp_bits_data_zeroed_2}};
  assign io_core_exe_1_iresp_valid = _io_core_exe_1_iresp_valid_output;
  assign io_core_exe_1_iresp_bits_uop_rob_idx = _GEN_1185 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_216 : casez_tmp_224) : casez_tmp_238;
  assign io_core_exe_1_iresp_bits_uop_pdst = _GEN_1185 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_219 : casez_tmp_226) : casez_tmp_241;
  assign io_core_exe_1_iresp_bits_uop_is_amo = _GEN_1185 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_221 : casez_tmp_227) : casez_tmp_243;
  assign io_core_exe_1_iresp_bits_uop_uses_stq = _GEN_1185 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_222 : casez_tmp_228) : casez_tmp_244;
  assign io_core_exe_1_iresp_bits_uop_dst_rtype = _GEN_1185 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_213 : casez_tmp_229) : casez_tmp_235;
  assign io_core_exe_1_iresp_bits_data = _GEN_1185 ? io_dmem_resp_1_bits_data : {_ldq_bits_debug_wb_data_T_46 ? {56{casez_tmp_242 & io_core_exe_1_iresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_37 ? {48{casez_tmp_242 & io_core_exe_1_iresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_28 ? {32{casez_tmp_242 & io_core_exe_1_iresp_bits_data_zeroed[31]}} : casez_tmp_233[63:32], io_core_exe_1_iresp_bits_data_zeroed[31:16]}, io_core_exe_1_iresp_bits_data_zeroed_1[15:8]}, io_core_exe_1_iresp_bits_data_zeroed_2};
  assign io_core_exe_1_fresp_valid = _io_core_exe_1_fresp_valid_output;
  assign io_core_exe_1_fresp_bits_uop_uopc = _GEN_1185 ? casez_tmp_214 : casez_tmp_237;
  assign io_core_exe_1_fresp_bits_uop_br_mask = _GEN_1185 ? casez_tmp_215 : casez_tmp_230;
  assign io_core_exe_1_fresp_bits_uop_rob_idx = _GEN_1185 ? casez_tmp_216 : casez_tmp_238;
  assign io_core_exe_1_fresp_bits_uop_stq_idx = _GEN_1185 ? casez_tmp_218 : casez_tmp_240;
  assign io_core_exe_1_fresp_bits_uop_pdst = _GEN_1185 ? casez_tmp_219 : casez_tmp_241;
  assign io_core_exe_1_fresp_bits_uop_mem_size = _GEN_1185 ? casez_tmp_220 : casez_tmp_234;
  assign io_core_exe_1_fresp_bits_uop_is_amo = _GEN_1185 ? casez_tmp_221 : casez_tmp_243;
  assign io_core_exe_1_fresp_bits_uop_uses_stq = _GEN_1185 ? casez_tmp_222 : casez_tmp_244;
  assign io_core_exe_1_fresp_bits_uop_dst_rtype = _GEN_1185 ? casez_tmp_213 : casez_tmp_235;
  assign io_core_exe_1_fresp_bits_uop_fp_val = _GEN_1185 ? casez_tmp_223 : casez_tmp_245;
  assign io_core_exe_1_fresp_bits_data = {1'h0, _GEN_1185 ? io_dmem_resp_1_bits_data : {_ldq_bits_debug_wb_data_T_46 ? {56{casez_tmp_242 & io_core_exe_1_fresp_bits_data_zeroed_2[7]}} : {_ldq_bits_debug_wb_data_T_37 ? {48{casez_tmp_242 & io_core_exe_1_fresp_bits_data_zeroed_1[15]}} : {_ldq_bits_debug_wb_data_T_28 ? {32{casez_tmp_242 & io_core_exe_1_fresp_bits_data_zeroed[31]}} : casez_tmp_233[63:32], io_core_exe_1_fresp_bits_data_zeroed[31:16]}, io_core_exe_1_fresp_bits_data_zeroed_1[15:8]}, io_core_exe_1_fresp_bits_data_zeroed_2}};
  assign io_core_dis_ldq_idx_0 = ldq_tail;
  assign io_core_dis_ldq_idx_1 = _GEN_66;
  assign io_core_dis_ldq_idx_2 = _GEN_164;
  assign io_core_dis_ldq_idx_3 = _GEN_231;
  assign io_core_dis_stq_idx_0 = stq_tail;
  assign io_core_dis_stq_idx_1 = _ldq_T_35_bits_youngest_stq_idx;
  assign io_core_dis_stq_idx_2 = _ldq_T_75_bits_youngest_stq_idx;
  assign io_core_dis_stq_idx_3 = _ldq_T_115_bits_youngest_stq_idx;
  assign io_core_ldq_full_0 = _GEN_0 == ldq_head;
  assign io_core_ldq_full_1 = _GEN_67 == ldq_head;
  assign io_core_ldq_full_2 = _GEN_165 == ldq_head;
  assign io_core_ldq_full_3 = _GEN_232 == ldq_head;
  assign io_core_stq_full_0 = _GEN_1 == stq_head;
  assign io_core_stq_full_1 = _GEN_68 == stq_head;
  assign io_core_stq_full_2 = _GEN_166 == stq_head;
  assign io_core_stq_full_3 = _GEN_233 == stq_head;
  assign io_core_fp_stdata_ready = _io_core_fp_stdata_ready_output;
  assign io_core_clr_bsy_0_valid = clr_bsy_valid_0 & (io_core_brupdate_b1_mispredict_mask & clr_bsy_brmask_0) == 20'h0 & ~io_core_exception & ~io_core_clr_bsy_0_valid_REG & ~io_core_clr_bsy_0_valid_REG_2;
  assign io_core_clr_bsy_0_bits = clr_bsy_rob_idx_0;
  assign io_core_clr_bsy_1_valid = clr_bsy_valid_1 & (io_core_brupdate_b1_mispredict_mask & clr_bsy_brmask_1) == 20'h0 & ~io_core_exception & ~io_core_clr_bsy_1_valid_REG & ~io_core_clr_bsy_1_valid_REG_2;
  assign io_core_clr_bsy_1_bits = clr_bsy_rob_idx_1;
  assign io_core_clr_bsy_2_valid = stdf_clr_bsy_valid & (io_core_brupdate_b1_mispredict_mask & stdf_clr_bsy_brmask) == 20'h0 & ~io_core_exception & ~io_core_clr_bsy_2_valid_REG & ~io_core_clr_bsy_2_valid_REG_2;
  assign io_core_clr_bsy_2_bits = stdf_clr_bsy_rob_idx;
  assign io_core_spec_ld_wakeup_0_valid = _io_core_spec_ld_wakeup_0_valid_output;
  assign io_core_spec_ld_wakeup_0_bits = mem_incoming_uop_0_pdst;
  assign io_core_spec_ld_wakeup_1_valid = _io_core_spec_ld_wakeup_1_valid_output;
  assign io_core_spec_ld_wakeup_1_bits = mem_incoming_uop_1_pdst;
  assign io_core_ld_miss = ~((~spec_ld_succeed_REG | _io_core_exe_0_iresp_valid_output & (_GEN_1181 ? (io_dmem_resp_0_bits_uop_uses_ldq ? casez_tmp_184 : casez_tmp_192) : casez_tmp_206) == spec_ld_succeed_REG_1) & (~spec_ld_succeed_REG_2 | _io_core_exe_1_iresp_valid_output & (_GEN_1185 ? (io_dmem_resp_1_bits_uop_uses_ldq ? casez_tmp_217 : casez_tmp_225) : casez_tmp_239) == spec_ld_succeed_REG_3)) & io_core_ld_miss_REG;
  assign io_core_fencei_rdy = ~(stq_0_valid | stq_1_valid | stq_2_valid | stq_3_valid | stq_4_valid | stq_5_valid | stq_6_valid | stq_7_valid | stq_8_valid | stq_9_valid | stq_10_valid | stq_11_valid | stq_12_valid | stq_13_valid | stq_14_valid | stq_15_valid | stq_16_valid | stq_17_valid | stq_18_valid | stq_19_valid | stq_20_valid | stq_21_valid | stq_22_valid | stq_23_valid | stq_24_valid | stq_25_valid | stq_26_valid | stq_27_valid | stq_28_valid | stq_29_valid | stq_30_valid | stq_31_valid) & io_dmem_ordered;
  assign io_core_lxcpt_valid = r_xcpt_valid & ~io_core_exception & (io_core_brupdate_b1_mispredict_mask & r_xcpt_uop_br_mask) == 20'h0;
  assign io_core_lxcpt_bits_uop_br_mask = r_xcpt_uop_br_mask;
  assign io_core_lxcpt_bits_uop_rob_idx = r_xcpt_uop_rob_idx;
  assign io_core_lxcpt_bits_cause = r_xcpt_cause;
  assign io_core_lxcpt_bits_badvaddr = r_xcpt_badvaddr;
  assign io_dmem_req_valid = _io_dmem_req_valid_output;
  assign io_dmem_req_bits_0_valid = dmem_req_0_valid;
  assign io_dmem_req_bits_0_bits_uop_br_mask = can_fire_load_incoming_0 ? exe_tlb_uop_0_br_mask : will_fire_store_commit_0 ? casez_tmp_84 : 20'h0;
  assign io_dmem_req_bits_0_bits_uop_ldq_idx = can_fire_load_incoming_0 ? (_exe_tlb_uop_T_2 ? ldq_incoming_idx_0 : 5'h0) : will_fire_store_commit_0 ? casez_tmp_85 : 5'h0;
  assign io_dmem_req_bits_0_bits_uop_stq_idx = can_fire_load_incoming_0 ? (_exe_tlb_uop_T_2 ? stq_incoming_idx_0 : 5'h0) : will_fire_store_commit_0 ? casez_tmp_86 : 5'h0;
  assign io_dmem_req_bits_0_bits_uop_mem_cmd = can_fire_load_incoming_0 ? (_exe_tlb_uop_T_2 ? mem_incoming_uop_out_mem_cmd : 5'h0) : will_fire_store_commit_0 ? casez_tmp_87 : 5'h0;
  assign io_dmem_req_bits_0_bits_uop_mem_size = can_fire_load_incoming_0 ? (_exe_tlb_uop_T_2 ? mem_incoming_uop_out_mem_size : 2'h0) : will_fire_store_commit_0 ? casez_tmp_81 : 2'h0;
  assign io_dmem_req_bits_0_bits_uop_mem_signed = can_fire_load_incoming_0 ? _exe_tlb_uop_T_2 & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_mem_signed : io_core_exe_0_req_bits_uop_mem_signed) : will_fire_store_commit_0 & casez_tmp_88;
  assign io_dmem_req_bits_0_bits_uop_is_amo = can_fire_load_incoming_0 ? _exe_tlb_uop_T_2 & (io_core_exe_1_req_bits_sfence_valid ? io_core_exe_1_req_bits_uop_is_amo : io_core_exe_0_req_bits_uop_is_amo) : will_fire_store_commit_0 & casez_tmp_51;
  assign io_dmem_req_bits_0_bits_uop_uses_ldq = can_fire_load_incoming_0 ? exe_tlb_uop_0_uses_ldq : will_fire_store_commit_0 & casez_tmp_89;
  assign io_dmem_req_bits_0_bits_uop_uses_stq = can_fire_load_incoming_0 ? exe_tlb_uop_0_uses_stq : will_fire_store_commit_0 & casez_tmp_90;
  assign io_dmem_req_bits_0_bits_addr = can_fire_load_incoming_0 ? _GEN_334 : will_fire_store_commit_0 ? casez_tmp_80 : 40'h0;
  assign io_dmem_req_bits_0_bits_data = can_fire_load_incoming_0 | ~will_fire_store_commit_0 ? 64'h0 : casez_tmp_83;
  assign io_dmem_req_bits_1_valid = dmem_req_1_valid;
  assign io_dmem_req_bits_1_bits_uop_br_mask = can_fire_load_incoming_1 ? exe_tlb_uop_1_br_mask : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_br_mask : casez_tmp_67) : will_fire_load_wakeup_1 ? casez_tmp_92 : 20'h0;
  assign io_dmem_req_bits_1_bits_uop_ldq_idx = can_fire_load_incoming_1 ? (_exe_tlb_uop_T_9 ? ldq_incoming_idx_1 : will_fire_load_retry_1 ? casez_tmp_69 : will_fire_sta_retry_1 ? casez_tmp_58 : 5'h0) : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? ldq_incoming_idx_1 : casez_tmp_69) : will_fire_load_wakeup_1 ? casez_tmp_93 : 5'h0;
  assign io_dmem_req_bits_1_bits_uop_stq_idx = can_fire_load_incoming_1 ? (_exe_tlb_uop_T_9 ? stq_incoming_idx_1 : will_fire_load_retry_1 ? casez_tmp_70 : will_fire_sta_retry_1 ? casez_tmp_59 : 5'h0) : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? stq_incoming_idx_1 : casez_tmp_70) : will_fire_load_wakeup_1 ? casez_tmp_94 : 5'h0;
  assign io_dmem_req_bits_1_bits_uop_mem_cmd = can_fire_load_incoming_1 ? exe_tlb_uop_1_mem_cmd : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_mem_cmd : casez_tmp_72) : will_fire_load_wakeup_1 ? casez_tmp_95 : _GEN_336 ? hella_req_cmd : 5'h0;
  assign io_dmem_req_bits_1_bits_uop_mem_size = can_fire_load_incoming_1 ? exe_tlb_uop_1_mem_size : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_mem_size : casez_tmp_73) : will_fire_load_wakeup_1 ? casez_tmp_96 : _GEN_336 ? hella_req_size : 2'h0;
  assign io_dmem_req_bits_1_bits_uop_mem_signed = can_fire_load_incoming_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_mem_signed : will_fire_load_retry_1 ? casez_tmp_74 : will_fire_sta_retry_1 & casez_tmp_63) : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_mem_signed : casez_tmp_74) : will_fire_load_wakeup_1 ? casez_tmp_97 : _GEN_336 & hella_req_signed;
  assign io_dmem_req_bits_1_bits_uop_is_amo = can_fire_load_incoming_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_is_amo : will_fire_load_retry_1 ? casez_tmp_75 : will_fire_sta_retry_1 & casez_tmp_64) : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_is_amo : casez_tmp_75) : will_fire_load_wakeup_1 & casez_tmp_98;
  assign io_dmem_req_bits_1_bits_uop_uses_ldq = can_fire_load_incoming_1 ? exe_tlb_uop_1_uses_ldq : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_uses_ldq : casez_tmp_76) : will_fire_load_wakeup_1 & casez_tmp_99;
  assign io_dmem_req_bits_1_bits_uop_uses_stq = can_fire_load_incoming_1 ? exe_tlb_uop_1_uses_stq : will_fire_load_retry_1 ? (_exe_tlb_uop_T_9 ? exe_req_1_bits_uop_uses_stq : casez_tmp_77) : will_fire_load_wakeup_1 & casez_tmp_100;
  assign io_dmem_req_bits_1_bits_addr = _GEN_339 ? _GEN_338 : will_fire_load_wakeup_1 ? casez_tmp_91 : _GEN_337;
  assign io_dmem_req_bits_1_bits_data = _GEN_340 | will_fire_hella_incoming_1 | ~will_fire_hella_wakeup_1 ? 64'h0 : casez_tmp_101;
  assign io_dmem_req_bits_1_bits_is_hella = ~_GEN_340 & (will_fire_hella_incoming_1 | will_fire_hella_wakeup_1);
  assign io_dmem_s1_kill_0 = _GEN_1171 ? (_GEN_113704 ? io_dmem_s1_kill_0_REG_125 : _GEN_1173 ? io_dmem_s1_kill_0_REG_126 : _GEN_113869 ? io_dmem_s1_kill_0_REG_127 : _GEN_113272) : _GEN_113272;
  assign io_dmem_s1_kill_1 = _GEN_1174 ? (_GEN_113938 ? io_dmem_s1_kill_1_REG_125 : _GEN_1176 ? io_dmem_s1_kill_1_REG_126 : _GEN_113869 ? io_dmem_s1_kill_1_REG_127 : _GEN_113506) : _GEN_113506;
  assign io_dmem_brupdate_b1_resolve_mask = io_core_brupdate_b1_resolve_mask;
  assign io_dmem_brupdate_b1_mispredict_mask = io_core_brupdate_b1_mispredict_mask;
  assign io_dmem_exception = io_core_exception;
  assign io_dmem_release_ready = will_fire_release_1;
  assign io_dmem_force_order = _GEN & _GEN_139807 | io_core_fence_dmem;
  assign io_hellacache_req_ready = ~(|hella_state);
  assign io_hellacache_s2_nack = ~(~(|hella_state) | _GEN_140251) & _GEN_140233;
  assign io_hellacache_resp_valid = ~(~(|hella_state) | _GEN_140251 | _GEN_140233 | _GEN_330) & _GEN_331 & (_GEN_1231 | _GEN_140185);
  assign io_hellacache_resp_bits_data = _GEN_1231 ? io_dmem_resp_1_bits_data : io_dmem_resp_0_bits_data;
  assign io_hellacache_s2_xcpt_ae_ld = ~(~(|hella_state) | _GEN_140251 | _GEN_140233) & _GEN_330 & hella_xcpt_ae_ld;
endmodule

