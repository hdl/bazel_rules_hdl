// Standard header to adapt well known macros to our needs.

// Users can define 'PRINTF_COND' to add an extra gate to prints.
`ifndef PRINTF_COND_
  `ifdef PRINTF_COND
    `define PRINTF_COND_ (`PRINTF_COND)
  `else  // PRINTF_COND
    `define PRINTF_COND_ 1
  `endif // PRINTF_COND
`endif // not def PRINTF_COND_

module TileResetDomain(
  input          auto_boom_tile_buffer_out_a_ready,
                 auto_boom_tile_buffer_out_b_valid,
  input  [2:0]   auto_boom_tile_buffer_out_b_bits_opcode,
  input  [1:0]   auto_boom_tile_buffer_out_b_bits_param,
  input  [3:0]   auto_boom_tile_buffer_out_b_bits_size,
  input  [4:0]   auto_boom_tile_buffer_out_b_bits_source,
  input  [31:0]  auto_boom_tile_buffer_out_b_bits_address,
  input  [15:0]  auto_boom_tile_buffer_out_b_bits_mask,
  input          auto_boom_tile_buffer_out_b_bits_corrupt,
                 auto_boom_tile_buffer_out_c_ready,
                 auto_boom_tile_buffer_out_d_valid,
  input  [2:0]   auto_boom_tile_buffer_out_d_bits_opcode,
  input  [1:0]   auto_boom_tile_buffer_out_d_bits_param,
  input  [3:0]   auto_boom_tile_buffer_out_d_bits_size,
  input  [4:0]   auto_boom_tile_buffer_out_d_bits_source,
  input  [3:0]   auto_boom_tile_buffer_out_d_bits_sink,
  input          auto_boom_tile_buffer_out_d_bits_denied,
  input  [127:0] auto_boom_tile_buffer_out_d_bits_data,
  input          auto_boom_tile_buffer_out_d_bits_corrupt,
                 auto_boom_tile_buffer_out_e_ready,
                 auto_boom_tile_int_local_in_3_0,
                 auto_boom_tile_int_local_in_2_0,
                 auto_boom_tile_int_local_in_1_0,
                 auto_boom_tile_int_local_in_1_1,
                 auto_boom_tile_int_local_in_0_0,
                 auto_clock_in_clock,
                 auto_clock_in_reset,
  output         auto_boom_tile_buffer_out_a_valid,
  output [2:0]   auto_boom_tile_buffer_out_a_bits_opcode,
                 auto_boom_tile_buffer_out_a_bits_param,
  output [3:0]   auto_boom_tile_buffer_out_a_bits_size,
  output [4:0]   auto_boom_tile_buffer_out_a_bits_source,
  output [31:0]  auto_boom_tile_buffer_out_a_bits_address,
  output [15:0]  auto_boom_tile_buffer_out_a_bits_mask,
  output [127:0] auto_boom_tile_buffer_out_a_bits_data,
  output         auto_boom_tile_buffer_out_b_ready,
                 auto_boom_tile_buffer_out_c_valid,
  output [2:0]   auto_boom_tile_buffer_out_c_bits_opcode,
                 auto_boom_tile_buffer_out_c_bits_param,
  output [3:0]   auto_boom_tile_buffer_out_c_bits_size,
  output [4:0]   auto_boom_tile_buffer_out_c_bits_source,
  output [31:0]  auto_boom_tile_buffer_out_c_bits_address,
  output [127:0] auto_boom_tile_buffer_out_c_bits_data,
  output         auto_boom_tile_buffer_out_d_ready,
                 auto_boom_tile_buffer_out_e_valid,
  output [3:0]   auto_boom_tile_buffer_out_e_bits_sink
);

  BoomTile boom_tile (
    .clock                          (auto_clock_in_clock),
    .reset                          (auto_clock_in_reset),
    .auto_buffer_out_a_ready        (auto_boom_tile_buffer_out_a_ready),
    .auto_buffer_out_b_valid        (auto_boom_tile_buffer_out_b_valid),
    .auto_buffer_out_b_bits_opcode  (auto_boom_tile_buffer_out_b_bits_opcode),
    .auto_buffer_out_b_bits_param   (auto_boom_tile_buffer_out_b_bits_param),
    .auto_buffer_out_b_bits_size    (auto_boom_tile_buffer_out_b_bits_size),
    .auto_buffer_out_b_bits_source  (auto_boom_tile_buffer_out_b_bits_source),
    .auto_buffer_out_b_bits_address (auto_boom_tile_buffer_out_b_bits_address),
    .auto_buffer_out_b_bits_mask    (auto_boom_tile_buffer_out_b_bits_mask),
    .auto_buffer_out_b_bits_corrupt (auto_boom_tile_buffer_out_b_bits_corrupt),
    .auto_buffer_out_c_ready        (auto_boom_tile_buffer_out_c_ready),
    .auto_buffer_out_d_valid        (auto_boom_tile_buffer_out_d_valid),
    .auto_buffer_out_d_bits_opcode  (auto_boom_tile_buffer_out_d_bits_opcode),
    .auto_buffer_out_d_bits_param   (auto_boom_tile_buffer_out_d_bits_param),
    .auto_buffer_out_d_bits_size    (auto_boom_tile_buffer_out_d_bits_size),
    .auto_buffer_out_d_bits_source  (auto_boom_tile_buffer_out_d_bits_source),
    .auto_buffer_out_d_bits_sink    (auto_boom_tile_buffer_out_d_bits_sink),
    .auto_buffer_out_d_bits_denied  (auto_boom_tile_buffer_out_d_bits_denied),
    .auto_buffer_out_d_bits_data    (auto_boom_tile_buffer_out_d_bits_data),
    .auto_buffer_out_d_bits_corrupt (auto_boom_tile_buffer_out_d_bits_corrupt),
    .auto_buffer_out_e_ready        (auto_boom_tile_buffer_out_e_ready),
    .auto_int_local_in_3_0          (auto_boom_tile_int_local_in_3_0),
    .auto_int_local_in_2_0          (auto_boom_tile_int_local_in_2_0),
    .auto_int_local_in_1_0          (auto_boom_tile_int_local_in_1_0),
    .auto_int_local_in_1_1          (auto_boom_tile_int_local_in_1_1),
    .auto_int_local_in_0_0          (auto_boom_tile_int_local_in_0_0),
    .auto_buffer_out_a_valid        (auto_boom_tile_buffer_out_a_valid),
    .auto_buffer_out_a_bits_opcode  (auto_boom_tile_buffer_out_a_bits_opcode),
    .auto_buffer_out_a_bits_param   (auto_boom_tile_buffer_out_a_bits_param),
    .auto_buffer_out_a_bits_size    (auto_boom_tile_buffer_out_a_bits_size),
    .auto_buffer_out_a_bits_source  (auto_boom_tile_buffer_out_a_bits_source),
    .auto_buffer_out_a_bits_address (auto_boom_tile_buffer_out_a_bits_address),
    .auto_buffer_out_a_bits_mask    (auto_boom_tile_buffer_out_a_bits_mask),
    .auto_buffer_out_a_bits_data    (auto_boom_tile_buffer_out_a_bits_data),
    .auto_buffer_out_b_ready        (auto_boom_tile_buffer_out_b_ready),
    .auto_buffer_out_c_valid        (auto_boom_tile_buffer_out_c_valid),
    .auto_buffer_out_c_bits_opcode  (auto_boom_tile_buffer_out_c_bits_opcode),
    .auto_buffer_out_c_bits_param   (auto_boom_tile_buffer_out_c_bits_param),
    .auto_buffer_out_c_bits_size    (auto_boom_tile_buffer_out_c_bits_size),
    .auto_buffer_out_c_bits_source  (auto_boom_tile_buffer_out_c_bits_source),
    .auto_buffer_out_c_bits_address (auto_boom_tile_buffer_out_c_bits_address),
    .auto_buffer_out_c_bits_data    (auto_boom_tile_buffer_out_c_bits_data),
    .auto_buffer_out_d_ready        (auto_boom_tile_buffer_out_d_ready),
    .auto_buffer_out_e_valid        (auto_boom_tile_buffer_out_e_valid),
    .auto_buffer_out_e_bits_sink    (auto_boom_tile_buffer_out_e_bits_sink)
  );
endmodule

